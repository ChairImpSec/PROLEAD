module circuit ( plaintext1, plaintext2, plaintext3, key1, key2, key3,
        reset1, reset2, reset3, ciphertext, done, clk );
  input [127:0] plaintext1;
  input [127:0] plaintext2;
  input [127:0] plaintext3;
  input [127:0] key1;
  input [127:0] key2;
  input [127:0] key3;
  output [127:0] ciphertext;
  input reset1, reset2, reset3, clk;
  output done;
  wire   done1, done2, done3, inst1_n1297, inst1_n1296, inst1_n1295,
         inst1_n1294, inst1_n1293, inst1_n1292, inst1_n1291, inst1_n1290,
         inst1_n1289, inst1_n1288, inst1_n1287, inst1_n1286, inst1_n1285,
         inst1_n1284, inst1_n1283, inst1_n1282, inst1_n1281, inst1_n1280,
         inst1_n1279, inst1_n1278, inst1_n1277, inst1_n1276, inst1_n1275,
         inst1_n1274, inst1_n1273, inst1_n1272, inst1_n1271, inst1_n1270,
         inst1_n1269, inst1_n1268, inst1_n1267, inst1_n1266, inst1_n1265,
         inst1_n1264, inst1_n1263, inst1_n1262, inst1_n1261, inst1_n1260,
         inst1_n1259, inst1_n1258, inst1_n1257, inst1_n1256, inst1_n1255,
         inst1_n1254, inst1_n1253, inst1_n1252, inst1_n1251, inst1_n1250,
         inst1_n1249, inst1_n1248, inst1_n1247, inst1_n1246, inst1_n1245,
         inst1_n1244, inst1_n1243, inst1_n1242, inst1_n1241, inst1_n1240,
         inst1_n1239, inst1_n1238, inst1_n1237, inst1_n1236, inst1_n1235,
         inst1_n1234, inst1_n1233, inst1_n1232, inst1_n1231, inst1_n1230,
         inst1_n1229, inst1_n1228, inst1_n1227, inst1_n1226, inst1_n1225,
         inst1_n1224, inst1_n1223, inst1_n1222, inst1_n1221, inst1_n1220,
         inst1_n1219, inst1_n1218, inst1_n1217, inst1_n1216, inst1_n1215,
         inst1_n1214, inst1_n1213, inst1_n1212, inst1_n1211, inst1_n1210,
         inst1_n1209, inst1_n1208, inst1_n1207, inst1_n1206, inst1_n1205,
         inst1_n1204, inst1_n1203, inst1_n1202, inst1_n1201, inst1_n1200,
         inst1_n1199, inst1_n1198, inst1_n1197, inst1_n1196, inst1_n1195,
         inst1_n1194, inst1_n1193, inst1_n1192, inst1_n1191, inst1_n1190,
         inst1_n1187, inst1_n1186, inst1_n1185, inst1_n1184, inst1_n1183,
         inst1_n1182, inst1_n1181, inst1_n1180, inst1_n1179, inst1_n1178,
         inst1_n1177, inst1_n1176, inst1_n1175, inst1_n1174, inst1_n1173,
         inst1_n1172, inst1_n1171, inst1_n1170, inst1_n1169, inst1_n1168,
         inst1_n1167, inst1_n1166, inst1_n1165, inst1_n1164, inst1_n1163,
         inst1_n1162, inst1_n1161, inst1_n1160, inst1_n1159, inst1_n1158,
         inst1_n1157, inst1_n1156, inst1_n1155, inst1_n1154, inst1_n1153,
         inst1_n1152, inst1_n1151, inst1_n1150, inst1_n1149, inst1_n1148,
         inst1_n1147, inst1_n1146, inst1_n1145, inst1_n1144, inst1_n1143,
         inst1_n1142, inst1_n1141, inst1_n1140, inst1_n1139, inst1_n1138,
         inst1_n1137, inst1_n1136, inst1_n1135, inst1_n1134, inst1_n1133,
         inst1_n1132, inst1_n1131, inst1_n1130, inst1_n1129, inst1_n1128,
         inst1_n1127, inst1_n1126, inst1_n1125, inst1_n1124, inst1_n1123,
         inst1_n1120, inst1_n1117, inst1_n1112, inst1_n1108, inst1_n1107,
         inst1_n1104, inst1_n1101, inst1_n1099, inst1_n1095, inst1_n1083,
         inst1_n1078, inst1_n1069, inst1_n1068, inst1_n1066, inst1_n1065,
         inst1_n1064, inst1_n1063, inst1_n1062, inst1_n1053, inst1_n1045,
         inst1_n1043, inst1_n1042, inst1_n1041, inst1_n1040, inst1_n1039,
         inst1_n1038, inst1_n1037, inst1_n1036, inst1_n1035, inst1_n1034,
         inst1_n1033, inst1_n1032, inst1_n1031, inst1_n1030, inst1_n1029,
         inst1_n1028, inst1_n1027, inst1_n1026, inst1_n1025, inst1_n1024,
         inst1_n1023, inst1_n1022, inst1_n1021, inst1_n1020, inst1_n1019,
         inst1_n1018, inst1_n1017, inst1_n1016, inst1_n1015, inst1_n1014,
         inst1_n1013, inst1_n1012, inst1_n1011, inst1_n1010, inst1_n1009,
         inst1_n1008, inst1_n1007, inst1_n1006, inst1_n1005, inst1_n1004,
         inst1_n1003, inst1_n1002, inst1_n1001, inst1_n1000, inst1_n999,
         inst1_n998, inst1_n997, inst1_n996, inst1_n995, inst1_n994,
         inst1_n993, inst1_n992, inst1_n991, inst1_n990, inst1_n989,
         inst1_n988, inst1_n987, inst1_n986, inst1_n985, inst1_n984,
         inst1_n983, inst1_n982, inst1_n981, inst1_n931, inst1_n930,
         inst1_n929, inst1_n928, inst1_n927, inst1_n926, inst1_n925,
         inst1_n924, inst1_n907, inst1_n906, inst1_n905, inst1_n904,
         inst1_n903, inst1_n902, inst1_n901, inst1_n900, inst1_n899,
         inst1_n898, inst1_n897, inst1_n896, inst1_n895, inst1_n894,
         inst1_n893, inst1_n892, inst1_n867, inst1_n866, inst1_n865,
         inst1_n864, inst1_n863, inst1_n862, inst1_n861, inst1_n860,
         inst1_n859, inst1_n858, inst1_n857, inst1_n856, inst1_n855,
         inst1_n854, inst1_n853, inst1_n852, inst1_n850, inst1_n849,
         inst1_n848, inst1_n847, inst1_n846, inst1_n845, inst1_n844,
         inst1_n843, inst1_n842, inst1_n841, inst1_n840, inst1_n839,
         inst1_n838, inst1_n837, inst1_n836, inst1_n835, inst1_n834,
         inst1_n833, inst1_n832, inst1_n831, inst1_n830, inst1_n829,
         inst1_n828, inst1_n827, inst1_n826, inst1_n825, inst1_n824,
         inst1_n823, inst1_n822, inst1_n821, inst1_n820, inst1_n819,
         inst1_n818, inst1_n817, inst1_n816, inst1_n815, inst1_n814,
         inst1_n813, inst1_n812, inst1_n811, inst1_n810, inst1_n809,
         inst1_n808, inst1_n807, inst1_n806, inst1_n805, inst1_n804,
         inst1_n803, inst1_n802, inst1_n801, inst1_n800, inst1_n799,
         inst1_n798, inst1_n797, inst1_n796, inst1_n795, inst1_n794,
         inst1_n793, inst1_n792, inst1_n791, inst1_n790, inst1_n789,
         inst1_n788, inst1_n787, inst1_n786, inst1_n785, inst1_n784,
         inst1_n783, inst1_n782, inst1_n781, inst1_n780, inst1_n779,
         inst1_n778, inst1_n777, inst1_n776, inst1_n775, inst1_n774,
         inst1_n773, inst1_n772, inst1_n771, inst1_n770, inst1_n769,
         inst1_n768, inst1_n767, inst1_n766, inst1_n765, inst1_n764,
         inst1_n763, inst1_n762, inst1_n761, inst1_n760, inst1_n759,
         inst1_n758, inst1_n757, inst1_n756, inst1_n755, inst1_n754,
         inst1_n753, inst1_n752, inst1_n751, inst1_n750, inst1_n749,
         inst1_n748, inst1_n747, inst1_n746, inst1_n745, inst1_n744,
         inst1_n743, inst1_n742, inst1_n741, inst1_n740, inst1_n739,
         inst1_n738, inst1_n737, inst1_n736, inst1_n735, inst1_n734,
         inst1_n733, inst1_n732, inst1_n731, inst1_n730, inst1_n729,
         inst1_n728, inst1_n727, inst1_n726, inst1_n725, inst1_n724,
         inst1_n723, inst1_n722, inst1_n721, inst1_n720, inst1_n719,
         inst1_n718, inst1_n717, inst1_n716, inst1_n715, inst1_n714,
         inst1_n713, inst1_n712, inst1_n711, inst1_n710, inst1_n709,
         inst1_n708, inst1_n707, inst1_n706, inst1_n705, inst1_n704,
         inst1_n703, inst1_n702, inst1_n701, inst1_n700, inst1_n699,
         inst1_n698, inst1_n697, inst1_n696, inst1_n695, inst1_n694,
         inst1_n693, inst1_n692, inst1_n691, inst1_n690, inst1_n689,
         inst1_n688, inst1_n687, inst1_n686, inst1_n685, inst1_n684,
         inst1_n683, inst1_n682, inst1_n681, inst1_n680, inst1_n679,
         inst1_n678, inst1_n677, inst1_n676, inst1_n675, inst1_n674,
         inst1_n673, inst1_n672, inst1_n671, inst1_n670, inst1_n669,
         inst1_n668, inst1_n667, inst1_n666, inst1_n665, inst1_n664,
         inst1_n663, inst1_n662, inst1_n661, inst1_n660, inst1_n659,
         inst1_n658, inst1_n657, inst1_n656, inst1_n655, inst1_n654,
         inst1_n653, inst1_n652, inst1_n651, inst1_n650, inst1_n649,
         inst1_n648, inst1_n647, inst1_n646, inst1_n645, inst1_n644,
         inst1_n643, inst1_n642, inst1_n641, inst1_n640, inst1_n639,
         inst1_n638, inst1_n637, inst1_n636, inst1_n635, inst1_n634,
         inst1_n633, inst1_n632, inst1_n631, inst1_n630, inst1_n629,
         inst1_n628, inst1_n627, inst1_n626, inst1_n625, inst1_n624,
         inst1_n623, inst1_n622, inst1_n621, inst1_n620, inst1_n619,
         inst1_n618, inst1_n617, inst1_n616, inst1_n615, inst1_n614,
         inst1_n613, inst1_n612, inst1_n611, inst1_n610, inst1_n609,
         inst1_n608, inst1_n607, inst1_n606, inst1_n605, inst1_n604,
         inst1_n603, inst1_n602, inst1_n601, inst1_n600, inst1_n599,
         inst1_n598, inst1_n597, inst1_n596, inst1_n595, inst1_n594,
         inst1_n593, inst1_n592, inst1_n591, inst1_n590, inst1_n589,
         inst1_n588, inst1_n587, inst1_n586, inst1_n585, inst1_n584,
         inst1_n583, inst1_n582, inst1_n581, inst1_n580, inst1_n579,
         inst1_n578, inst1_n577, inst1_n576, inst1_n575, inst1_n574,
         inst1_n573, inst1_n572, inst1_n571, inst1_n570, inst1_n569,
         inst1_n568, inst1_n567, inst1_n566, inst1_n565, inst1_n564,
         inst1_n563, inst1_n562, inst1_n561, inst1_n560, inst1_n559,
         inst1_n558, inst1_n557, inst1_n556, inst1_n555, inst1_n554,
         inst1_n553, inst1_n552, inst1_n551, inst1_n550, inst1_n549,
         inst1_n548, inst1_n547, inst1_n546, inst1_n545, inst1_n544,
         inst1_n543, inst1_n542, inst1_n541, inst1_n540, inst1_n539,
         inst1_n538, inst1_n537, inst1_n536, inst1_n535, inst1_n534,
         inst1_n533, inst1_n532, inst1_n531, inst1_n530, inst1_n529,
         inst1_n528, inst1_n527, inst1_n526, inst1_n525, inst1_n524,
         inst1_n523, inst1_n522, inst1_n521, inst1_n520, inst1_n519,
         inst1_n518, inst1_n517, inst1_n516, inst1_n515, inst1_n514,
         inst1_n513, inst1_n512, inst1_n511, inst1_n510, inst1_n509,
         inst1_n508, inst1_n507, inst1_n506, inst1_n505, inst1_n504,
         inst1_n503, inst1_n502, inst1_n501, inst1_n500, inst1_n499,
         inst1_n498, inst1_n497, inst1_n496, inst1_n495, inst1_n494,
         inst1_n493, inst1_n492, inst1_n491, inst1_n490, inst1_n489,
         inst1_n488, inst1_n487, inst1_n486, inst1_n485, inst1_n484,
         inst1_n483, inst1_n482, inst1_n481, inst1_n480, inst1_n479,
         inst1_n478, inst1_n477, inst1_n476, inst1_n475, inst1_n474,
         inst1_n473, inst1_n472, inst1_n471, inst1_n470, inst1_n469,
         inst1_n468, inst1_n467, inst1_n466, inst1_n465, inst1_n464,
         inst1_n463, inst1_n462, inst1_n461, inst1_n460, inst1_n459,
         inst1_n458, inst1_n457, inst1_n456, inst1_n455, inst1_n454,
         inst1_n453, inst1_n452, inst1_n451, inst1_n450, inst1_n449,
         inst1_n448, inst1_n447, inst1_n446, inst1_n445, inst1_n444,
         inst1_n443, inst1_n442, inst1_n441, inst1_n440, inst1_n439,
         inst1_n438, inst1_n437, inst1_n436, inst1_n435, inst1_n434,
         inst1_n433, inst1_n432, inst1_n431, inst1_n430, inst1_n429,
         inst1_n428, inst1_n427, inst1_n426, inst1_n425, inst1_n424,
         inst1_n423, inst1_n422, inst1_n421, inst1_n420, inst1_n419,
         inst1_n418, inst1_n417, inst1_n416, inst1_n415, inst1_n414,
         inst1_n413, inst1_n412, inst1_n411, inst1_n410, inst1_n409,
         inst1_n408, inst1_n407, inst1_n406, inst1_n405, inst1_n404,
         inst1_n403, inst1_n402, inst1_n401, inst1_n400, inst1_n399,
         inst1_n398, inst1_n397, inst1_n396, inst1_n395, inst1_n394,
         inst1_n393, inst1_n392, inst1_n391, inst1_n390, inst1_n389,
         inst1_n388, inst1_n387, inst1_n386, inst1_n385, inst1_n384,
         inst1_n383, inst1_n382, inst1_n381, inst1_n380, inst1_n379,
         inst1_n378, inst1_n377, inst1_n376, inst1_n375, inst1_n374,
         inst1_n373, inst1_n372, inst1_n371, inst1_n370, inst1_n369,
         inst1_n368, inst1_n367, inst1_n366, inst1_n365, inst1_n364,
         inst1_n363, inst1_n362, inst1_n361, inst1_n360, inst1_n359,
         inst1_n358, inst1_n357, inst1_n356, inst1_n355, inst1_n354,
         inst1_n353, inst1_n352, inst1_n351, inst1_n350, inst1_n349,
         inst1_n348, inst1_n347, inst1_n346, inst1_n345, inst1_n344,
         inst1_n343, inst1_n342, inst1_n341, inst1_n340, inst1_n339,
         inst1_n338, inst1_n337, inst1_n336, inst1_n335, inst1_n334,
         inst1_n333, inst1_n332, inst1_n331, inst1_n330, inst1_n329,
         inst1_n328, inst1_n327, inst1_n326, inst1_n325, inst1_n324,
         inst1_n323, inst1_n322, inst1_n321, inst1_n320, inst1_n319,
         inst1_n318, inst1_n317, inst1_n316, inst1_n315, inst1_n314,
         inst1_n313, inst1_n312, inst1_n311, inst1_n310, inst1_n309,
         inst1_n308, inst1_n307, inst1_n306, inst1_n305, inst1_n304,
         inst1_n303, inst1_n302, inst1_n301, inst1_n300, inst1_n299,
         inst1_n298, inst1_n297, inst1_n296, inst1_n295, inst1_n294,
         inst1_n293, inst1_n292, inst1_n291, inst1_n290, inst1_n289,
         inst1_n288, inst1_n287, inst1_n286, inst1_n285, inst1_n284,
         inst1_n283, inst1_n282, inst1_n281, inst1_n280, inst1_n279,
         inst1_n278, inst1_n277, inst1_n276, inst1_n275, inst1_n274,
         inst1_n273, inst1_n272, inst1_n271, inst1_n270, inst1_n269,
         inst1_n268, inst1_n267, inst1_n266, inst1_n265, inst1_n264,
         inst1_n263, inst1_n262, inst1_n261, inst1_n260, inst1_n259,
         inst1_n258, inst1_n257, inst1_n256, inst1_n255, inst1_n254,
         inst1_n253, inst1_n252, inst1_n251, inst1_n250, inst1_n249,
         inst1_n248, inst1_n247, inst1_n246, inst1_n245, inst1_n244,
         inst1_n243, inst1_n242, inst1_n241, inst1_n240, inst1_n239,
         inst1_n238, inst1_n237, inst1_n236, inst1_n235, inst1_n234,
         inst1_n233, inst1_n232, inst1_n231, inst1_n230, inst1_n229,
         inst1_n228, inst1_n227, inst1_n226, inst1_n225, inst1_n224,
         inst1_n223, inst1_n222, inst1_n221, inst1_n220, inst1_n219,
         inst1_n218, inst1_n217, inst1_n216, inst1_n215, inst1_n214,
         inst1_n213, inst1_n212, inst1_n211, inst1_n210, inst1_n209,
         inst1_n208, inst1_n207, inst1_n206, inst1_n205, inst1_n204,
         inst1_n203, inst1_n202, inst1_n201, inst1_n200, inst1_n199,
         inst1_n198, inst1_n197, inst1_n196, inst1_n195, inst1_n194,
         inst1_n193, inst1_n192, inst1_n191, inst1_n190, inst1_n189,
         inst1_n188, inst1_n1189, inst1_n1188, inst1_n143, inst1_n137,
         inst1_n136, inst1_n135, inst1_n134, inst1_n133, inst1_n132,
         inst1_n131, inst1_n130, inst1_n129, inst1_n128, inst1_n127,
         inst1_n126, inst1_n125, inst1_n124, inst1_n123, inst1_n122,
         inst1_n121, inst1_n120, inst1_n119, inst1_n118, inst1_n117,
         inst1_n116, inst1_n115, inst1_n114, inst1_n113, inst1_n112,
         inst1_n111, inst1_n110, inst1_n109, inst1_n108, inst1_n107, inst1_n98,
         inst1_n97, inst1_n96, inst1_n95, inst1_n94, inst1_n93, inst1_n92,
         inst1_n91, inst1_n90, inst1_n89, inst1_n88, inst1_n87, inst1_n86,
         inst1_n85, inst1_n84, inst1_n83, inst1_n82, inst1_n81, inst1_n80,
         inst1_n79, inst1_n78, inst1_n77, inst1_n76, inst1_n75, inst1_n74,
         inst1_n73, inst1_n72, inst1_n71, inst1_n70, inst1_n69, inst1_n68,
         inst1_n67, inst1_n65, inst1_n57, inst1_n24, inst1_n22, inst1_n17,
         inst1_n14, inst1_n12, inst1_n11, inst1_n10, inst1_n9, inst1_n6,
         inst1_n1122, inst1_n1121, inst1_n1119, inst1_n1118, inst1_n1116,
         inst1_n1115, inst1_n1114, inst1_n1113, inst1_n1111, inst1_n1110,
         inst1_n1109, inst1_n1106, inst1_n1105, inst1_n1103, inst1_n1102,
         inst1_n1100, inst1_n1098, inst1_n1097, inst1_n1096, inst1_n1094,
         inst1_n1093, inst1_n1092, inst1_n1091, inst1_n1090, inst1_n1089,
         inst1_n1088, inst1_n1087, inst1_n1086, inst1_n1085, inst1_n1084,
         inst1_n1082, inst1_n1081, inst1_n1080, inst1_n1079, inst1_n1077,
         inst1_n1076, inst1_n1075, inst1_n1074, inst1_n1073, inst1_n1072,
         inst1_n1071, inst1_n1070, inst1_n1061, inst1_n1060, inst1_n1059,
         inst1_n1058, inst1_n1057, inst1_n1056, inst1_n1055, inst1_n1054,
         inst1_n1052, inst1_n1051, inst1_n1050, inst1_n1049, inst1_n1048,
         inst1_n1047, inst1_n1046, inst1_n1044, inst1_n980, inst1_n979,
         inst1_n978, inst1_n977, inst1_n976, inst1_n975, inst1_n974,
         inst1_n973, inst1_n972, inst1_n971, inst1_n970, inst1_n969,
         inst1_n968, inst1_n967, inst1_n966, inst1_n965, inst1_n964,
         inst1_n963, inst1_n962, inst1_n961, inst1_n960, inst1_n959,
         inst1_n958, inst1_n957, inst1_n956, inst1_n955, inst1_n954,
         inst1_n953, inst1_n952, inst1_n951, inst1_n950, inst1_n949,
         inst1_n948, inst1_n947, inst1_n946, inst1_n945, inst1_n944,
         inst1_n943, inst1_n942, inst1_n941, inst1_n940, inst1_n939,
         inst1_n938, inst1_n937, inst1_n936, inst1_n935, inst1_n934,
         inst1_n933, inst1_n932, inst1_n923, inst1_n922, inst1_n921,
         inst1_n920, inst1_n919, inst1_n918, inst1_n917, inst1_n916,
         inst1_n915, inst1_n914, inst1_n913, inst1_n912, inst1_n911,
         inst1_n910, inst1_n909, inst1_n908, inst1_n891, inst1_n890,
         inst1_n889, inst1_n888, inst1_n887, inst1_n886, inst1_n885,
         inst1_n884, inst1_n883, inst1_n882, inst1_n881, inst1_n880,
         inst1_n879, inst1_n878, inst1_n877, inst1_n876, inst1_n875,
         inst1_n874, inst1_n873, inst1_n872, inst1_n871, inst1_n870,
         inst1_n869, inst1_n868, inst1_n851, inst1_calcRCon_n44,
         inst1_calcRCon_n45, inst1_calcRCon_n46, inst1_calcRCon_n47,
         inst1_calcRCon_n48, inst1_calcRCon_n49, inst1_calcRCon_n50,
         inst1_calcRCon_n51, inst1_KeyArray_S33reg_gff_1_SFF_7_n5,
         inst1_KeyArray_S33reg_gff_1_SFF_6_n5,
         inst1_KeyArray_S33reg_gff_1_SFF_5_n5,
         inst1_KeyArray_S33reg_gff_1_SFF_4_n5,
         inst1_KeyArray_S33reg_gff_1_SFF_3_n5,
         inst1_KeyArray_S33reg_gff_1_SFF_2_n5,
         inst1_KeyArray_S33reg_gff_1_SFF_1_n5,
         inst1_KeyArray_S33reg_gff_1_SFF_0_n5,
         inst1_KeyArray_S32reg_gff_1_SFF_7_n5,
         inst1_KeyArray_S32reg_gff_1_SFF_6_n5,
         inst1_KeyArray_S32reg_gff_1_SFF_5_n5,
         inst1_KeyArray_S32reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S32reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S32reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S32reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S32reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S31reg_gff_1_SFF_7_n6,
         inst1_KeyArray_S31reg_gff_1_SFF_6_n6,
         inst1_KeyArray_S31reg_gff_1_SFF_5_n6,
         inst1_KeyArray_S31reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S31reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S31reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S31reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S31reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S30reg_gff_1_SFF_7_n6,
         inst1_KeyArray_S30reg_gff_1_SFF_6_n6,
         inst1_KeyArray_S30reg_gff_1_SFF_5_n6,
         inst1_KeyArray_S30reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S30reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S30reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S30reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S30reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S23reg_gff_1_SFF_7_n5,
         inst1_KeyArray_S23reg_gff_1_SFF_6_n5,
         inst1_KeyArray_S23reg_gff_1_SFF_5_n5,
         inst1_KeyArray_S23reg_gff_1_SFF_4_n5,
         inst1_KeyArray_S23reg_gff_1_SFF_3_n5,
         inst1_KeyArray_S23reg_gff_1_SFF_2_n5,
         inst1_KeyArray_S23reg_gff_1_SFF_1_n5,
         inst1_KeyArray_S23reg_gff_1_SFF_0_n5,
         inst1_KeyArray_S22reg_gff_1_SFF_7_n5,
         inst1_KeyArray_S22reg_gff_1_SFF_6_n5,
         inst1_KeyArray_S22reg_gff_1_SFF_5_n5,
         inst1_KeyArray_S22reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S22reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S22reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S22reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S22reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S21reg_gff_1_SFF_7_n6,
         inst1_KeyArray_S21reg_gff_1_SFF_6_n6,
         inst1_KeyArray_S21reg_gff_1_SFF_5_n6,
         inst1_KeyArray_S21reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S21reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S21reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S21reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S21reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S20reg_gff_1_SFF_7_n6,
         inst1_KeyArray_S20reg_gff_1_SFF_6_n6,
         inst1_KeyArray_S20reg_gff_1_SFF_5_n6,
         inst1_KeyArray_S20reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S20reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S20reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S20reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S20reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S13reg_gff_1_SFF_7_n5,
         inst1_KeyArray_S13reg_gff_1_SFF_6_n5,
         inst1_KeyArray_S13reg_gff_1_SFF_5_n5,
         inst1_KeyArray_S13reg_gff_1_SFF_4_n5,
         inst1_KeyArray_S13reg_gff_1_SFF_3_n5,
         inst1_KeyArray_S13reg_gff_1_SFF_2_n5,
         inst1_KeyArray_S13reg_gff_1_SFF_1_n5,
         inst1_KeyArray_S13reg_gff_1_SFF_0_n5,
         inst1_KeyArray_S12reg_gff_1_SFF_7_n5,
         inst1_KeyArray_S12reg_gff_1_SFF_6_n5,
         inst1_KeyArray_S12reg_gff_1_SFF_5_n5,
         inst1_KeyArray_S12reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S12reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S12reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S12reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S12reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S11reg_gff_1_SFF_7_n6,
         inst1_KeyArray_S11reg_gff_1_SFF_6_n6,
         inst1_KeyArray_S11reg_gff_1_SFF_5_n6,
         inst1_KeyArray_S11reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S11reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S11reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S11reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S11reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S10reg_gff_1_SFF_7_n6,
         inst1_KeyArray_S10reg_gff_1_SFF_6_n6,
         inst1_KeyArray_S10reg_gff_1_SFF_5_n6,
         inst1_KeyArray_S10reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S10reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S10reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S10reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S10reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S03reg_gff_1_SFF_7_n5,
         inst1_KeyArray_S03reg_gff_1_SFF_6_n5,
         inst1_KeyArray_S03reg_gff_1_SFF_5_n5,
         inst1_KeyArray_S03reg_gff_1_SFF_4_n5,
         inst1_KeyArray_S03reg_gff_1_SFF_3_n5,
         inst1_KeyArray_S03reg_gff_1_SFF_2_n5,
         inst1_KeyArray_S03reg_gff_1_SFF_1_n5,
         inst1_KeyArray_S03reg_gff_1_SFF_0_n5,
         inst1_KeyArray_S02reg_gff_1_SFF_7_n5,
         inst1_KeyArray_S02reg_gff_1_SFF_6_n5,
         inst1_KeyArray_S02reg_gff_1_SFF_5_n5,
         inst1_KeyArray_S02reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S02reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S02reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S02reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S02reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S01reg_gff_1_SFF_7_n6,
         inst1_KeyArray_S01reg_gff_1_SFF_6_n6,
         inst1_KeyArray_S01reg_gff_1_SFF_5_n6,
         inst1_KeyArray_S01reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S01reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S01reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S01reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S01reg_gff_1_SFF_0_n6,
         inst1_KeyArray_S00reg_gff_1_SFF_7_n6,
         inst1_KeyArray_S00reg_gff_1_SFF_6_n6,
         inst1_KeyArray_S00reg_gff_1_SFF_5_n6,
         inst1_KeyArray_S00reg_gff_1_SFF_4_n6,
         inst1_KeyArray_S00reg_gff_1_SFF_3_n6,
         inst1_KeyArray_S00reg_gff_1_SFF_2_n6,
         inst1_KeyArray_S00reg_gff_1_SFF_1_n6,
         inst1_KeyArray_S00reg_gff_1_SFF_0_n6,
         inst1_stateArray_S33reg_gff_1_SFF_7_n5,
         inst1_stateArray_S33reg_gff_1_SFF_6_n5,
         inst1_stateArray_S33reg_gff_1_SFF_5_n5,
         inst1_stateArray_S33reg_gff_1_SFF_4_n5,
         inst1_stateArray_S33reg_gff_1_SFF_3_n5,
         inst1_stateArray_S33reg_gff_1_SFF_2_n5,
         inst1_stateArray_S33reg_gff_1_SFF_1_n5,
         inst1_stateArray_S33reg_gff_1_SFF_0_n5,
         inst1_stateArray_S32reg_gff_1_SFF_7_n5,
         inst1_stateArray_S32reg_gff_1_SFF_6_n5,
         inst1_stateArray_S32reg_gff_1_SFF_5_n5,
         inst1_stateArray_S32reg_gff_1_SFF_4_n6,
         inst1_stateArray_S32reg_gff_1_SFF_3_n6,
         inst1_stateArray_S32reg_gff_1_SFF_2_n6,
         inst1_stateArray_S32reg_gff_1_SFF_1_n6,
         inst1_stateArray_S32reg_gff_1_SFF_0_n6,
         inst1_stateArray_S31reg_gff_1_SFF_7_n6,
         inst1_stateArray_S31reg_gff_1_SFF_6_n6,
         inst1_stateArray_S31reg_gff_1_SFF_5_n6,
         inst1_stateArray_S31reg_gff_1_SFF_4_n6,
         inst1_stateArray_S31reg_gff_1_SFF_3_n6,
         inst1_stateArray_S31reg_gff_1_SFF_2_n6,
         inst1_stateArray_S31reg_gff_1_SFF_1_n6,
         inst1_stateArray_S31reg_gff_1_SFF_0_n6,
         inst1_stateArray_S30reg_gff_1_SFF_7_n5,
         inst1_stateArray_S30reg_gff_1_SFF_6_n5,
         inst1_stateArray_S30reg_gff_1_SFF_5_n5,
         inst1_stateArray_S30reg_gff_1_SFF_4_n5,
         inst1_stateArray_S30reg_gff_1_SFF_3_n5,
         inst1_stateArray_S30reg_gff_1_SFF_2_n5,
         inst1_stateArray_S30reg_gff_1_SFF_1_n5,
         inst1_stateArray_S30reg_gff_1_SFF_0_n5,
         inst1_stateArray_S23reg_gff_1_SFF_7_n5,
         inst1_stateArray_S23reg_gff_1_SFF_6_n5,
         inst1_stateArray_S23reg_gff_1_SFF_5_n5,
         inst1_stateArray_S23reg_gff_1_SFF_4_n6,
         inst1_stateArray_S23reg_gff_1_SFF_3_n6,
         inst1_stateArray_S23reg_gff_1_SFF_2_n6,
         inst1_stateArray_S23reg_gff_1_SFF_1_n6,
         inst1_stateArray_S23reg_gff_1_SFF_0_n6,
         inst1_stateArray_S22reg_gff_1_SFF_7_n6,
         inst1_stateArray_S22reg_gff_1_SFF_6_n6,
         inst1_stateArray_S22reg_gff_1_SFF_5_n6,
         inst1_stateArray_S22reg_gff_1_SFF_4_n6,
         inst1_stateArray_S22reg_gff_1_SFF_3_n6,
         inst1_stateArray_S22reg_gff_1_SFF_2_n6,
         inst1_stateArray_S22reg_gff_1_SFF_1_n6,
         inst1_stateArray_S22reg_gff_1_SFF_0_n6,
         inst1_stateArray_S21reg_gff_1_SFF_7_n6,
         inst1_stateArray_S21reg_gff_1_SFF_6_n6,
         inst1_stateArray_S21reg_gff_1_SFF_5_n6,
         inst1_stateArray_S21reg_gff_1_SFF_4_n6,
         inst1_stateArray_S21reg_gff_1_SFF_3_n6,
         inst1_stateArray_S21reg_gff_1_SFF_2_n6,
         inst1_stateArray_S21reg_gff_1_SFF_1_n6,
         inst1_stateArray_S21reg_gff_1_SFF_0_n6,
         inst1_stateArray_S20reg_gff_1_SFF_7_n5,
         inst1_stateArray_S20reg_gff_1_SFF_6_n5,
         inst1_stateArray_S20reg_gff_1_SFF_5_n5,
         inst1_stateArray_S20reg_gff_1_SFF_4_n5,
         inst1_stateArray_S20reg_gff_1_SFF_3_n5,
         inst1_stateArray_S20reg_gff_1_SFF_2_n5,
         inst1_stateArray_S20reg_gff_1_SFF_1_n5,
         inst1_stateArray_S20reg_gff_1_SFF_0_n5,
         inst1_stateArray_S13reg_gff_1_SFF_7_n5,
         inst1_stateArray_S13reg_gff_1_SFF_6_n5,
         inst1_stateArray_S13reg_gff_1_SFF_5_n5,
         inst1_stateArray_S13reg_gff_1_SFF_4_n6,
         inst1_stateArray_S13reg_gff_1_SFF_3_n6,
         inst1_stateArray_S13reg_gff_1_SFF_2_n6,
         inst1_stateArray_S13reg_gff_1_SFF_1_n6,
         inst1_stateArray_S13reg_gff_1_SFF_0_n6,
         inst1_stateArray_S12reg_gff_1_SFF_7_n6,
         inst1_stateArray_S12reg_gff_1_SFF_6_n6,
         inst1_stateArray_S12reg_gff_1_SFF_5_n6,
         inst1_stateArray_S12reg_gff_1_SFF_4_n6,
         inst1_stateArray_S12reg_gff_1_SFF_3_n6,
         inst1_stateArray_S12reg_gff_1_SFF_2_n6,
         inst1_stateArray_S12reg_gff_1_SFF_1_n6,
         inst1_stateArray_S12reg_gff_1_SFF_0_n6,
         inst1_stateArray_S11reg_gff_1_SFF_7_n6,
         inst1_stateArray_S11reg_gff_1_SFF_6_n6,
         inst1_stateArray_S11reg_gff_1_SFF_5_n6,
         inst1_stateArray_S11reg_gff_1_SFF_4_n6,
         inst1_stateArray_S11reg_gff_1_SFF_3_n6,
         inst1_stateArray_S11reg_gff_1_SFF_2_n6,
         inst1_stateArray_S11reg_gff_1_SFF_1_n6,
         inst1_stateArray_S11reg_gff_1_SFF_0_n6,
         inst1_stateArray_S10reg_gff_1_SFF_7_n5,
         inst1_stateArray_S10reg_gff_1_SFF_6_n5,
         inst1_stateArray_S10reg_gff_1_SFF_5_n5,
         inst1_stateArray_S10reg_gff_1_SFF_4_n5,
         inst1_stateArray_S10reg_gff_1_SFF_3_n5,
         inst1_stateArray_S10reg_gff_1_SFF_2_n5,
         inst1_stateArray_S10reg_gff_1_SFF_1_n5,
         inst1_stateArray_S10reg_gff_1_SFF_0_n5,
         inst1_stateArray_S03reg_gff_1_SFF_7_n5,
         inst1_stateArray_S03reg_gff_1_SFF_6_n5,
         inst1_stateArray_S03reg_gff_1_SFF_5_n5,
         inst1_stateArray_S03reg_gff_1_SFF_4_n6,
         inst1_stateArray_S03reg_gff_1_SFF_3_n6,
         inst1_stateArray_S03reg_gff_1_SFF_2_n6,
         inst1_stateArray_S03reg_gff_1_SFF_1_n6,
         inst1_stateArray_S03reg_gff_1_SFF_0_n6,
         inst1_stateArray_S02reg_gff_1_SFF_7_n6,
         inst1_stateArray_S02reg_gff_1_SFF_6_n6,
         inst1_stateArray_S02reg_gff_1_SFF_5_n6,
         inst1_stateArray_S02reg_gff_1_SFF_4_n6,
         inst1_stateArray_S02reg_gff_1_SFF_3_n6,
         inst1_stateArray_S02reg_gff_1_SFF_2_n6,
         inst1_stateArray_S02reg_gff_1_SFF_1_n6,
         inst1_stateArray_S02reg_gff_1_SFF_0_n6,
         inst1_stateArray_S01reg_gff_1_SFF_7_n6,
         inst1_stateArray_S01reg_gff_1_SFF_6_n6,
         inst1_stateArray_S01reg_gff_1_SFF_5_n6,
         inst1_stateArray_S01reg_gff_1_SFF_4_n6,
         inst1_stateArray_S01reg_gff_1_SFF_3_n6,
         inst1_stateArray_S01reg_gff_1_SFF_2_n6,
         inst1_stateArray_S01reg_gff_1_SFF_1_n6,
         inst1_stateArray_S01reg_gff_1_SFF_0_n6,
         inst1_stateArray_S00reg_gff_1_SFF_7_n6,
         inst1_stateArray_S00reg_gff_1_SFF_6_n6,
         inst1_stateArray_S00reg_gff_1_SFF_5_n6,
         inst1_stateArray_S00reg_gff_1_SFF_4_n6,
         inst1_stateArray_S00reg_gff_1_SFF_3_n6,
         inst1_stateArray_S00reg_gff_1_SFF_2_n6,
         inst1_stateArray_S00reg_gff_1_SFF_1_n6,
         inst1_stateArray_S00reg_gff_1_SFF_0_n6, inst1_ctrl_seq4_SFF_1_n5,
         inst1_ctrl_seq4_SFF_0_n5, inst1_ctrl_seq6_SFF_4_n5,
         inst1_ctrl_seq6_SFF_3_n5, inst1_ctrl_seq6_SFF_2_n5,
         inst1_ctrl_seq6_SFF_1_n5, inst1_ctrl_seq6_SFF_0_n5, inst1_ctrl_n6,
         inst2_n2872, inst2_n2871, inst2_n2870, inst2_n2869, inst2_n2868,
         inst2_n2867, inst2_n2866, inst2_n2865, inst2_n2864, inst2_n2863,
         inst2_n2862, inst2_n2861, inst2_n2860, inst2_n2859, inst2_n2858,
         inst2_n2857, inst2_n2856, inst2_n2855, inst2_n2854, inst2_n2853,
         inst2_n2852, inst2_n2851, inst2_n2850, inst2_n2849, inst2_n2848,
         inst2_n2847, inst2_n2846, inst2_n2845, inst2_n2844, inst2_n2843,
         inst2_n2842, inst2_n2841, inst2_n2840, inst2_n2839, inst2_n2838,
         inst2_n2837, inst2_n2836, inst2_n2835, inst2_n2834, inst2_n2833,
         inst2_n2832, inst2_n2831, inst2_n2830, inst2_n2829, inst2_n2828,
         inst2_n2827, inst2_n2826, inst2_n2825, inst2_n2824, inst2_n2823,
         inst2_n2822, inst2_n2821, inst2_n2820, inst2_n2819, inst2_n2818,
         inst2_n2817, inst2_n2816, inst2_n2815, inst2_n2814, inst2_n2813,
         inst2_n2812, inst2_n2811, inst2_n2810, inst2_n2809, inst2_n2808,
         inst2_n2807, inst2_n2806, inst2_n2805, inst2_n2804, inst2_n2803,
         inst2_n2802, inst2_n2801, inst2_n2800, inst2_n2799, inst2_n2798,
         inst2_n2797, inst2_n2796, inst2_n2795, inst2_n2794, inst2_n2793,
         inst2_n2792, inst2_n2791, inst2_n2790, inst2_n2789, inst2_n2788,
         inst2_n2787, inst2_n2786, inst2_n2785, inst2_n2784, inst2_n2783,
         inst2_n2782, inst2_n2781, inst2_n2780, inst2_n2779, inst2_n2778,
         inst2_n2777, inst2_n2776, inst2_n2775, inst2_n2774, inst2_n2773,
         inst2_n2772, inst2_n2771, inst2_n2770, inst2_n2769, inst2_n2768,
         inst2_n2767, inst2_n2766, inst2_n2765, inst2_n2764, inst2_n2763,
         inst2_n2762, inst2_n2761, inst2_n2760, inst2_n2759, inst2_n2758,
         inst2_n2757, inst2_n2756, inst2_n2755, inst2_n2754, inst2_n2753,
         inst2_n2752, inst2_n2751, inst2_n2750, inst2_n2749, inst2_n2748,
         inst2_n2747, inst2_n2746, inst2_n2745, inst2_n2744, inst2_n2743,
         inst2_n2742, inst2_n2741, inst2_n2740, inst2_n2739, inst2_n2738,
         inst2_n2737, inst2_n2736, inst2_n2735, inst2_n2734, inst2_n2733,
         inst2_n2732, inst2_n2731, inst2_n2730, inst2_n2729, inst2_n2728,
         inst2_n2727, inst2_n2726, inst2_n2725, inst2_n2724, inst2_n2723,
         inst2_n2722, inst2_n2721, inst2_n2720, inst2_n2719, inst2_n2718,
         inst2_n2717, inst2_n2716, inst2_n2715, inst2_n2714, inst2_n2713,
         inst2_n2712, inst2_n2711, inst2_n2710, inst2_n2709, inst2_n2708,
         inst2_n2707, inst2_n2706, inst2_n2705, inst2_n2704, inst2_n2703,
         inst2_n2702, inst2_n2701, inst2_n2700, inst2_n2699, inst2_n2698,
         inst2_n2697, inst2_n2696, inst2_n2695, inst2_n2694, inst2_n2693,
         inst2_n2692, inst2_n2691, inst2_n2690, inst2_n2689, inst2_n2688,
         inst2_n2687, inst2_n2685, inst2_n2684, inst2_n2683, inst2_n2682,
         inst2_n2681, inst2_n2680, inst2_n2679, inst2_n2678, inst2_n2677,
         inst2_n2676, inst2_n2675, inst2_n2674, inst2_n2673, inst2_n2672,
         inst2_n2671, inst2_n2670, inst2_n2669, inst2_n2668, inst2_n2667,
         inst2_n2666, inst2_n2665, inst2_n2664, inst2_n2663, inst2_n2662,
         inst2_n2661, inst2_n2660, inst2_n2659, inst2_n2658, inst2_n2657,
         inst2_n2656, inst2_n2655, inst2_n2654, inst2_n2653, inst2_n2652,
         inst2_n2651, inst2_n2650, inst2_n2649, inst2_n2648, inst2_n2647,
         inst2_n2646, inst2_n2645, inst2_n2644, inst2_n2643, inst2_n2642,
         inst2_n2641, inst2_n2640, inst2_n2639, inst2_n2638, inst2_n2637,
         inst2_n2636, inst2_n2635, inst2_n2634, inst2_n2633, inst2_n2632,
         inst2_n2631, inst2_n2630, inst2_n2629, inst2_n2628, inst2_n2627,
         inst2_n2626, inst2_n2625, inst2_n2624, inst2_n2623, inst2_n2622,
         inst2_n2621, inst2_n2620, inst2_n2619, inst2_n2618, inst2_n2617,
         inst2_n2616, inst2_n2615, inst2_n2614, inst2_n2613, inst2_n2612,
         inst2_n2611, inst2_n2610, inst2_n2609, inst2_n2608, inst2_n2607,
         inst2_n2606, inst2_n2605, inst2_n2604, inst2_n2603, inst2_n2602,
         inst2_n2601, inst2_n2600, inst2_n2599, inst2_n2598, inst2_n2597,
         inst2_n2596, inst2_n2595, inst2_n2594, inst2_n2593, inst2_n2592,
         inst2_n2591, inst2_n2590, inst2_n2589, inst2_n2588, inst2_n2587,
         inst2_n2586, inst2_n2585, inst2_n2584, inst2_n2583, inst2_n2582,
         inst2_n2581, inst2_n2580, inst2_n2579, inst2_n2578, inst2_n2577,
         inst2_n2576, inst2_n2575, inst2_n2574, inst2_n2573, inst2_n2572,
         inst2_n2571, inst2_n2570, inst2_n2569, inst2_n2568, inst2_n2567,
         inst2_n2566, inst2_n2565, inst2_n2564, inst2_n2563, inst2_n2562,
         inst2_n2561, inst2_n2560, inst2_n2559, inst2_n2558, inst2_n2557,
         inst2_n2556, inst2_n2555, inst2_n2554, inst2_n2553, inst2_n2552,
         inst2_n2551, inst2_n2550, inst2_n2549, inst2_n2548, inst2_n2547,
         inst2_n2546, inst2_n2545, inst2_n2544, inst2_n2543, inst2_n2542,
         inst2_n2541, inst2_n2540, inst2_n2539, inst2_n2538, inst2_n2537,
         inst2_n2536, inst2_n2535, inst2_n2534, inst2_n2533, inst2_n2532,
         inst2_n2531, inst2_n2530, inst2_n2529, inst2_n2528, inst2_n2527,
         inst2_n2526, inst2_n2525, inst2_n2524, inst2_n2523, inst2_n2522,
         inst2_n2521, inst2_n2520, inst2_n2519, inst2_n2518, inst2_n2517,
         inst2_n2516, inst2_n2515, inst2_n2514, inst2_n2513, inst2_n2512,
         inst2_n2511, inst2_n2510, inst2_n2509, inst2_n2508, inst2_n2507,
         inst2_n2506, inst2_n2505, inst2_n2504, inst2_n2503, inst2_n2502,
         inst2_n2501, inst2_n2500, inst2_n2499, inst2_n2498, inst2_n2497,
         inst2_n2496, inst2_n2495, inst2_n2494, inst2_n2493, inst2_n2492,
         inst2_n2491, inst2_n2490, inst2_n2489, inst2_n2488, inst2_n2487,
         inst2_n2486, inst2_n2485, inst2_n2484, inst2_n2483, inst2_n2482,
         inst2_n2481, inst2_n2480, inst2_n2479, inst2_n2478, inst2_n2477,
         inst2_n2476, inst2_n2475, inst2_n2474, inst2_n2473, inst2_n2472,
         inst2_n2471, inst2_n2470, inst2_n2469, inst2_n2468, inst2_n2467,
         inst2_n2466, inst2_n2465, inst2_n2464, inst2_n2463, inst2_n2462,
         inst2_n2461, inst2_n2460, inst2_n2459, inst2_n2458, inst2_n2457,
         inst2_n2456, inst2_n2455, inst2_n2454, inst2_n2453, inst2_n2452,
         inst2_n2451, inst2_n2450, inst2_n2449, inst2_n2448, inst2_n2447,
         inst2_n2446, inst2_n2445, inst2_n2444, inst2_n2443, inst2_n2442,
         inst2_n2441, inst2_n2440, inst2_n2439, inst2_n2438, inst2_n2437,
         inst2_n2436, inst2_n2435, inst2_n2434, inst2_n2433, inst2_n2432,
         inst2_n2431, inst2_n2430, inst2_n2429, inst2_n2428, inst2_n2427,
         inst2_n2426, inst2_n2425, inst2_n2424, inst2_n2423, inst2_n2422,
         inst2_n2421, inst2_n2420, inst2_n2419, inst2_n2418, inst2_n2417,
         inst2_n2416, inst2_n2415, inst2_n2414, inst2_n2413, inst2_n2412,
         inst2_n2411, inst2_n2410, inst2_n2409, inst2_n2408, inst2_n2407,
         inst2_n2406, inst2_n2405, inst2_n2404, inst2_n2403, inst2_n2402,
         inst2_n2401, inst2_n2400, inst2_n2399, inst2_n2398, inst2_n2397,
         inst2_n2396, inst2_n2395, inst2_n2394, inst2_n2393, inst2_n2392,
         inst2_n2391, inst2_n2390, inst2_n2389, inst2_n2388, inst2_n2387,
         inst2_n2386, inst2_n2385, inst2_n2384, inst2_n2383, inst2_n2382,
         inst2_n2381, inst2_n2380, inst2_n2379, inst2_n2378, inst2_n2377,
         inst2_n2376, inst2_n2375, inst2_n2374, inst2_n2373, inst2_n2372,
         inst2_n2371, inst2_n2370, inst2_n2369, inst2_n2368, inst2_n2367,
         inst2_n2366, inst2_n2365, inst2_n2364, inst2_n2363, inst2_n2362,
         inst2_n2361, inst2_n2360, inst2_n2359, inst2_n2358, inst2_n2357,
         inst2_n2356, inst2_n2355, inst2_n2354, inst2_n2353, inst2_n2352,
         inst2_n2351, inst2_n2350, inst2_n2349, inst2_n2348, inst2_n2347,
         inst2_n2346, inst2_n2345, inst2_n2344, inst2_n2343, inst2_n2342,
         inst2_n2341, inst2_n2340, inst2_n2339, inst2_n2338, inst2_n2337,
         inst2_n2336, inst2_n2335, inst2_n2334, inst2_n2333, inst2_n2332,
         inst2_n2331, inst2_n2330, inst2_n2329, inst2_n2328, inst2_n2327,
         inst2_n2326, inst2_n2325, inst2_n2324, inst2_n2323, inst2_n2322,
         inst2_n2321, inst2_n2320, inst2_n2319, inst2_n2318, inst2_n2317,
         inst2_n2316, inst2_n2315, inst2_n2314, inst2_n2313, inst2_n2312,
         inst2_n2311, inst2_n2310, inst2_n2309, inst2_n2308, inst2_n2307,
         inst2_n2306, inst2_n2305, inst2_n2304, inst2_n2303, inst2_n2302,
         inst2_n2301, inst2_n2300, inst2_n2299, inst2_n2298, inst2_n2297,
         inst2_n2296, inst2_n2295, inst2_n2294, inst2_n2293, inst2_n2292,
         inst2_n2291, inst2_n2290, inst2_n2289, inst2_n2288, inst2_n2287,
         inst2_n2286, inst2_n2285, inst2_n2284, inst2_n2283, inst2_n2282,
         inst2_n2281, inst2_n2280, inst2_n2279, inst2_n2278, inst2_n2277,
         inst2_n2276, inst2_n2275, inst2_n2274, inst2_n2273, inst2_n2272,
         inst2_n2271, inst2_n2270, inst2_n2269, inst2_n2268, inst2_n2267,
         inst2_n2266, inst2_n2265, inst2_n2264, inst2_n2263, inst2_n2262,
         inst2_n2261, inst2_n2260, inst2_n2259, inst2_n2258, inst2_n2257,
         inst2_n2256, inst2_n2255, inst2_n2254, inst2_n2253, inst2_n2252,
         inst2_n2251, inst2_n2250, inst2_n2249, inst2_n2248, inst2_n2247,
         inst2_n2246, inst2_n2245, inst2_n2244, inst2_n2243, inst2_n2242,
         inst2_n2241, inst2_n2240, inst2_n2239, inst2_n2238, inst2_n2237,
         inst2_n2236, inst2_n2235, inst2_n2234, inst2_n2233, inst2_n2232,
         inst2_n2231, inst2_n2230, inst2_n2229, inst2_n2228, inst2_n2227,
         inst2_n2226, inst2_n2225, inst2_n2224, inst2_n2223, inst2_n2222,
         inst2_n2221, inst2_n2220, inst2_n2219, inst2_n2218, inst2_n2217,
         inst2_n2216, inst2_n2215, inst2_n2214, inst2_n2213, inst2_n2212,
         inst2_n2211, inst2_n2210, inst2_n2209, inst2_n2208, inst2_n2207,
         inst2_n2206, inst2_n2205, inst2_n2204, inst2_n2203, inst2_n2202,
         inst2_n2201, inst2_n2200, inst2_n2199, inst2_n2198, inst2_n2197,
         inst2_n2196, inst2_n2195, inst2_n2194, inst2_n2193, inst2_n2192,
         inst2_n2191, inst2_n2190, inst2_n2189, inst2_n2188, inst2_n2187,
         inst2_n2186, inst2_n2185, inst2_n2184, inst2_n2183, inst2_n2182,
         inst2_n2181, inst2_n2180, inst2_n2179, inst2_n2178, inst2_n2177,
         inst2_n2176, inst2_n2175, inst2_n2174, inst2_n2173, inst2_n2172,
         inst2_n2171, inst2_n2170, inst2_n2169, inst2_n2168, inst2_n2167,
         inst2_n2166, inst2_n2165, inst2_n2164, inst2_n2163, inst2_n2162,
         inst2_n2161, inst2_n2160, inst2_n2159, inst2_n2158, inst2_n2157,
         inst2_n2156, inst2_n2155, inst2_n2154, inst2_n2153, inst2_n2152,
         inst2_n2151, inst2_n2150, inst2_n2149, inst2_n2148, inst2_n2147,
         inst2_n2146, inst2_n2145, inst2_n2144, inst2_n2143, inst2_n2142,
         inst2_n2141, inst2_n2140, inst2_n2139, inst2_n2138, inst2_n2137,
         inst2_n2136, inst2_n2135, inst2_n2134, inst2_n2133, inst2_n2132,
         inst2_n2131, inst2_n2130, inst2_n2129, inst2_n2128, inst2_n2127,
         inst2_n2126, inst2_n2125, inst2_n2124, inst2_n2123, inst2_n2122,
         inst2_n2121, inst2_n2120, inst2_n2119, inst2_n2118, inst2_n2117,
         inst2_n2116, inst2_n2115, inst2_n2114, inst2_n2113, inst2_n2112,
         inst2_n2111, inst2_n2110, inst2_n2109, inst2_n2108, inst2_n2107,
         inst2_n2106, inst2_n2105, inst2_n2104, inst2_n2103, inst2_n2102,
         inst2_n2101, inst2_n2100, inst2_n2099, inst2_n2098, inst2_n2097,
         inst2_n2096, inst2_n2095, inst2_n2094, inst2_n2093, inst2_n2092,
         inst2_n2091, inst2_n2090, inst2_n2089, inst2_n2088, inst2_n2087,
         inst2_n2086, inst2_n2085, inst2_n2084, inst2_n2083, inst2_n2082,
         inst2_n2081, inst2_n2080, inst2_n2079, inst2_n2078, inst2_n2077,
         inst2_n2076, inst2_n2075, inst2_n2074, inst2_n2073, inst2_n2072,
         inst2_n2071, inst2_n2070, inst2_n2069, inst2_n2068, inst2_n2067,
         inst2_n2066, inst2_n2065, inst2_n2064, inst2_n2063, inst2_n2062,
         inst2_n2061, inst2_n2060, inst2_n2059, inst2_n2058, inst2_n2057,
         inst2_n2056, inst2_n2055, inst2_n2054, inst2_n2053, inst2_n2052,
         inst2_n2051, inst2_n2050, inst2_n2049, inst2_n2048, inst2_n2047,
         inst2_n2046, inst2_n2045, inst2_n2044, inst2_n2043, inst2_n2042,
         inst2_n2041, inst2_n2040, inst2_n2039, inst2_n2038, inst2_n2037,
         inst2_n2036, inst2_n2035, inst2_n2034, inst2_n2033, inst2_n2032,
         inst2_n2031, inst2_n2030, inst2_n2029, inst2_n2028, inst2_n2027,
         inst2_n2026, inst2_n2025, inst2_n2024, inst2_n2023, inst2_n2022,
         inst2_n2021, inst2_n2020, inst2_n2019, inst2_n2018, inst2_n2017,
         inst2_n2016, inst2_n2015, inst2_n2014, inst2_n2013, inst2_n2012,
         inst2_n2011, inst2_n2010, inst2_n2009, inst2_n2008, inst2_n2007,
         inst2_n2006, inst2_n2005, inst2_n2004, inst2_n2003, inst2_n2002,
         inst2_n2001, inst2_n2000, inst2_n1999, inst2_n1998, inst2_n1997,
         inst2_n1996, inst2_n1995, inst2_n1994, inst2_n1993, inst2_n1992,
         inst2_n1991, inst2_n1990, inst2_n1989, inst2_n1988, inst2_n1987,
         inst2_n1986, inst2_n1985, inst2_n1984, inst2_n1983, inst2_n1982,
         inst2_n1981, inst2_n1980, inst2_n1979, inst2_n1978, inst2_n1977,
         inst2_n1976, inst2_n1975, inst2_n1974, inst2_n1973, inst2_n1972,
         inst2_n1971, inst2_n1970, inst2_n1969, inst2_n1968, inst2_n1967,
         inst2_n1966, inst2_n1965, inst2_n1964, inst2_n1963, inst2_n1962,
         inst2_n1961, inst2_n1960, inst2_n1959, inst2_n1958, inst2_n1957,
         inst2_n1956, inst2_n1955, inst2_n1954, inst2_n1953, inst2_n1952,
         inst2_n1951, inst2_n1950, inst2_n1949, inst2_n1948, inst2_n1947,
         inst2_n1946, inst2_n1945, inst2_n1944, inst2_n1943, inst2_n1942,
         inst2_n1941, inst2_n1940, inst2_n1939, inst2_n1938, inst2_n1937,
         inst2_n1936, inst2_n1935, inst2_n1934, inst2_n1933, inst2_n1932,
         inst2_n1931, inst2_n1930, inst2_n1929, inst2_n1928, inst2_n1927,
         inst2_n1926, inst2_n1925, inst2_n1924, inst2_n1923, inst2_n1922,
         inst2_n1921, inst2_n1920, inst2_n1919, inst2_n1918, inst2_n1917,
         inst2_n1916, inst2_n1915, inst2_n1914, inst2_n1096, inst2_n1088,
         inst2_n1290, inst2_n1273, inst2_n1272, inst2_n1271, inst2_n1270,
         inst2_n1269, inst2_n1268, inst2_n1267, inst2_n1266, inst2_n1265,
         inst2_n1264, inst2_n1263, inst2_n1262, inst2_n1261, inst2_n1260,
         inst2_n1259, inst2_n1258, inst2_n1257, inst2_n1256, inst2_n1255,
         inst2_n1254, inst2_n1253, inst2_n1252, inst2_n1251, inst2_n1250,
         inst2_n1233, inst2_n1232, inst2_n1231, inst2_n1230, inst2_n1229,
         inst2_n1228, inst2_n1227, inst2_n1226, inst2_n1225, inst2_n1224,
         inst2_n1223, inst2_n1222, inst2_n1221, inst2_n1220, inst2_n1219,
         inst2_n1218, inst2_n1209, inst2_n1208, inst2_n1207, inst2_n1206,
         inst2_n1205, inst2_n1204, inst2_n1203, inst2_n1202, inst2_n1201,
         inst2_n1200, inst2_n1199, inst2_n1198, inst2_n1197, inst2_n1196,
         inst2_n1195, inst2_n1194, inst2_n1193, inst2_n1192, inst2_n1191,
         inst2_n1190, inst2_n1189, inst2_n1188, inst2_n1187, inst2_n1186,
         inst2_n1185, inst2_n1184, inst2_n1183, inst2_n1182, inst2_n1181,
         inst2_n1180, inst2_n1179, inst2_n1178, inst2_n1177, inst2_n1176,
         inst2_n1175, inst2_n1174, inst2_n1173, inst2_n1172, inst2_n1171,
         inst2_n1170, inst2_n1169, inst2_n1168, inst2_n1167, inst2_n1166,
         inst2_n1165, inst2_n1164, inst2_n1163, inst2_n1162, inst2_n1161,
         inst2_n1097, inst2_n1095, inst2_n1094, inst2_n1093, inst2_n1092,
         inst2_n1091, inst2_n1090, inst2_n1089, inst2_n1087, inst2_n1086,
         inst2_n1085, inst2_n1084, inst2_n1083, inst2_n1082, inst2_n1081,
         inst2_n1080, inst2_n1071, inst2_n718, inst2_n706, inst2_n581,
         inst2_n499, inst2_n444, inst2_n321, inst2_n236, inst2_n233,
         inst2_n232, inst2_n231, inst2_n230, inst2_n228, inst2_n227,
         inst2_n226, inst2_n225, inst2_n224, inst2_n223, inst2_n222,
         inst2_n221, inst2_n220, inst2_n219, inst2_n218, inst2_n216,
         inst2_n215, inst2_n214, inst2_n212, inst2_n210, inst2_n209,
         inst2_n207, inst2_n206, inst2_n203, inst2_n202, inst2_n201,
         inst2_n199, inst2_n198, inst2_n197, inst2_n196, inst2_n194,
         inst2_n193, inst2_n191, inst2_n190, inst2_n143, inst2_n137,
         inst2_n136, inst2_n135, inst2_n134, inst2_n133, inst2_n132,
         inst2_n131, inst2_n130, inst2_n129, inst2_n128, inst2_n127,
         inst2_n126, inst2_n125, inst2_n124, inst2_n123, inst2_n122,
         inst2_n121, inst2_n120, inst2_n119, inst2_n118, inst2_n117,
         inst2_n116, inst2_n115, inst2_n114, inst2_n113, inst2_n112,
         inst2_n111, inst2_n110, inst2_n109, inst2_n108, inst2_n107, inst2_n98,
         inst2_n97, inst2_n96, inst2_n95, inst2_n94, inst2_n93, inst2_n92,
         inst2_n91, inst2_n90, inst2_n89, inst2_n88, inst2_n87, inst2_n86,
         inst2_n85, inst2_n84, inst2_n83, inst2_n82, inst2_n81, inst2_n80,
         inst2_n79, inst2_n78, inst2_n77, inst2_n76, inst2_n75, inst2_n74,
         inst2_n73, inst2_n72, inst2_n71, inst2_n70, inst2_n69, inst2_n68,
         inst2_n67, inst2_n65, inst2_n57, inst2_n24, inst2_n22, inst2_n17,
         inst2_n14, inst2_n12, inst2_n11, inst2_n10, inst2_n9, inst2_n6,
         inst2_calcRCon_n44, inst2_calcRCon_n45, inst2_calcRCon_n46,
         inst2_calcRCon_n47, inst2_calcRCon_n48, inst2_calcRCon_n49,
         inst2_calcRCon_n50, inst2_calcRCon_n51,
         inst2_KeyArray_S33reg_gff_1_SFF_7_n5,
         inst2_KeyArray_S33reg_gff_1_SFF_6_n5,
         inst2_KeyArray_S33reg_gff_1_SFF_5_n5,
         inst2_KeyArray_S33reg_gff_1_SFF_4_n5,
         inst2_KeyArray_S33reg_gff_1_SFF_3_n5,
         inst2_KeyArray_S33reg_gff_1_SFF_2_n5,
         inst2_KeyArray_S33reg_gff_1_SFF_1_n5,
         inst2_KeyArray_S33reg_gff_1_SFF_0_n5,
         inst2_KeyArray_S32reg_gff_1_SFF_7_n5,
         inst2_KeyArray_S32reg_gff_1_SFF_6_n5,
         inst2_KeyArray_S32reg_gff_1_SFF_5_n5,
         inst2_KeyArray_S32reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S32reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S32reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S32reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S32reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S31reg_gff_1_SFF_7_n6,
         inst2_KeyArray_S31reg_gff_1_SFF_6_n6,
         inst2_KeyArray_S31reg_gff_1_SFF_5_n6,
         inst2_KeyArray_S31reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S31reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S31reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S31reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S31reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S30reg_gff_1_SFF_7_n6,
         inst2_KeyArray_S30reg_gff_1_SFF_6_n6,
         inst2_KeyArray_S30reg_gff_1_SFF_5_n6,
         inst2_KeyArray_S30reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S30reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S30reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S30reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S30reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S23reg_gff_1_SFF_7_n5,
         inst2_KeyArray_S23reg_gff_1_SFF_6_n5,
         inst2_KeyArray_S23reg_gff_1_SFF_5_n5,
         inst2_KeyArray_S23reg_gff_1_SFF_4_n5,
         inst2_KeyArray_S23reg_gff_1_SFF_3_n5,
         inst2_KeyArray_S23reg_gff_1_SFF_2_n5,
         inst2_KeyArray_S23reg_gff_1_SFF_1_n5,
         inst2_KeyArray_S23reg_gff_1_SFF_0_n5,
         inst2_KeyArray_S22reg_gff_1_SFF_7_n5,
         inst2_KeyArray_S22reg_gff_1_SFF_6_n5,
         inst2_KeyArray_S22reg_gff_1_SFF_5_n5,
         inst2_KeyArray_S22reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S22reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S22reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S22reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S22reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S21reg_gff_1_SFF_7_n6,
         inst2_KeyArray_S21reg_gff_1_SFF_6_n6,
         inst2_KeyArray_S21reg_gff_1_SFF_5_n6,
         inst2_KeyArray_S21reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S21reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S21reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S21reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S21reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S20reg_gff_1_SFF_7_n6,
         inst2_KeyArray_S20reg_gff_1_SFF_6_n6,
         inst2_KeyArray_S20reg_gff_1_SFF_5_n6,
         inst2_KeyArray_S20reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S20reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S20reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S20reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S20reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S13reg_gff_1_SFF_7_n5,
         inst2_KeyArray_S13reg_gff_1_SFF_6_n5,
         inst2_KeyArray_S13reg_gff_1_SFF_5_n5,
         inst2_KeyArray_S13reg_gff_1_SFF_4_n5,
         inst2_KeyArray_S13reg_gff_1_SFF_3_n5,
         inst2_KeyArray_S13reg_gff_1_SFF_2_n5,
         inst2_KeyArray_S13reg_gff_1_SFF_1_n5,
         inst2_KeyArray_S13reg_gff_1_SFF_0_n5,
         inst2_KeyArray_S12reg_gff_1_SFF_7_n5,
         inst2_KeyArray_S12reg_gff_1_SFF_6_n5,
         inst2_KeyArray_S12reg_gff_1_SFF_5_n5,
         inst2_KeyArray_S12reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S12reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S12reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S12reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S12reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S11reg_gff_1_SFF_7_n6,
         inst2_KeyArray_S11reg_gff_1_SFF_6_n6,
         inst2_KeyArray_S11reg_gff_1_SFF_5_n6,
         inst2_KeyArray_S11reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S11reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S11reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S11reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S11reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S10reg_gff_1_SFF_7_n6,
         inst2_KeyArray_S10reg_gff_1_SFF_6_n6,
         inst2_KeyArray_S10reg_gff_1_SFF_5_n6,
         inst2_KeyArray_S10reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S10reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S10reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S10reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S10reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S03reg_gff_1_SFF_7_n5,
         inst2_KeyArray_S03reg_gff_1_SFF_6_n5,
         inst2_KeyArray_S03reg_gff_1_SFF_5_n5,
         inst2_KeyArray_S03reg_gff_1_SFF_4_n5,
         inst2_KeyArray_S03reg_gff_1_SFF_3_n5,
         inst2_KeyArray_S03reg_gff_1_SFF_2_n5,
         inst2_KeyArray_S03reg_gff_1_SFF_1_n5,
         inst2_KeyArray_S03reg_gff_1_SFF_0_n5,
         inst2_KeyArray_S02reg_gff_1_SFF_7_n5,
         inst2_KeyArray_S02reg_gff_1_SFF_6_n5,
         inst2_KeyArray_S02reg_gff_1_SFF_5_n5,
         inst2_KeyArray_S02reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S02reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S02reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S02reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S02reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S01reg_gff_1_SFF_7_n6,
         inst2_KeyArray_S01reg_gff_1_SFF_6_n6,
         inst2_KeyArray_S01reg_gff_1_SFF_5_n6,
         inst2_KeyArray_S01reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S01reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S01reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S01reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S01reg_gff_1_SFF_0_n6,
         inst2_KeyArray_S00reg_gff_1_SFF_7_n6,
         inst2_KeyArray_S00reg_gff_1_SFF_6_n6,
         inst2_KeyArray_S00reg_gff_1_SFF_5_n6,
         inst2_KeyArray_S00reg_gff_1_SFF_4_n6,
         inst2_KeyArray_S00reg_gff_1_SFF_3_n6,
         inst2_KeyArray_S00reg_gff_1_SFF_2_n6,
         inst2_KeyArray_S00reg_gff_1_SFF_1_n6,
         inst2_KeyArray_S00reg_gff_1_SFF_0_n6,
         inst2_stateArray_S33reg_gff_1_SFF_7_n5,
         inst2_stateArray_S33reg_gff_1_SFF_6_n5,
         inst2_stateArray_S33reg_gff_1_SFF_5_n5,
         inst2_stateArray_S33reg_gff_1_SFF_4_n5,
         inst2_stateArray_S33reg_gff_1_SFF_3_n5,
         inst2_stateArray_S33reg_gff_1_SFF_2_n5,
         inst2_stateArray_S33reg_gff_1_SFF_1_n5,
         inst2_stateArray_S33reg_gff_1_SFF_0_n5,
         inst2_stateArray_S32reg_gff_1_SFF_7_n5,
         inst2_stateArray_S32reg_gff_1_SFF_6_n5,
         inst2_stateArray_S32reg_gff_1_SFF_5_n5,
         inst2_stateArray_S32reg_gff_1_SFF_4_n6,
         inst2_stateArray_S32reg_gff_1_SFF_3_n6,
         inst2_stateArray_S32reg_gff_1_SFF_2_n6,
         inst2_stateArray_S32reg_gff_1_SFF_1_n6,
         inst2_stateArray_S32reg_gff_1_SFF_0_n6,
         inst2_stateArray_S31reg_gff_1_SFF_7_n6,
         inst2_stateArray_S31reg_gff_1_SFF_6_n6,
         inst2_stateArray_S31reg_gff_1_SFF_5_n6,
         inst2_stateArray_S31reg_gff_1_SFF_4_n6,
         inst2_stateArray_S31reg_gff_1_SFF_3_n6,
         inst2_stateArray_S31reg_gff_1_SFF_2_n6,
         inst2_stateArray_S31reg_gff_1_SFF_1_n6,
         inst2_stateArray_S31reg_gff_1_SFF_0_n6,
         inst2_stateArray_S30reg_gff_1_SFF_7_n5,
         inst2_stateArray_S30reg_gff_1_SFF_6_n5,
         inst2_stateArray_S30reg_gff_1_SFF_5_n5,
         inst2_stateArray_S30reg_gff_1_SFF_4_n5,
         inst2_stateArray_S30reg_gff_1_SFF_3_n5,
         inst2_stateArray_S30reg_gff_1_SFF_2_n5,
         inst2_stateArray_S30reg_gff_1_SFF_1_n5,
         inst2_stateArray_S30reg_gff_1_SFF_0_n5,
         inst2_stateArray_S23reg_gff_1_SFF_7_n5,
         inst2_stateArray_S23reg_gff_1_SFF_6_n5,
         inst2_stateArray_S23reg_gff_1_SFF_5_n5,
         inst2_stateArray_S23reg_gff_1_SFF_4_n6,
         inst2_stateArray_S23reg_gff_1_SFF_3_n6,
         inst2_stateArray_S23reg_gff_1_SFF_2_n6,
         inst2_stateArray_S23reg_gff_1_SFF_1_n6,
         inst2_stateArray_S23reg_gff_1_SFF_0_n6,
         inst2_stateArray_S22reg_gff_1_SFF_7_n6,
         inst2_stateArray_S22reg_gff_1_SFF_6_n6,
         inst2_stateArray_S22reg_gff_1_SFF_5_n6,
         inst2_stateArray_S22reg_gff_1_SFF_4_n6,
         inst2_stateArray_S22reg_gff_1_SFF_3_n6,
         inst2_stateArray_S22reg_gff_1_SFF_2_n6,
         inst2_stateArray_S22reg_gff_1_SFF_1_n6,
         inst2_stateArray_S22reg_gff_1_SFF_0_n6,
         inst2_stateArray_S21reg_gff_1_SFF_7_n6,
         inst2_stateArray_S21reg_gff_1_SFF_6_n6,
         inst2_stateArray_S21reg_gff_1_SFF_5_n6,
         inst2_stateArray_S21reg_gff_1_SFF_4_n6,
         inst2_stateArray_S21reg_gff_1_SFF_3_n6,
         inst2_stateArray_S21reg_gff_1_SFF_2_n6,
         inst2_stateArray_S21reg_gff_1_SFF_1_n6,
         inst2_stateArray_S21reg_gff_1_SFF_0_n6,
         inst2_stateArray_S20reg_gff_1_SFF_7_n5,
         inst2_stateArray_S20reg_gff_1_SFF_6_n5,
         inst2_stateArray_S20reg_gff_1_SFF_5_n5,
         inst2_stateArray_S20reg_gff_1_SFF_4_n5,
         inst2_stateArray_S20reg_gff_1_SFF_3_n5,
         inst2_stateArray_S20reg_gff_1_SFF_2_n5,
         inst2_stateArray_S20reg_gff_1_SFF_1_n5,
         inst2_stateArray_S20reg_gff_1_SFF_0_n5,
         inst2_stateArray_S13reg_gff_1_SFF_7_n5,
         inst2_stateArray_S13reg_gff_1_SFF_6_n5,
         inst2_stateArray_S13reg_gff_1_SFF_5_n5,
         inst2_stateArray_S13reg_gff_1_SFF_4_n6,
         inst2_stateArray_S13reg_gff_1_SFF_3_n6,
         inst2_stateArray_S13reg_gff_1_SFF_2_n6,
         inst2_stateArray_S13reg_gff_1_SFF_1_n6,
         inst2_stateArray_S13reg_gff_1_SFF_0_n6,
         inst2_stateArray_S12reg_gff_1_SFF_7_n6,
         inst2_stateArray_S12reg_gff_1_SFF_6_n6,
         inst2_stateArray_S12reg_gff_1_SFF_5_n6,
         inst2_stateArray_S12reg_gff_1_SFF_4_n6,
         inst2_stateArray_S12reg_gff_1_SFF_3_n6,
         inst2_stateArray_S12reg_gff_1_SFF_2_n6,
         inst2_stateArray_S12reg_gff_1_SFF_1_n6,
         inst2_stateArray_S12reg_gff_1_SFF_0_n6,
         inst2_stateArray_S11reg_gff_1_SFF_7_n6,
         inst2_stateArray_S11reg_gff_1_SFF_6_n6,
         inst2_stateArray_S11reg_gff_1_SFF_5_n6,
         inst2_stateArray_S11reg_gff_1_SFF_4_n6,
         inst2_stateArray_S11reg_gff_1_SFF_3_n6,
         inst2_stateArray_S11reg_gff_1_SFF_2_n6,
         inst2_stateArray_S11reg_gff_1_SFF_1_n6,
         inst2_stateArray_S11reg_gff_1_SFF_0_n6,
         inst2_stateArray_S10reg_gff_1_SFF_7_n5,
         inst2_stateArray_S10reg_gff_1_SFF_6_n5,
         inst2_stateArray_S10reg_gff_1_SFF_5_n5,
         inst2_stateArray_S10reg_gff_1_SFF_4_n5,
         inst2_stateArray_S10reg_gff_1_SFF_3_n5,
         inst2_stateArray_S10reg_gff_1_SFF_2_n5,
         inst2_stateArray_S10reg_gff_1_SFF_1_n5,
         inst2_stateArray_S10reg_gff_1_SFF_0_n5,
         inst2_stateArray_S03reg_gff_1_SFF_7_n5,
         inst2_stateArray_S03reg_gff_1_SFF_6_n5,
         inst2_stateArray_S03reg_gff_1_SFF_5_n5,
         inst2_stateArray_S03reg_gff_1_SFF_4_n6,
         inst2_stateArray_S03reg_gff_1_SFF_3_n6,
         inst2_stateArray_S03reg_gff_1_SFF_2_n6,
         inst2_stateArray_S03reg_gff_1_SFF_1_n6,
         inst2_stateArray_S03reg_gff_1_SFF_0_n6,
         inst2_stateArray_S02reg_gff_1_SFF_7_n6,
         inst2_stateArray_S02reg_gff_1_SFF_6_n6,
         inst2_stateArray_S02reg_gff_1_SFF_5_n6,
         inst2_stateArray_S02reg_gff_1_SFF_4_n6,
         inst2_stateArray_S02reg_gff_1_SFF_3_n6,
         inst2_stateArray_S02reg_gff_1_SFF_2_n6,
         inst2_stateArray_S02reg_gff_1_SFF_1_n6,
         inst2_stateArray_S02reg_gff_1_SFF_0_n6,
         inst2_stateArray_S01reg_gff_1_SFF_7_n6,
         inst2_stateArray_S01reg_gff_1_SFF_6_n6,
         inst2_stateArray_S01reg_gff_1_SFF_5_n6,
         inst2_stateArray_S01reg_gff_1_SFF_4_n6,
         inst2_stateArray_S01reg_gff_1_SFF_3_n6,
         inst2_stateArray_S01reg_gff_1_SFF_2_n6,
         inst2_stateArray_S01reg_gff_1_SFF_1_n6,
         inst2_stateArray_S01reg_gff_1_SFF_0_n6,
         inst2_stateArray_S00reg_gff_1_SFF_7_n6,
         inst2_stateArray_S00reg_gff_1_SFF_6_n6,
         inst2_stateArray_S00reg_gff_1_SFF_5_n6,
         inst2_stateArray_S00reg_gff_1_SFF_4_n6,
         inst2_stateArray_S00reg_gff_1_SFF_3_n6,
         inst2_stateArray_S00reg_gff_1_SFF_2_n6,
         inst2_stateArray_S00reg_gff_1_SFF_1_n6,
         inst2_stateArray_S00reg_gff_1_SFF_0_n6, inst2_ctrl_seq4_SFF_1_n5,
         inst2_ctrl_seq4_SFF_0_n5, inst2_ctrl_seq6_SFF_4_n5,
         inst2_ctrl_seq6_SFF_3_n5, inst2_ctrl_seq6_SFF_2_n5,
         inst2_ctrl_seq6_SFF_1_n5, inst2_ctrl_seq6_SFF_0_n5, inst2_ctrl_n6,
         inst3_n2873, inst3_n2872, inst3_n2871, inst3_n2870, inst3_n2869,
         inst3_n2868, inst3_n2867, inst3_n2866, inst3_n2865, inst3_n2864,
         inst3_n2863, inst3_n2862, inst3_n2861, inst3_n2860, inst3_n2859,
         inst3_n2858, inst3_n2857, inst3_n2856, inst3_n2855, inst3_n2854,
         inst3_n2853, inst3_n2852, inst3_n2851, inst3_n2850, inst3_n2849,
         inst3_n2848, inst3_n2847, inst3_n2846, inst3_n2845, inst3_n2844,
         inst3_n2843, inst3_n2842, inst3_n2841, inst3_n2840, inst3_n2839,
         inst3_n2838, inst3_n2837, inst3_n2836, inst3_n2835, inst3_n2834,
         inst3_n2833, inst3_n2832, inst3_n2831, inst3_n2830, inst3_n2829,
         inst3_n2828, inst3_n2827, inst3_n2826, inst3_n2825, inst3_n2824,
         inst3_n2823, inst3_n2822, inst3_n2821, inst3_n2820, inst3_n2819,
         inst3_n2818, inst3_n2817, inst3_n2816, inst3_n2815, inst3_n2814,
         inst3_n2813, inst3_n2812, inst3_n2811, inst3_n2810, inst3_n2809,
         inst3_n2808, inst3_n2807, inst3_n2806, inst3_n2805, inst3_n2804,
         inst3_n2803, inst3_n2802, inst3_n2801, inst3_n2800, inst3_n2799,
         inst3_n2798, inst3_n2797, inst3_n2796, inst3_n2795, inst3_n2794,
         inst3_n2793, inst3_n2792, inst3_n2791, inst3_n2790, inst3_n2789,
         inst3_n2788, inst3_n2787, inst3_n2786, inst3_n2785, inst3_n2784,
         inst3_n2783, inst3_n2782, inst3_n2781, inst3_n2780, inst3_n2779,
         inst3_n2778, inst3_n2777, inst3_n2776, inst3_n2775, inst3_n2774,
         inst3_n2773, inst3_n2772, inst3_n2771, inst3_n2770, inst3_n2769,
         inst3_n2768, inst3_n2767, inst3_n2766, inst3_n2765, inst3_n2764,
         inst3_n2763, inst3_n2762, inst3_n2761, inst3_n2760, inst3_n2759,
         inst3_n2758, inst3_n2757, inst3_n2756, inst3_n2755, inst3_n2754,
         inst3_n2753, inst3_n2752, inst3_n2751, inst3_n2750, inst3_n2749,
         inst3_n2748, inst3_n2747, inst3_n2746, inst3_n2745, inst3_n2744,
         inst3_n2743, inst3_n2742, inst3_n2741, inst3_n2740, inst3_n2739,
         inst3_n2738, inst3_n2737, inst3_n2736, inst3_n2735, inst3_n2734,
         inst3_n2733, inst3_n2732, inst3_n2731, inst3_n2730, inst3_n2729,
         inst3_n2728, inst3_n2727, inst3_n2726, inst3_n2725, inst3_n2724,
         inst3_n2723, inst3_n2722, inst3_n2721, inst3_n2720, inst3_n2719,
         inst3_n2718, inst3_n2717, inst3_n2716, inst3_n2715, inst3_n2714,
         inst3_n2713, inst3_n2712, inst3_n2711, inst3_n2710, inst3_n2709,
         inst3_n2708, inst3_n2707, inst3_n2706, inst3_n2705, inst3_n2704,
         inst3_n2703, inst3_n2702, inst3_n2701, inst3_n2700, inst3_n2699,
         inst3_n2698, inst3_n2697, inst3_n2696, inst3_n2695, inst3_n2694,
         inst3_n2693, inst3_n2692, inst3_n2691, inst3_n2690, inst3_n2689,
         inst3_n2688, inst3_n2687, inst3_n2686, inst3_n2685, inst3_n2684,
         inst3_n2683, inst3_n2682, inst3_n2681, inst3_n2680, inst3_n2679,
         inst3_n2678, inst3_n2677, inst3_n2676, inst3_n2675, inst3_n2674,
         inst3_n2673, inst3_n2672, inst3_n2671, inst3_n2670, inst3_n2669,
         inst3_n2668, inst3_n2667, inst3_n2666, inst3_n2665, inst3_n2664,
         inst3_n2663, inst3_n2662, inst3_n2661, inst3_n2660, inst3_n2659,
         inst3_n2658, inst3_n2657, inst3_n2656, inst3_n2655, inst3_n2654,
         inst3_n2653, inst3_n2652, inst3_n2651, inst3_n2650, inst3_n2649,
         inst3_n2648, inst3_n2647, inst3_n2646, inst3_n2645, inst3_n2644,
         inst3_n2643, inst3_n2642, inst3_n2641, inst3_n2640, inst3_n2639,
         inst3_n2638, inst3_n2637, inst3_n2636, inst3_n2635, inst3_n2634,
         inst3_n2633, inst3_n2632, inst3_n2631, inst3_n2630, inst3_n2629,
         inst3_n2628, inst3_n2627, inst3_n2626, inst3_n2625, inst3_n2624,
         inst3_n2623, inst3_n2622, inst3_n2621, inst3_n2620, inst3_n2619,
         inst3_n2618, inst3_n2617, inst3_n2616, inst3_n2615, inst3_n2614,
         inst3_n2613, inst3_n2612, inst3_n2611, inst3_n2610, inst3_n2609,
         inst3_n2608, inst3_n2607, inst3_n2606, inst3_n2605, inst3_n2604,
         inst3_n2603, inst3_n2602, inst3_n2601, inst3_n2600, inst3_n2599,
         inst3_n2598, inst3_n2597, inst3_n2596, inst3_n2595, inst3_n2594,
         inst3_n2593, inst3_n2592, inst3_n2591, inst3_n2590, inst3_n2589,
         inst3_n2588, inst3_n2587, inst3_n2586, inst3_n2585, inst3_n2584,
         inst3_n2583, inst3_n2582, inst3_n2581, inst3_n2580, inst3_n2579,
         inst3_n2578, inst3_n2577, inst3_n2576, inst3_n2575, inst3_n2574,
         inst3_n2573, inst3_n2572, inst3_n2571, inst3_n2570, inst3_n2569,
         inst3_n2568, inst3_n2567, inst3_n2566, inst3_n2565, inst3_n2564,
         inst3_n2563, inst3_n2562, inst3_n2561, inst3_n2560, inst3_n2559,
         inst3_n2558, inst3_n2557, inst3_n2556, inst3_n2555, inst3_n2554,
         inst3_n2553, inst3_n2552, inst3_n2551, inst3_n2550, inst3_n2549,
         inst3_n2548, inst3_n2547, inst3_n2546, inst3_n2545, inst3_n2544,
         inst3_n2543, inst3_n2542, inst3_n2541, inst3_n2540, inst3_n2539,
         inst3_n2538, inst3_n2537, inst3_n2536, inst3_n2535, inst3_n2534,
         inst3_n2533, inst3_n2532, inst3_n2531, inst3_n2530, inst3_n2529,
         inst3_n2528, inst3_n2527, inst3_n2526, inst3_n2525, inst3_n2524,
         inst3_n2523, inst3_n2522, inst3_n2521, inst3_n2520, inst3_n2519,
         inst3_n2518, inst3_n2517, inst3_n2516, inst3_n2515, inst3_n2514,
         inst3_n2513, inst3_n2512, inst3_n2511, inst3_n2510, inst3_n2509,
         inst3_n2508, inst3_n2507, inst3_n2506, inst3_n2505, inst3_n2504,
         inst3_n2503, inst3_n2502, inst3_n2501, inst3_n2500, inst3_n2499,
         inst3_n2498, inst3_n2497, inst3_n2496, inst3_n2495, inst3_n2494,
         inst3_n2493, inst3_n2492, inst3_n2491, inst3_n2490, inst3_n2489,
         inst3_n2488, inst3_n2487, inst3_n2486, inst3_n2485, inst3_n2484,
         inst3_n2483, inst3_n2482, inst3_n2481, inst3_n2480, inst3_n2479,
         inst3_n2478, inst3_n2477, inst3_n2476, inst3_n2475, inst3_n2474,
         inst3_n2473, inst3_n2472, inst3_n2471, inst3_n2470, inst3_n2469,
         inst3_n2468, inst3_n2467, inst3_n2466, inst3_n2465, inst3_n2464,
         inst3_n2463, inst3_n2462, inst3_n2461, inst3_n2460, inst3_n2459,
         inst3_n2458, inst3_n2457, inst3_n2456, inst3_n2455, inst3_n2454,
         inst3_n2453, inst3_n2452, inst3_n2451, inst3_n2450, inst3_n2449,
         inst3_n2448, inst3_n2447, inst3_n2446, inst3_n2445, inst3_n2444,
         inst3_n2443, inst3_n2442, inst3_n2441, inst3_n2440, inst3_n2439,
         inst3_n2438, inst3_n2437, inst3_n2436, inst3_n2435, inst3_n2434,
         inst3_n2433, inst3_n2432, inst3_n2431, inst3_n2430, inst3_n2429,
         inst3_n2428, inst3_n2427, inst3_n2426, inst3_n2425, inst3_n2424,
         inst3_n2423, inst3_n2422, inst3_n2421, inst3_n2420, inst3_n2419,
         inst3_n2418, inst3_n2417, inst3_n2416, inst3_n2415, inst3_n2414,
         inst3_n2413, inst3_n2412, inst3_n2411, inst3_n2410, inst3_n2409,
         inst3_n2408, inst3_n2407, inst3_n2406, inst3_n2405, inst3_n2404,
         inst3_n2403, inst3_n2402, inst3_n2401, inst3_n2400, inst3_n2399,
         inst3_n2398, inst3_n2397, inst3_n2396, inst3_n2395, inst3_n2394,
         inst3_n2393, inst3_n2392, inst3_n2391, inst3_n2390, inst3_n2389,
         inst3_n2388, inst3_n2387, inst3_n2386, inst3_n2385, inst3_n2384,
         inst3_n2383, inst3_n2382, inst3_n2381, inst3_n2380, inst3_n2379,
         inst3_n2378, inst3_n2377, inst3_n2376, inst3_n2375, inst3_n2374,
         inst3_n2373, inst3_n2372, inst3_n2371, inst3_n2370, inst3_n2369,
         inst3_n2368, inst3_n2367, inst3_n2366, inst3_n2365, inst3_n2364,
         inst3_n2363, inst3_n2362, inst3_n2361, inst3_n2360, inst3_n2359,
         inst3_n2358, inst3_n2357, inst3_n2356, inst3_n2355, inst3_n2354,
         inst3_n2353, inst3_n2352, inst3_n2351, inst3_n2350, inst3_n2349,
         inst3_n2348, inst3_n2347, inst3_n2346, inst3_n2345, inst3_n2344,
         inst3_n2343, inst3_n2342, inst3_n2341, inst3_n2340, inst3_n2339,
         inst3_n2338, inst3_n2337, inst3_n2336, inst3_n2335, inst3_n2334,
         inst3_n2333, inst3_n2332, inst3_n2331, inst3_n2330, inst3_n2329,
         inst3_n2328, inst3_n2327, inst3_n2326, inst3_n2325, inst3_n2324,
         inst3_n2323, inst3_n2322, inst3_n2321, inst3_n2320, inst3_n2319,
         inst3_n2318, inst3_n2317, inst3_n2316, inst3_n2315, inst3_n2314,
         inst3_n2313, inst3_n2312, inst3_n2311, inst3_n2310, inst3_n2309,
         inst3_n2308, inst3_n2307, inst3_n2306, inst3_n2305, inst3_n2304,
         inst3_n2303, inst3_n2302, inst3_n2301, inst3_n2300, inst3_n2299,
         inst3_n2298, inst3_n2297, inst3_n2296, inst3_n2295, inst3_n2294,
         inst3_n2293, inst3_n2292, inst3_n2291, inst3_n2290, inst3_n2289,
         inst3_n2288, inst3_n2287, inst3_n2286, inst3_n2285, inst3_n2284,
         inst3_n2283, inst3_n2282, inst3_n2281, inst3_n2280, inst3_n2279,
         inst3_n2278, inst3_n2277, inst3_n2276, inst3_n2275, inst3_n2274,
         inst3_n2273, inst3_n2272, inst3_n2271, inst3_n2270, inst3_n2269,
         inst3_n2268, inst3_n2267, inst3_n2266, inst3_n2265, inst3_n2264,
         inst3_n2263, inst3_n2262, inst3_n2261, inst3_n2260, inst3_n2259,
         inst3_n2258, inst3_n2257, inst3_n2256, inst3_n2255, inst3_n2254,
         inst3_n2253, inst3_n2252, inst3_n2251, inst3_n2250, inst3_n2249,
         inst3_n2248, inst3_n2247, inst3_n2246, inst3_n2245, inst3_n2244,
         inst3_n2243, inst3_n2242, inst3_n2241, inst3_n2240, inst3_n2239,
         inst3_n2238, inst3_n2237, inst3_n2236, inst3_n2235, inst3_n2234,
         inst3_n2233, inst3_n2232, inst3_n2231, inst3_n2230, inst3_n2229,
         inst3_n2228, inst3_n2227, inst3_n2226, inst3_n2225, inst3_n2224,
         inst3_n2223, inst3_n2222, inst3_n2221, inst3_n2220, inst3_n2219,
         inst3_n2218, inst3_n2217, inst3_n2216, inst3_n2215, inst3_n2214,
         inst3_n2213, inst3_n2212, inst3_n2211, inst3_n2210, inst3_n2209,
         inst3_n2208, inst3_n2207, inst3_n2206, inst3_n2205, inst3_n2204,
         inst3_n2203, inst3_n2202, inst3_n2201, inst3_n2200, inst3_n2199,
         inst3_n2198, inst3_n2197, inst3_n2196, inst3_n2195, inst3_n2194,
         inst3_n2193, inst3_n2192, inst3_n2191, inst3_n2190, inst3_n2189,
         inst3_n2188, inst3_n2187, inst3_n2186, inst3_n2185, inst3_n2184,
         inst3_n2183, inst3_n2182, inst3_n2181, inst3_n2180, inst3_n2179,
         inst3_n2178, inst3_n2177, inst3_n2176, inst3_n2175, inst3_n2174,
         inst3_n2173, inst3_n2172, inst3_n2171, inst3_n2170, inst3_n2169,
         inst3_n2168, inst3_n2167, inst3_n2166, inst3_n2165, inst3_n2164,
         inst3_n2163, inst3_n2162, inst3_n2161, inst3_n2160, inst3_n2159,
         inst3_n2158, inst3_n2157, inst3_n2156, inst3_n2155, inst3_n2154,
         inst3_n2153, inst3_n2152, inst3_n2151, inst3_n2150, inst3_n2149,
         inst3_n2148, inst3_n2147, inst3_n2146, inst3_n2145, inst3_n2144,
         inst3_n2143, inst3_n2142, inst3_n2141, inst3_n2140, inst3_n2139,
         inst3_n2138, inst3_n2137, inst3_n2136, inst3_n2135, inst3_n2134,
         inst3_n2133, inst3_n2132, inst3_n2131, inst3_n2130, inst3_n2129,
         inst3_n2128, inst3_n2127, inst3_n2126, inst3_n2125, inst3_n2124,
         inst3_n2123, inst3_n2122, inst3_n2121, inst3_n2120, inst3_n2119,
         inst3_n2118, inst3_n2117, inst3_n2116, inst3_n2115, inst3_n2114,
         inst3_n2113, inst3_n2112, inst3_n2111, inst3_n2110, inst3_n2109,
         inst3_n2108, inst3_n2107, inst3_n2106, inst3_n2105, inst3_n2104,
         inst3_n2103, inst3_n2102, inst3_n2101, inst3_n2100, inst3_n2099,
         inst3_n2098, inst3_n2097, inst3_n2096, inst3_n2095, inst3_n2094,
         inst3_n2093, inst3_n2092, inst3_n2091, inst3_n2090, inst3_n2089,
         inst3_n2088, inst3_n2087, inst3_n2086, inst3_n2085, inst3_n2084,
         inst3_n2083, inst3_n2082, inst3_n2081, inst3_n2080, inst3_n2079,
         inst3_n2078, inst3_n2077, inst3_n2076, inst3_n2075, inst3_n2074,
         inst3_n2073, inst3_n2072, inst3_n2071, inst3_n2070, inst3_n2069,
         inst3_n2068, inst3_n2067, inst3_n2066, inst3_n2065, inst3_n2064,
         inst3_n2063, inst3_n2062, inst3_n2061, inst3_n2060, inst3_n2059,
         inst3_n2058, inst3_n2057, inst3_n2056, inst3_n2055, inst3_n2054,
         inst3_n2053, inst3_n2052, inst3_n2051, inst3_n2050, inst3_n2049,
         inst3_n2048, inst3_n2047, inst3_n2046, inst3_n2045, inst3_n2044,
         inst3_n2043, inst3_n2042, inst3_n2041, inst3_n2040, inst3_n2039,
         inst3_n2038, inst3_n2037, inst3_n2036, inst3_n2035, inst3_n2034,
         inst3_n2033, inst3_n2032, inst3_n2031, inst3_n2030, inst3_n2029,
         inst3_n2028, inst3_n2027, inst3_n2026, inst3_n2025, inst3_n2024,
         inst3_n2023, inst3_n2022, inst3_n2021, inst3_n2020, inst3_n2019,
         inst3_n2018, inst3_n2017, inst3_n2016, inst3_n2015, inst3_n2014,
         inst3_n2013, inst3_n2012, inst3_n2011, inst3_n2010, inst3_n2009,
         inst3_n2008, inst3_n2007, inst3_n2006, inst3_n2005, inst3_n2004,
         inst3_n2003, inst3_n2002, inst3_n2001, inst3_n2000, inst3_n1999,
         inst3_n1998, inst3_n1997, inst3_n1996, inst3_n1995, inst3_n1994,
         inst3_n1993, inst3_n1992, inst3_n1991, inst3_n1990, inst3_n1989,
         inst3_n1988, inst3_n1987, inst3_n1986, inst3_n1985, inst3_n1984,
         inst3_n1983, inst3_n1982, inst3_n1981, inst3_n1980, inst3_n1979,
         inst3_n1978, inst3_n1977, inst3_n1976, inst3_n1975, inst3_n1974,
         inst3_n1973, inst3_n1972, inst3_n1971, inst3_n1970, inst3_n1969,
         inst3_n1968, inst3_n1967, inst3_n1966, inst3_n1965, inst3_n1964,
         inst3_n1963, inst3_n1962, inst3_n1961, inst3_n1960, inst3_n1959,
         inst3_n1958, inst3_n1957, inst3_n1956, inst3_n1955, inst3_n1954,
         inst3_n1953, inst3_n1952, inst3_n1951, inst3_n1950, inst3_n1949,
         inst3_n1948, inst3_n1947, inst3_n1946, inst3_n1945, inst3_n1944,
         inst3_n1943, inst3_n1942, inst3_n1941, inst3_n1940, inst3_n1939,
         inst3_n1938, inst3_n1937, inst3_n1936, inst3_n1935, inst3_n1934,
         inst3_n1933, inst3_n1932, inst3_n1931, inst3_n1930, inst3_n1929,
         inst3_n1928, inst3_n1927, inst3_n1926, inst3_n1925, inst3_n1924,
         inst3_n1923, inst3_n1922, inst3_n1921, inst3_n1920, inst3_n1919,
         inst3_n1918, inst3_n1917, inst3_n1916, inst3_n1914, inst3_n1096,
         inst3_n1088, inst3_n1290, inst3_n1273, inst3_n1272, inst3_n1271,
         inst3_n1270, inst3_n1269, inst3_n1268, inst3_n1267, inst3_n1266,
         inst3_n1265, inst3_n1264, inst3_n1263, inst3_n1262, inst3_n1261,
         inst3_n1260, inst3_n1259, inst3_n1258, inst3_n1257, inst3_n1256,
         inst3_n1255, inst3_n1254, inst3_n1253, inst3_n1252, inst3_n1251,
         inst3_n1250, inst3_n1233, inst3_n1232, inst3_n1231, inst3_n1230,
         inst3_n1229, inst3_n1228, inst3_n1227, inst3_n1226, inst3_n1225,
         inst3_n1224, inst3_n1223, inst3_n1222, inst3_n1221, inst3_n1220,
         inst3_n1219, inst3_n1218, inst3_n1209, inst3_n1208, inst3_n1207,
         inst3_n1206, inst3_n1205, inst3_n1204, inst3_n1203, inst3_n1202,
         inst3_n1201, inst3_n1200, inst3_n1199, inst3_n1198, inst3_n1197,
         inst3_n1196, inst3_n1195, inst3_n1194, inst3_n1193, inst3_n1192,
         inst3_n1191, inst3_n1190, inst3_n1189, inst3_n1188, inst3_n1187,
         inst3_n1186, inst3_n1185, inst3_n1184, inst3_n1183, inst3_n1182,
         inst3_n1181, inst3_n1180, inst3_n1179, inst3_n1178, inst3_n1177,
         inst3_n1176, inst3_n1175, inst3_n1174, inst3_n1173, inst3_n1172,
         inst3_n1171, inst3_n1170, inst3_n1169, inst3_n1168, inst3_n1167,
         inst3_n1166, inst3_n1165, inst3_n1164, inst3_n1163, inst3_n1162,
         inst3_n1161, inst3_n1097, inst3_n1095, inst3_n1094, inst3_n1093,
         inst3_n1092, inst3_n1091, inst3_n1090, inst3_n1089, inst3_n1087,
         inst3_n1086, inst3_n1085, inst3_n1084, inst3_n1083, inst3_n1082,
         inst3_n1081, inst3_n1080, inst3_n1071, inst3_n718, inst3_n706,
         inst3_n581, inst3_n499, inst3_n444, inst3_n321, inst3_n233,
         inst3_n232, inst3_n231, inst3_n230, inst3_n228, inst3_n227,
         inst3_n226, inst3_n225, inst3_n224, inst3_n223, inst3_n222,
         inst3_n221, inst3_n220, inst3_n219, inst3_n218, inst3_n216,
         inst3_n215, inst3_n214, inst3_n212, inst3_n210, inst3_n209,
         inst3_n207, inst3_n206, inst3_n203, inst3_n202, inst3_n201,
         inst3_n199, inst3_n198, inst3_n197, inst3_n196, inst3_n194,
         inst3_n193, inst3_n191, inst3_n190, inst3_n143, inst3_n137,
         inst3_n136, inst3_n135, inst3_n134, inst3_n133, inst3_n132,
         inst3_n131, inst3_n130, inst3_n129, inst3_n128, inst3_n127,
         inst3_n126, inst3_n125, inst3_n124, inst3_n123, inst3_n122,
         inst3_n121, inst3_n120, inst3_n119, inst3_n118, inst3_n117,
         inst3_n116, inst3_n115, inst3_n114, inst3_n113, inst3_n112,
         inst3_n111, inst3_n110, inst3_n109, inst3_n108, inst3_n107, inst3_n98,
         inst3_n97, inst3_n96, inst3_n95, inst3_n94, inst3_n93, inst3_n92,
         inst3_n91, inst3_n90, inst3_n89, inst3_n88, inst3_n87, inst3_n86,
         inst3_n85, inst3_n84, inst3_n83, inst3_n82, inst3_n81, inst3_n80,
         inst3_n79, inst3_n78, inst3_n77, inst3_n76, inst3_n75, inst3_n74,
         inst3_n73, inst3_n72, inst3_n71, inst3_n70, inst3_n69, inst3_n68,
         inst3_n67, inst3_n65, inst3_n57, inst3_n25, inst3_n24, inst3_n22,
         inst3_n17, inst3_n14, inst3_n12, inst3_n11, inst3_n10, inst3_n9,
         inst3_n6, inst3_calcRCon_n44, inst3_calcRCon_n45, inst3_calcRCon_n46,
         inst3_calcRCon_n47, inst3_calcRCon_n48, inst3_calcRCon_n49,
         inst3_calcRCon_n50, inst3_calcRCon_n51,
         inst3_KeyArray_S33reg_gff_1_SFF_7_n5,
         inst3_KeyArray_S33reg_gff_1_SFF_6_n5,
         inst3_KeyArray_S33reg_gff_1_SFF_5_n5,
         inst3_KeyArray_S33reg_gff_1_SFF_4_n5,
         inst3_KeyArray_S33reg_gff_1_SFF_3_n5,
         inst3_KeyArray_S33reg_gff_1_SFF_2_n5,
         inst3_KeyArray_S33reg_gff_1_SFF_1_n5,
         inst3_KeyArray_S33reg_gff_1_SFF_0_n5,
         inst3_KeyArray_S32reg_gff_1_SFF_7_n5,
         inst3_KeyArray_S32reg_gff_1_SFF_6_n5,
         inst3_KeyArray_S32reg_gff_1_SFF_5_n5,
         inst3_KeyArray_S32reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S32reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S32reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S32reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S32reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S31reg_gff_1_SFF_7_n6,
         inst3_KeyArray_S31reg_gff_1_SFF_6_n6,
         inst3_KeyArray_S31reg_gff_1_SFF_5_n6,
         inst3_KeyArray_S31reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S31reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S31reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S31reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S31reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S30reg_gff_1_SFF_7_n6,
         inst3_KeyArray_S30reg_gff_1_SFF_6_n6,
         inst3_KeyArray_S30reg_gff_1_SFF_5_n6,
         inst3_KeyArray_S30reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S30reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S30reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S30reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S30reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S23reg_gff_1_SFF_7_n5,
         inst3_KeyArray_S23reg_gff_1_SFF_6_n5,
         inst3_KeyArray_S23reg_gff_1_SFF_5_n5,
         inst3_KeyArray_S23reg_gff_1_SFF_4_n5,
         inst3_KeyArray_S23reg_gff_1_SFF_3_n5,
         inst3_KeyArray_S23reg_gff_1_SFF_2_n5,
         inst3_KeyArray_S23reg_gff_1_SFF_1_n5,
         inst3_KeyArray_S23reg_gff_1_SFF_0_n5,
         inst3_KeyArray_S22reg_gff_1_SFF_7_n5,
         inst3_KeyArray_S22reg_gff_1_SFF_6_n5,
         inst3_KeyArray_S22reg_gff_1_SFF_5_n5,
         inst3_KeyArray_S22reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S22reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S22reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S22reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S22reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S21reg_gff_1_SFF_7_n6,
         inst3_KeyArray_S21reg_gff_1_SFF_6_n6,
         inst3_KeyArray_S21reg_gff_1_SFF_5_n6,
         inst3_KeyArray_S21reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S21reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S21reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S21reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S21reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S20reg_gff_1_SFF_7_n6,
         inst3_KeyArray_S20reg_gff_1_SFF_6_n6,
         inst3_KeyArray_S20reg_gff_1_SFF_5_n6,
         inst3_KeyArray_S20reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S20reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S20reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S20reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S20reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S13reg_gff_1_SFF_7_n5,
         inst3_KeyArray_S13reg_gff_1_SFF_6_n5,
         inst3_KeyArray_S13reg_gff_1_SFF_5_n5,
         inst3_KeyArray_S13reg_gff_1_SFF_4_n5,
         inst3_KeyArray_S13reg_gff_1_SFF_3_n5,
         inst3_KeyArray_S13reg_gff_1_SFF_2_n5,
         inst3_KeyArray_S13reg_gff_1_SFF_1_n5,
         inst3_KeyArray_S13reg_gff_1_SFF_0_n5,
         inst3_KeyArray_S12reg_gff_1_SFF_7_n5,
         inst3_KeyArray_S12reg_gff_1_SFF_6_n5,
         inst3_KeyArray_S12reg_gff_1_SFF_5_n5,
         inst3_KeyArray_S12reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S12reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S12reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S12reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S12reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S11reg_gff_1_SFF_7_n6,
         inst3_KeyArray_S11reg_gff_1_SFF_6_n6,
         inst3_KeyArray_S11reg_gff_1_SFF_5_n6,
         inst3_KeyArray_S11reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S11reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S11reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S11reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S11reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S10reg_gff_1_SFF_7_n6,
         inst3_KeyArray_S10reg_gff_1_SFF_6_n6,
         inst3_KeyArray_S10reg_gff_1_SFF_5_n6,
         inst3_KeyArray_S10reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S10reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S10reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S10reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S10reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S03reg_gff_1_SFF_7_n5,
         inst3_KeyArray_S03reg_gff_1_SFF_6_n5,
         inst3_KeyArray_S03reg_gff_1_SFF_5_n5,
         inst3_KeyArray_S03reg_gff_1_SFF_4_n5,
         inst3_KeyArray_S03reg_gff_1_SFF_3_n5,
         inst3_KeyArray_S03reg_gff_1_SFF_2_n5,
         inst3_KeyArray_S03reg_gff_1_SFF_1_n5,
         inst3_KeyArray_S03reg_gff_1_SFF_0_n5,
         inst3_KeyArray_S02reg_gff_1_SFF_7_n5,
         inst3_KeyArray_S02reg_gff_1_SFF_6_n5,
         inst3_KeyArray_S02reg_gff_1_SFF_5_n5,
         inst3_KeyArray_S02reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S02reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S02reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S02reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S02reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S01reg_gff_1_SFF_7_n6,
         inst3_KeyArray_S01reg_gff_1_SFF_6_n6,
         inst3_KeyArray_S01reg_gff_1_SFF_5_n6,
         inst3_KeyArray_S01reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S01reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S01reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S01reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S01reg_gff_1_SFF_0_n6,
         inst3_KeyArray_S00reg_gff_1_SFF_7_n6,
         inst3_KeyArray_S00reg_gff_1_SFF_6_n6,
         inst3_KeyArray_S00reg_gff_1_SFF_5_n6,
         inst3_KeyArray_S00reg_gff_1_SFF_4_n6,
         inst3_KeyArray_S00reg_gff_1_SFF_3_n6,
         inst3_KeyArray_S00reg_gff_1_SFF_2_n6,
         inst3_KeyArray_S00reg_gff_1_SFF_1_n6,
         inst3_KeyArray_S00reg_gff_1_SFF_0_n6,
         inst3_stateArray_S33reg_gff_1_SFF_7_n5,
         inst3_stateArray_S33reg_gff_1_SFF_6_n5,
         inst3_stateArray_S33reg_gff_1_SFF_5_n5,
         inst3_stateArray_S33reg_gff_1_SFF_4_n5,
         inst3_stateArray_S33reg_gff_1_SFF_3_n5,
         inst3_stateArray_S33reg_gff_1_SFF_2_n5,
         inst3_stateArray_S33reg_gff_1_SFF_1_n5,
         inst3_stateArray_S33reg_gff_1_SFF_0_n5,
         inst3_stateArray_S32reg_gff_1_SFF_7_n5,
         inst3_stateArray_S32reg_gff_1_SFF_6_n5,
         inst3_stateArray_S32reg_gff_1_SFF_5_n5,
         inst3_stateArray_S32reg_gff_1_SFF_4_n6,
         inst3_stateArray_S32reg_gff_1_SFF_3_n6,
         inst3_stateArray_S32reg_gff_1_SFF_2_n6,
         inst3_stateArray_S32reg_gff_1_SFF_1_n6,
         inst3_stateArray_S32reg_gff_1_SFF_0_n6,
         inst3_stateArray_S31reg_gff_1_SFF_7_n6,
         inst3_stateArray_S31reg_gff_1_SFF_6_n6,
         inst3_stateArray_S31reg_gff_1_SFF_5_n6,
         inst3_stateArray_S31reg_gff_1_SFF_4_n6,
         inst3_stateArray_S31reg_gff_1_SFF_3_n6,
         inst3_stateArray_S31reg_gff_1_SFF_2_n6,
         inst3_stateArray_S31reg_gff_1_SFF_1_n6,
         inst3_stateArray_S31reg_gff_1_SFF_0_n6,
         inst3_stateArray_S30reg_gff_1_SFF_7_n5,
         inst3_stateArray_S30reg_gff_1_SFF_6_n5,
         inst3_stateArray_S30reg_gff_1_SFF_5_n5,
         inst3_stateArray_S30reg_gff_1_SFF_4_n5,
         inst3_stateArray_S30reg_gff_1_SFF_3_n5,
         inst3_stateArray_S30reg_gff_1_SFF_2_n5,
         inst3_stateArray_S30reg_gff_1_SFF_1_n5,
         inst3_stateArray_S30reg_gff_1_SFF_0_n5,
         inst3_stateArray_S23reg_gff_1_SFF_7_n5,
         inst3_stateArray_S23reg_gff_1_SFF_6_n5,
         inst3_stateArray_S23reg_gff_1_SFF_5_n5,
         inst3_stateArray_S23reg_gff_1_SFF_4_n6,
         inst3_stateArray_S23reg_gff_1_SFF_3_n6,
         inst3_stateArray_S23reg_gff_1_SFF_2_n6,
         inst3_stateArray_S23reg_gff_1_SFF_1_n6,
         inst3_stateArray_S23reg_gff_1_SFF_0_n6,
         inst3_stateArray_S22reg_gff_1_SFF_7_n6,
         inst3_stateArray_S22reg_gff_1_SFF_6_n6,
         inst3_stateArray_S22reg_gff_1_SFF_5_n6,
         inst3_stateArray_S22reg_gff_1_SFF_4_n6,
         inst3_stateArray_S22reg_gff_1_SFF_3_n6,
         inst3_stateArray_S22reg_gff_1_SFF_2_n6,
         inst3_stateArray_S22reg_gff_1_SFF_1_n6,
         inst3_stateArray_S22reg_gff_1_SFF_0_n6,
         inst3_stateArray_S21reg_gff_1_SFF_7_n6,
         inst3_stateArray_S21reg_gff_1_SFF_6_n6,
         inst3_stateArray_S21reg_gff_1_SFF_5_n6,
         inst3_stateArray_S21reg_gff_1_SFF_4_n6,
         inst3_stateArray_S21reg_gff_1_SFF_3_n6,
         inst3_stateArray_S21reg_gff_1_SFF_2_n6,
         inst3_stateArray_S21reg_gff_1_SFF_1_n6,
         inst3_stateArray_S21reg_gff_1_SFF_0_n6,
         inst3_stateArray_S20reg_gff_1_SFF_7_n5,
         inst3_stateArray_S20reg_gff_1_SFF_6_n5,
         inst3_stateArray_S20reg_gff_1_SFF_5_n5,
         inst3_stateArray_S20reg_gff_1_SFF_4_n5,
         inst3_stateArray_S20reg_gff_1_SFF_3_n5,
         inst3_stateArray_S20reg_gff_1_SFF_2_n5,
         inst3_stateArray_S20reg_gff_1_SFF_1_n5,
         inst3_stateArray_S20reg_gff_1_SFF_0_n5,
         inst3_stateArray_S13reg_gff_1_SFF_7_n5,
         inst3_stateArray_S13reg_gff_1_SFF_6_n5,
         inst3_stateArray_S13reg_gff_1_SFF_5_n5,
         inst3_stateArray_S13reg_gff_1_SFF_4_n6,
         inst3_stateArray_S13reg_gff_1_SFF_3_n6,
         inst3_stateArray_S13reg_gff_1_SFF_2_n6,
         inst3_stateArray_S13reg_gff_1_SFF_1_n6,
         inst3_stateArray_S13reg_gff_1_SFF_0_n6,
         inst3_stateArray_S12reg_gff_1_SFF_7_n6,
         inst3_stateArray_S12reg_gff_1_SFF_6_n6,
         inst3_stateArray_S12reg_gff_1_SFF_5_n6,
         inst3_stateArray_S12reg_gff_1_SFF_4_n6,
         inst3_stateArray_S12reg_gff_1_SFF_3_n6,
         inst3_stateArray_S12reg_gff_1_SFF_2_n6,
         inst3_stateArray_S12reg_gff_1_SFF_1_n6,
         inst3_stateArray_S12reg_gff_1_SFF_0_n6,
         inst3_stateArray_S11reg_gff_1_SFF_7_n6,
         inst3_stateArray_S11reg_gff_1_SFF_6_n6,
         inst3_stateArray_S11reg_gff_1_SFF_5_n6,
         inst3_stateArray_S11reg_gff_1_SFF_4_n6,
         inst3_stateArray_S11reg_gff_1_SFF_3_n6,
         inst3_stateArray_S11reg_gff_1_SFF_2_n6,
         inst3_stateArray_S11reg_gff_1_SFF_1_n6,
         inst3_stateArray_S11reg_gff_1_SFF_0_n6,
         inst3_stateArray_S10reg_gff_1_SFF_7_n5,
         inst3_stateArray_S10reg_gff_1_SFF_6_n5,
         inst3_stateArray_S10reg_gff_1_SFF_5_n5,
         inst3_stateArray_S10reg_gff_1_SFF_4_n5,
         inst3_stateArray_S10reg_gff_1_SFF_3_n5,
         inst3_stateArray_S10reg_gff_1_SFF_2_n5,
         inst3_stateArray_S10reg_gff_1_SFF_1_n5,
         inst3_stateArray_S10reg_gff_1_SFF_0_n5,
         inst3_stateArray_S03reg_gff_1_SFF_7_n5,
         inst3_stateArray_S03reg_gff_1_SFF_6_n5,
         inst3_stateArray_S03reg_gff_1_SFF_5_n5,
         inst3_stateArray_S03reg_gff_1_SFF_4_n6,
         inst3_stateArray_S03reg_gff_1_SFF_3_n6,
         inst3_stateArray_S03reg_gff_1_SFF_2_n6,
         inst3_stateArray_S03reg_gff_1_SFF_1_n6,
         inst3_stateArray_S03reg_gff_1_SFF_0_n6,
         inst3_stateArray_S02reg_gff_1_SFF_7_n6,
         inst3_stateArray_S02reg_gff_1_SFF_6_n6,
         inst3_stateArray_S02reg_gff_1_SFF_5_n6,
         inst3_stateArray_S02reg_gff_1_SFF_4_n6,
         inst3_stateArray_S02reg_gff_1_SFF_3_n6,
         inst3_stateArray_S02reg_gff_1_SFF_2_n6,
         inst3_stateArray_S02reg_gff_1_SFF_1_n6,
         inst3_stateArray_S02reg_gff_1_SFF_0_n6,
         inst3_stateArray_S01reg_gff_1_SFF_7_n6,
         inst3_stateArray_S01reg_gff_1_SFF_6_n6,
         inst3_stateArray_S01reg_gff_1_SFF_5_n6,
         inst3_stateArray_S01reg_gff_1_SFF_4_n6,
         inst3_stateArray_S01reg_gff_1_SFF_3_n6,
         inst3_stateArray_S01reg_gff_1_SFF_2_n6,
         inst3_stateArray_S01reg_gff_1_SFF_1_n6,
         inst3_stateArray_S01reg_gff_1_SFF_0_n6,
         inst3_stateArray_S00reg_gff_1_SFF_7_n6,
         inst3_stateArray_S00reg_gff_1_SFF_6_n6,
         inst3_stateArray_S00reg_gff_1_SFF_5_n6,
         inst3_stateArray_S00reg_gff_1_SFF_4_n6,
         inst3_stateArray_S00reg_gff_1_SFF_3_n6,
         inst3_stateArray_S00reg_gff_1_SFF_2_n6,
         inst3_stateArray_S00reg_gff_1_SFF_1_n6,
         inst3_stateArray_S00reg_gff_1_SFF_0_n6, inst3_ctrl_seq4_SFF_1_n5,
         inst3_ctrl_seq4_SFF_0_n5, inst3_ctrl_seq6_SFF_4_n5,
         inst3_ctrl_seq6_SFF_3_n5, inst3_ctrl_seq6_SFF_2_n5,
         inst3_ctrl_seq6_SFF_1_n5, inst3_ctrl_seq6_SFF_0_n5, inst3_ctrl_n6,
         mv_0_n256, mv_0_n255, mv_0_n254, mv_0_n253, mv_0_n252, mv_0_n251,
         mv_0_n250, mv_0_n249, mv_0_n248, mv_0_n247, mv_0_n246, mv_0_n245,
         mv_0_n244, mv_0_n243, mv_0_n242, mv_0_n241, mv_0_n240, mv_0_n239,
         mv_0_n238, mv_0_n237, mv_0_n236, mv_0_n235, mv_0_n234, mv_0_n233,
         mv_0_n232, mv_0_n231, mv_0_n230, mv_0_n229, mv_0_n228, mv_0_n227,
         mv_0_n226, mv_0_n225, mv_0_n224, mv_0_n223, mv_0_n222, mv_0_n221,
         mv_0_n220, mv_0_n219, mv_0_n218, mv_0_n217, mv_0_n216, mv_0_n215,
         mv_0_n214, mv_0_n213, mv_0_n212, mv_0_n211, mv_0_n210, mv_0_n209,
         mv_0_n208, mv_0_n207, mv_0_n206, mv_0_n205, mv_0_n204, mv_0_n203,
         mv_0_n202, mv_0_n201, mv_0_n200, mv_0_n199, mv_0_n198, mv_0_n197,
         mv_0_n196, mv_0_n195, mv_0_n194, mv_0_n193, mv_0_n192, mv_0_n191,
         mv_0_n190, mv_0_n189, mv_0_n188, mv_0_n187, mv_0_n186, mv_0_n185,
         mv_0_n184, mv_0_n183, mv_0_n182, mv_0_n181, mv_0_n180, mv_0_n179,
         mv_0_n178, mv_0_n177, mv_0_n176, mv_0_n175, mv_0_n174, mv_0_n173,
         mv_0_n172, mv_0_n171, mv_0_n170, mv_0_n169, mv_0_n168, mv_0_n167,
         mv_0_n166, mv_0_n165, mv_0_n164, mv_0_n163, mv_0_n162, mv_0_n161,
         mv_0_n160, mv_0_n159, mv_0_n158, mv_0_n157, mv_0_n156, mv_0_n155,
         mv_0_n154, mv_0_n153, mv_0_n152, mv_0_n151, mv_0_n150, mv_0_n149,
         mv_0_n148, mv_0_n147, mv_0_n146, mv_0_n145, mv_0_n144, mv_0_n143,
         mv_0_n142, mv_0_n141, mv_0_n140, mv_0_n139, mv_0_n138, mv_0_n137,
         mv_0_n136, mv_0_n135, mv_0_n134, mv_0_n133, mv_0_n132, mv_0_n131,
         mv_0_n130, mv_0_n129, mv_0_n128, mv_0_n127, mv_0_n126, mv_0_n125,
         mv_0_n124, mv_0_n123, mv_0_n122, mv_0_n121, mv_0_n120, mv_0_n119,
         mv_0_n118, mv_0_n117, mv_0_n116, mv_0_n115, mv_0_n114, mv_0_n113,
         mv_0_n112, mv_0_n111, mv_0_n110, mv_0_n109, mv_0_n108, mv_0_n107,
         mv_0_n106, mv_0_n105, mv_0_n104, mv_0_n103, mv_0_n102, mv_0_n101,
         mv_0_n100, mv_0_n99, mv_0_n98, mv_0_n97, mv_0_n96, mv_0_n95, mv_0_n94,
         mv_0_n93, mv_0_n92, mv_0_n91, mv_0_n90, mv_0_n89, mv_0_n88, mv_0_n87,
         mv_0_n86, mv_0_n85, mv_0_n84, mv_0_n83, mv_0_n82, mv_0_n81, mv_0_n80,
         mv_0_n79, mv_0_n78, mv_0_n77, mv_0_n76, mv_0_n75, mv_0_n74, mv_0_n73,
         mv_0_n72, mv_0_n71, mv_0_n70, mv_0_n69, mv_0_n68, mv_0_n67, mv_0_n66,
         mv_0_n65, mv_0_n64, mv_0_n63, mv_0_n62, mv_0_n61, mv_0_n60, mv_0_n59,
         mv_0_n58, mv_0_n57, mv_0_n56, mv_0_n55, mv_0_n54, mv_0_n53, mv_0_n52,
         mv_0_n51, mv_0_n50, mv_0_n49, mv_0_n48, mv_0_n47, mv_0_n46, mv_0_n45,
         mv_0_n44, mv_0_n43, mv_0_n42, mv_0_n41, mv_0_n40, mv_0_n39, mv_0_n38,
         mv_0_n37, mv_0_n36, mv_0_n35, mv_0_n34, mv_0_n33, mv_0_n32, mv_0_n31,
         mv_0_n30, mv_0_n29, mv_0_n28, mv_0_n27, mv_0_n26, mv_0_n25, mv_0_n24,
         mv_0_n23, mv_0_n22, mv_0_n21, mv_0_n20, mv_0_n19, mv_0_n18, mv_0_n17,
         mv_0_n16, mv_0_n15, mv_0_n14, mv_0_n13, mv_0_n12, mv_0_n11, mv_0_n10,
         mv_0_n9, mv_0_n8, mv_0_n7, mv_0_n6, mv_0_n5, mv_0_n4, mv_0_n3,
         mv_0_n2, mv_0_n1, mv_1_n2, mv_1_n1;
  wire   [127:0] ciphertext1;
  wire   [127:0] ciphertext2;
  wire   [127:0] ciphertext3;

  OAI21_X1 inst1_U1162 ( .B1(inst1_n1224), .B2(inst1_n1223), .A(inst1_n1222),
        .ZN(inst1_n1188) );
  NOR2_X1 inst1_U1161 ( .A1(inst1_n143), .A2(inst1_n1250), .ZN(inst1_n1224) );
  OAI211_X1 inst1_U1160 ( .C1(inst1_n1221), .C2(inst1_n1220), .A(inst1_n1219),
        .B(inst1_n1218), .ZN(inst1_stateArray_S23reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst1_U1159 ( .B1(inst1_n1217), .B2(ciphertext1[49]), .A(
        inst1_n1216), .ZN(inst1_n1218) );
  OAI22_X1 inst1_U1158 ( .A1(inst1_n1121), .A2(inst1_n1035), .B1(inst1_n1215),
        .B2(inst1_n1235), .ZN(inst1_n1216) );
  AOI22_X1 inst1_U1157 ( .A1(done1), .A2(ciphertext1[33]), .B1(plaintext1[33]),
        .B2(inst1_n1228), .ZN(inst1_n1219) );
  XNOR2_X1 inst1_U1156 ( .A(inst1_n1214), .B(inst1_n1213), .ZN(inst1_n1221) );
  AOI22_X1 inst1_U1155 ( .A1(inst1_n1121), .A2(inst1_n1212), .B1(inst1_n1211),
        .B2(ciphertext1[25]), .ZN(inst1_n1213) );
  XNOR2_X1 inst1_U1154 ( .A(inst1_n1210), .B(inst1_n1209), .ZN(inst1_n1214) );
  OAI211_X1 inst1_U1153 ( .C1(inst1_n1208), .C2(inst1_n1207), .A(inst1_n1206),
        .B(inst1_n1205), .ZN(inst1_stateArray_S23reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst1_U1152 ( .B1(inst1_n1217), .B2(ciphertext1[50]), .A(
        inst1_n1204), .ZN(inst1_n1205) );
  OAI22_X1 inst1_U1151 ( .A1(inst1_n1109), .A2(inst1_n1203), .B1(inst1_n1119),
        .B2(inst1_n1215), .ZN(inst1_n1204) );
  AOI22_X1 inst1_U1150 ( .A1(inst1_n677), .A2(ciphertext1[34]), .B1(
        plaintext1[34]), .B2(inst1_n1228), .ZN(inst1_n1206) );
  XNOR2_X1 inst1_U1149 ( .A(inst1_n1202), .B(inst1_n1201), .ZN(inst1_n1208) );
  AOI22_X1 inst1_U1148 ( .A1(inst1_n1200), .A2(ciphertext1[90]), .B1(
        inst1_n1118), .B2(inst1_n1199), .ZN(inst1_n1201) );
  NOR2_X1 inst1_U1147 ( .A1(inst1_n1198), .A2(inst1_n1236), .ZN(
        inst1_ctrl_seq4_SFF_1_n5) );
  NOR2_X1 inst1_U1146 ( .A1(inst1_n1080), .A2(inst1_n732), .ZN(
        inst1_ctrl_seq6_SFF_1_n5) );
  NOR2_X1 inst1_U1145 ( .A1(inst1_n1079), .A2(inst1_n830), .ZN(
        inst1_ctrl_seq6_SFF_3_n5) );
  OAI211_X1 inst1_U1144 ( .C1(inst1_n1220), .C2(inst1_n1197), .A(inst1_n1196),
        .B(inst1_n1195), .ZN(inst1_stateArray_S23reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst1_U1143 ( .B1(inst1_n1217), .B2(ciphertext1[52]), .A(
        inst1_n1194), .ZN(inst1_n1195) );
  OAI22_X1 inst1_U1142 ( .A1(inst1_n1105), .A2(inst1_n1203), .B1(inst1_n1215),
        .B2(inst1_n1234), .ZN(inst1_n1194) );
  AOI22_X1 inst1_U1141 ( .A1(inst1_n677), .A2(ciphertext1[36]), .B1(
        plaintext1[36]), .B2(inst1_n1228), .ZN(inst1_n1196) );
  XNOR2_X1 inst1_U1140 ( .A(inst1_n1193), .B(inst1_n1192), .ZN(inst1_n1197) );
  AOI22_X1 inst1_U1139 ( .A1(inst1_n1100), .A2(inst1_n1191), .B1(inst1_n1190),
        .B2(ciphertext1[92]), .ZN(inst1_n1192) );
  AOI22_X1 inst1_U1138 ( .A1(inst1_n1212), .A2(inst1_n1187), .B1(inst1_n1186),
        .B2(inst1_n1211), .ZN(inst1_n1193) );
  OAI22_X1 inst1_U1137 ( .A1(inst1_n1061), .A2(inst1_n1185), .B1(inst1_n1071),
        .B2(inst1_n1184), .ZN(inst1_calcRCon_n45) );
  OAI21_X1 inst1_U1136 ( .B1(inst1_n1074), .B2(inst1_n1184), .A(inst1_n1183),
        .ZN(inst1_calcRCon_n50) );
  OAI221_X1 inst1_U1135 ( .B1(inst1_n1070), .B2(inst1_n1075), .C1(inst1_n1226),
        .C2(inst1_n1264), .A(inst1_n1217), .ZN(inst1_n1183) );
  OAI22_X1 inst1_U1134 ( .A1(inst1_n1061), .A2(inst1_n1184), .B1(inst1_n1060),
        .B2(inst1_n1182), .ZN(inst1_calcRCon_n46) );
  OAI21_X1 inst1_U1133 ( .B1(inst1_n1060), .B2(inst1_n1184), .A(inst1_n1181),
        .ZN(inst1_calcRCon_n47) );
  OAI221_X1 inst1_U1132 ( .B1(inst1_n1072), .B2(inst1_n1070), .C1(inst1_n1240),
        .C2(inst1_n1226), .A(inst1_n1217), .ZN(inst1_n1181) );
  NAND2_X1 inst1_U1131 ( .A1(inst1_n6), .A2(inst1_n1182), .ZN(inst1_n1184) );
  OAI211_X1 inst1_U1130 ( .C1(inst1_n908), .C2(inst1_n1185), .A(inst1_n1180),
        .B(inst1_n1179), .ZN(inst1_stateArray_S20reg_gff_1_SFF_0_n5) );
  NAND2_X1 inst1_U1129 ( .A1(inst1_n191), .A2(ciphertext1[48]), .ZN(
        inst1_n1179) );
  AOI22_X1 inst1_U1128 ( .A1(ciphertext1[56]), .A2(inst1_n385), .B1(
        plaintext1[56]), .B2(inst1_n1228), .ZN(inst1_n1180) );
  OAI211_X1 inst1_U1127 ( .C1(inst1_n909), .C2(inst1_n1185), .A(inst1_n1178),
        .B(inst1_n1177), .ZN(inst1_stateArray_S20reg_gff_1_SFF_1_n5) );
  NAND2_X1 inst1_U1126 ( .A1(inst1_n191), .A2(ciphertext1[49]), .ZN(
        inst1_n1177) );
  AOI22_X1 inst1_U1125 ( .A1(ciphertext1[57]), .A2(inst1_n385), .B1(
        plaintext1[57]), .B2(inst1_n1228), .ZN(inst1_n1178) );
  OAI211_X1 inst1_U1124 ( .C1(inst1_n910), .C2(inst1_n1182), .A(inst1_n1176),
        .B(inst1_n1175), .ZN(inst1_stateArray_S20reg_gff_1_SFF_2_n5) );
  NAND2_X1 inst1_U1123 ( .A1(inst1_n191), .A2(ciphertext1[50]), .ZN(
        inst1_n1175) );
  AOI22_X1 inst1_U1122 ( .A1(inst1_n677), .A2(ciphertext1[58]), .B1(
        plaintext1[58]), .B2(inst1_n1228), .ZN(inst1_n1176) );
  OAI211_X1 inst1_U1121 ( .C1(inst1_n911), .C2(inst1_n1185), .A(inst1_n1174),
        .B(inst1_n1173), .ZN(inst1_stateArray_S20reg_gff_1_SFF_3_n5) );
  NAND2_X1 inst1_U1120 ( .A1(inst1_n191), .A2(ciphertext1[51]), .ZN(
        inst1_n1173) );
  AOI22_X1 inst1_U1119 ( .A1(inst1_n677), .A2(ciphertext1[59]), .B1(
        plaintext1[59]), .B2(inst1_n1228), .ZN(inst1_n1174) );
  OAI211_X1 inst1_U1118 ( .C1(inst1_n912), .C2(inst1_n1185), .A(inst1_n1172),
        .B(inst1_n1171), .ZN(inst1_stateArray_S20reg_gff_1_SFF_4_n5) );
  NAND2_X1 inst1_U1117 ( .A1(inst1_n191), .A2(ciphertext1[52]), .ZN(
        inst1_n1171) );
  AOI22_X1 inst1_U1116 ( .A1(ciphertext1[60]), .A2(done1), .B1(plaintext1[60]),
        .B2(inst1_n1228), .ZN(inst1_n1172) );
  OAI211_X1 inst1_U1115 ( .C1(inst1_n913), .C2(inst1_n1185), .A(inst1_n1170),
        .B(inst1_n1169), .ZN(inst1_stateArray_S20reg_gff_1_SFF_5_n5) );
  NAND2_X1 inst1_U1114 ( .A1(inst1_n191), .A2(ciphertext1[53]), .ZN(
        inst1_n1169) );
  AOI22_X1 inst1_U1113 ( .A1(ciphertext1[61]), .A2(inst1_n677), .B1(
        plaintext1[61]), .B2(inst1_n1228), .ZN(inst1_n1170) );
  OAI211_X1 inst1_U1112 ( .C1(inst1_n914), .C2(inst1_n1185), .A(inst1_n1168),
        .B(inst1_n1167), .ZN(inst1_stateArray_S20reg_gff_1_SFF_6_n5) );
  NAND2_X1 inst1_U1111 ( .A1(inst1_n191), .A2(ciphertext1[54]), .ZN(
        inst1_n1167) );
  AOI22_X1 inst1_U1110 ( .A1(ciphertext1[62]), .A2(done1), .B1(plaintext1[62]),
        .B2(inst1_n1228), .ZN(inst1_n1168) );
  OAI211_X1 inst1_U1109 ( .C1(inst1_n915), .C2(inst1_n1182), .A(inst1_n1166),
        .B(inst1_n1165), .ZN(inst1_stateArray_S20reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst1_U1108 ( .A1(inst1_n191), .A2(ciphertext1[55]), .ZN(
        inst1_n1165) );
  AOI22_X1 inst1_U1107 ( .A1(done1), .A2(ciphertext1[63]), .B1(plaintext1[63]),
        .B2(inst1_n1228), .ZN(inst1_n1166) );
  OAI211_X1 inst1_U1106 ( .C1(inst1_n908), .C2(inst1_n1198), .A(inst1_n1164),
        .B(inst1_n1163), .ZN(inst1_stateArray_S21reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst1_U1105 ( .A1(plaintext1[48]), .A2(inst1_n710), .ZN(inst1_n1163) );
  AOI22_X1 inst1_U1104 ( .A1(inst1_n677), .A2(ciphertext1[48]), .B1(
        inst1_n1217), .B2(ciphertext1[32]), .ZN(inst1_n1164) );
  OAI211_X1 inst1_U1103 ( .C1(inst1_n909), .C2(inst1_n1198), .A(inst1_n1162),
        .B(inst1_n1161), .ZN(inst1_stateArray_S21reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst1_U1102 ( .A1(plaintext1[49]), .A2(inst1_n830), .ZN(inst1_n1161) );
  AOI22_X1 inst1_U1101 ( .A1(done1), .A2(ciphertext1[49]), .B1(inst1_n1217),
        .B2(ciphertext1[33]), .ZN(inst1_n1162) );
  OAI211_X1 inst1_U1100 ( .C1(inst1_n910), .C2(inst1_n1198), .A(inst1_n1160),
        .B(inst1_n1159), .ZN(inst1_stateArray_S21reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst1_U1099 ( .A1(plaintext1[50]), .A2(inst1_n1156), .ZN(
        inst1_n1159) );
  AOI22_X1 inst1_U1098 ( .A1(inst1_n677), .A2(ciphertext1[50]), .B1(
        inst1_n1217), .B2(ciphertext1[34]), .ZN(inst1_n1160) );
  OAI211_X1 inst1_U1097 ( .C1(inst1_n911), .C2(inst1_n1198), .A(inst1_n1158),
        .B(inst1_n1157), .ZN(inst1_stateArray_S21reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst1_U1096 ( .A1(plaintext1[51]), .A2(inst1_n1156), .ZN(
        inst1_n1157) );
  AOI22_X1 inst1_U1095 ( .A1(done1), .A2(ciphertext1[51]), .B1(inst1_n1217),
        .B2(ciphertext1[35]), .ZN(inst1_n1158) );
  OAI211_X1 inst1_U1094 ( .C1(inst1_n912), .C2(inst1_n1198), .A(inst1_n1155),
        .B(inst1_n1154), .ZN(inst1_stateArray_S21reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst1_U1093 ( .A1(plaintext1[52]), .A2(inst1_n522), .ZN(inst1_n1154) );
  AOI22_X1 inst1_U1092 ( .A1(inst1_n677), .A2(ciphertext1[52]), .B1(
        inst1_n1217), .B2(ciphertext1[36]), .ZN(inst1_n1155) );
  OAI211_X1 inst1_U1091 ( .C1(inst1_n913), .C2(inst1_n1198), .A(inst1_n1153),
        .B(inst1_n1152), .ZN(inst1_stateArray_S21reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst1_U1090 ( .A1(plaintext1[53]), .A2(inst1_n1156), .ZN(
        inst1_n1152) );
  AOI22_X1 inst1_U1089 ( .A1(done1), .A2(ciphertext1[53]), .B1(inst1_n1217),
        .B2(ciphertext1[37]), .ZN(inst1_n1153) );
  OAI211_X1 inst1_U1088 ( .C1(inst1_n914), .C2(inst1_n1198), .A(inst1_n1151),
        .B(inst1_n1150), .ZN(inst1_stateArray_S21reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst1_U1087 ( .A1(plaintext1[54]), .A2(inst1_n596), .ZN(inst1_n1150) );
  AOI22_X1 inst1_U1086 ( .A1(inst1_n677), .A2(ciphertext1[54]), .B1(
        inst1_n1217), .B2(ciphertext1[38]), .ZN(inst1_n1151) );
  OAI211_X1 inst1_U1085 ( .C1(inst1_n915), .C2(inst1_n1198), .A(inst1_n1149),
        .B(inst1_n1148), .ZN(inst1_stateArray_S21reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst1_U1084 ( .A1(plaintext1[55]), .A2(inst1_n1156), .ZN(
        inst1_n1148) );
  AOI22_X1 inst1_U1083 ( .A1(done1), .A2(ciphertext1[55]), .B1(inst1_n1217),
        .B2(ciphertext1[39]), .ZN(inst1_n1149) );
  OAI21_X1 inst1_U1082 ( .B1(inst1_n920), .B2(inst1_n1198), .A(inst1_n1147),
        .ZN(inst1_stateArray_S22reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst1_U1081 ( .B1(plaintext1[44]), .B2(inst1_n830), .A(inst1_n1146),
        .ZN(inst1_n1147) );
  OAI22_X1 inst1_U1080 ( .A1(inst1_n912), .A2(inst1_n1145), .B1(inst1_n1185),
        .B2(inst1_n1234), .ZN(inst1_n1146) );
  OAI21_X1 inst1_U1079 ( .B1(inst1_n1198), .B2(inst1_n1258), .A(inst1_n1144),
        .ZN(inst1_stateArray_S30reg_gff_1_SFF_0_n5) );
  AOI21_X1 inst1_U1078 ( .B1(plaintext1[24]), .B2(inst1_n710), .A(inst1_n1143),
        .ZN(inst1_n1144) );
  OAI22_X1 inst1_U1077 ( .A1(inst1_n1113), .A2(inst1_n1142), .B1(inst1_n940),
        .B2(inst1_n1182), .ZN(inst1_n1143) );
  OAI21_X1 inst1_U1076 ( .B1(inst1_n1198), .B2(inst1_n1257), .A(inst1_n1141),
        .ZN(inst1_stateArray_S30reg_gff_1_SFF_1_n5) );
  AOI21_X1 inst1_U1075 ( .B1(plaintext1[25]), .B2(inst1_n494), .A(inst1_n1140),
        .ZN(inst1_n1141) );
  OAI22_X1 inst1_U1074 ( .A1(inst1_n1121), .A2(inst1_n1145), .B1(inst1_n941),
        .B2(inst1_n1182), .ZN(inst1_n1140) );
  OAI21_X1 inst1_U1073 ( .B1(inst1_n1198), .B2(inst1_n1256), .A(inst1_n1139),
        .ZN(inst1_stateArray_S30reg_gff_1_SFF_2_n5) );
  AOI21_X1 inst1_U1072 ( .B1(plaintext1[26]), .B2(inst1_n830), .A(inst1_n1138),
        .ZN(inst1_n1139) );
  OAI22_X1 inst1_U1071 ( .A1(inst1_n1109), .A2(inst1_n1142), .B1(inst1_n942),
        .B2(inst1_n1182), .ZN(inst1_n1138) );
  OAI21_X1 inst1_U1070 ( .B1(inst1_n1198), .B2(inst1_n1255), .A(inst1_n1137),
        .ZN(inst1_stateArray_S30reg_gff_1_SFF_3_n5) );
  AOI21_X1 inst1_U1069 ( .B1(plaintext1[27]), .B2(inst1_n507), .A(inst1_n1136),
        .ZN(inst1_n1137) );
  OAI22_X1 inst1_U1068 ( .A1(inst1_n943), .A2(inst1_n1185), .B1(inst1_n1135),
        .B2(inst1_n1231), .ZN(inst1_n1136) );
  OAI21_X1 inst1_U1067 ( .B1(inst1_n1198), .B2(inst1_n1254), .A(inst1_n1134),
        .ZN(inst1_stateArray_S30reg_gff_1_SFF_4_n5) );
  AOI21_X1 inst1_U1066 ( .B1(plaintext1[28]), .B2(inst1_n1133), .A(inst1_n1132), .ZN(inst1_n1134) );
  OAI22_X1 inst1_U1065 ( .A1(inst1_n1105), .A2(inst1_n1145), .B1(inst1_n944),
        .B2(inst1_n1182), .ZN(inst1_n1132) );
  OAI21_X1 inst1_U1064 ( .B1(inst1_n1198), .B2(inst1_n1253), .A(inst1_n1131),
        .ZN(inst1_stateArray_S30reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst1_U1063 ( .B1(plaintext1[29]), .B2(inst1_n507), .A(inst1_n1130),
        .ZN(inst1_n1131) );
  OAI22_X1 inst1_U1062 ( .A1(inst1_n945), .A2(inst1_n1185), .B1(inst1_n1135),
        .B2(inst1_n1229), .ZN(inst1_n1130) );
  OAI21_X1 inst1_U1061 ( .B1(inst1_n1198), .B2(inst1_n1251), .A(inst1_n1129),
        .ZN(inst1_stateArray_S30reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst1_U1060 ( .B1(plaintext1[30]), .B2(inst1_n732), .A(inst1_n1128),
        .ZN(inst1_n1129) );
  OAI22_X1 inst1_U1059 ( .A1(inst1_n1097), .A2(inst1_n1145), .B1(inst1_n946),
        .B2(inst1_n1182), .ZN(inst1_n1128) );
  OAI21_X1 inst1_U1058 ( .B1(inst1_n1198), .B2(inst1_n1252), .A(inst1_n1127),
        .ZN(inst1_stateArray_S30reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst1_U1057 ( .B1(plaintext1[31]), .B2(inst1_n899), .A(inst1_n1126),
        .ZN(inst1_n1127) );
  OAI22_X1 inst1_U1056 ( .A1(inst1_n947), .A2(inst1_n1185), .B1(inst1_n1135),
        .B2(inst1_n1230), .ZN(inst1_n1126) );
  OAI21_X1 inst1_U1055 ( .B1(inst1_n940), .B2(inst1_n1198), .A(inst1_n1125),
        .ZN(inst1_stateArray_S32reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst1_U1054 ( .B1(plaintext1[8]), .B2(inst1_n596), .A(inst1_n1124),
        .ZN(inst1_n1125) );
  OAI22_X1 inst1_U1053 ( .A1(inst1_n932), .A2(inst1_n1145), .B1(inst1_n1182),
        .B2(inst1_n1258), .ZN(inst1_n1124) );
  OAI21_X1 inst1_U1052 ( .B1(inst1_n941), .B2(inst1_n1198), .A(inst1_n1123),
        .ZN(inst1_stateArray_S32reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst1_U1051 ( .B1(plaintext1[9]), .B2(inst1_n732), .A(inst1_n1120),
        .ZN(inst1_n1123) );
  OAI22_X1 inst1_U1050 ( .A1(inst1_n933), .A2(inst1_n1145), .B1(inst1_n1182),
        .B2(inst1_n1257), .ZN(inst1_n1120) );
  OAI21_X1 inst1_U1049 ( .B1(inst1_n942), .B2(inst1_n1198), .A(inst1_n1117),
        .ZN(inst1_stateArray_S32reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst1_U1048 ( .B1(plaintext1[10]), .B2(inst1_n830), .A(inst1_n1112),
        .ZN(inst1_n1117) );
  OAI22_X1 inst1_U1047 ( .A1(inst1_n934), .A2(inst1_n1145), .B1(inst1_n1182),
        .B2(inst1_n1256), .ZN(inst1_n1112) );
  OAI21_X1 inst1_U1046 ( .B1(inst1_n943), .B2(inst1_n1198), .A(inst1_n1108),
        .ZN(inst1_stateArray_S32reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst1_U1045 ( .B1(plaintext1[11]), .B2(inst1_n522), .A(inst1_n1107),
        .ZN(inst1_n1108) );
  OAI22_X1 inst1_U1044 ( .A1(inst1_n935), .A2(inst1_n1145), .B1(inst1_n1185),
        .B2(inst1_n1255), .ZN(inst1_n1107) );
  OAI21_X1 inst1_U1043 ( .B1(inst1_n944), .B2(inst1_n1198), .A(inst1_n1104),
        .ZN(inst1_stateArray_S32reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst1_U1042 ( .B1(plaintext1[12]), .B2(inst1_n732), .A(inst1_n1101),
        .ZN(inst1_n1104) );
  OAI22_X1 inst1_U1041 ( .A1(inst1_n936), .A2(inst1_n1145), .B1(inst1_n1182),
        .B2(inst1_n1254), .ZN(inst1_n1101) );
  OAI21_X1 inst1_U1040 ( .B1(inst1_n945), .B2(inst1_n1198), .A(inst1_n1099),
        .ZN(inst1_stateArray_S32reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst1_U1039 ( .B1(plaintext1[13]), .B2(inst1_n522), .A(inst1_n1095),
        .ZN(inst1_n1099) );
  OAI22_X1 inst1_U1038 ( .A1(inst1_n937), .A2(inst1_n1145), .B1(inst1_n1182),
        .B2(inst1_n1253), .ZN(inst1_n1095) );
  OAI21_X1 inst1_U1037 ( .B1(inst1_n946), .B2(inst1_n1198), .A(inst1_n1083),
        .ZN(inst1_stateArray_S32reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst1_U1036 ( .B1(plaintext1[14]), .B2(inst1_n596), .A(inst1_n1078),
        .ZN(inst1_n1083) );
  OAI22_X1 inst1_U1035 ( .A1(inst1_n938), .A2(inst1_n1145), .B1(inst1_n1182),
        .B2(inst1_n1251), .ZN(inst1_n1078) );
  OAI21_X1 inst1_U1034 ( .B1(inst1_n947), .B2(inst1_n1198), .A(inst1_n1069),
        .ZN(inst1_stateArray_S32reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst1_U1033 ( .B1(plaintext1[15]), .B2(inst1_n596), .A(inst1_n1068),
        .ZN(inst1_n1069) );
  OAI22_X1 inst1_U1032 ( .A1(inst1_n939), .A2(inst1_n1145), .B1(inst1_n1185),
        .B2(inst1_n1252), .ZN(inst1_n1068) );
  INV_X1 inst1_U1031 ( .A(inst1_n1135), .ZN(done1) );
  OAI211_X1 inst1_U1030 ( .C1(inst1_n1072), .C2(inst1_n1217), .A(inst1_n6),
        .B(inst1_n1066), .ZN(inst1_calcRCon_n48) );
  OAI221_X1 inst1_U1029 ( .B1(inst1_n1073), .B2(inst1_n1070), .C1(inst1_n1263),
        .C2(inst1_n1226), .A(inst1_n1217), .ZN(inst1_n1066) );
  OAI21_X1 inst1_U1028 ( .B1(inst1_n916), .B2(inst1_n1198), .A(inst1_n1065),
        .ZN(inst1_stateArray_S22reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst1_U1027 ( .B1(plaintext1[40]), .B2(inst1_n710), .A(inst1_n1064),
        .ZN(inst1_n1065) );
  OAI22_X1 inst1_U1026 ( .A1(inst1_n908), .A2(inst1_n1145), .B1(inst1_n1182),
        .B2(inst1_n1233), .ZN(inst1_n1064) );
  OAI211_X1 inst1_U1025 ( .C1(inst1_n937), .C2(inst1_n1198), .A(inst1_n1063),
        .B(inst1_n1062), .ZN(inst1_stateArray_S31reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst1_U1024 ( .A1(plaintext1[21]), .A2(inst1_n710), .ZN(inst1_n1062) );
  AOI22_X1 inst1_U1023 ( .A1(inst1_n677), .A2(ciphertext1[21]), .B1(
        inst1_n1217), .B2(ciphertext1[29]), .ZN(inst1_n1063) );
  OAI21_X1 inst1_U1022 ( .B1(inst1_n917), .B2(inst1_n1198), .A(inst1_n1053),
        .ZN(inst1_stateArray_S22reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst1_U1021 ( .B1(plaintext1[41]), .B2(inst1_n732), .A(inst1_n1045),
        .ZN(inst1_n1053) );
  OAI22_X1 inst1_U1020 ( .A1(inst1_n909), .A2(inst1_n1145), .B1(inst1_n1182),
        .B2(inst1_n1235), .ZN(inst1_n1045) );
  OAI21_X1 inst1_U1019 ( .B1(inst1_n918), .B2(inst1_n1198), .A(inst1_n1043),
        .ZN(inst1_stateArray_S22reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst1_U1018 ( .B1(plaintext1[42]), .B2(inst1_n830), .A(inst1_n1042),
        .ZN(inst1_n1043) );
  OAI22_X1 inst1_U1017 ( .A1(inst1_n1119), .A2(inst1_n1185), .B1(inst1_n910),
        .B2(inst1_n1142), .ZN(inst1_n1042) );
  OAI21_X1 inst1_U1016 ( .B1(inst1_n919), .B2(inst1_n1198), .A(inst1_n1041),
        .ZN(inst1_stateArray_S22reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst1_U1015 ( .B1(plaintext1[43]), .B2(inst1_n1133), .A(inst1_n1040), .ZN(inst1_n1041) );
  OAI22_X1 inst1_U1014 ( .A1(inst1_n1116), .A2(inst1_n1185), .B1(inst1_n911),
        .B2(inst1_n1142), .ZN(inst1_n1040) );
  OAI21_X1 inst1_U1013 ( .B1(inst1_n922), .B2(inst1_n1198), .A(inst1_n1039),
        .ZN(inst1_stateArray_S22reg_gff_1_SFF_6_n6) );
  AOI21_X1 inst1_U1012 ( .B1(plaintext1[46]), .B2(inst1_n1133), .A(inst1_n1038), .ZN(inst1_n1039) );
  OAI22_X1 inst1_U1011 ( .A1(inst1_n914), .A2(inst1_n1145), .B1(inst1_n1185),
        .B2(inst1_n1232), .ZN(inst1_n1038) );
  OAI21_X1 inst1_U1010 ( .B1(inst1_n923), .B2(inst1_n1198), .A(inst1_n1037),
        .ZN(inst1_stateArray_S22reg_gff_1_SFF_7_n6) );
  AOI21_X1 inst1_U1009 ( .B1(plaintext1[47]), .B2(inst1_n1133), .A(inst1_n1036), .ZN(inst1_n1037) );
  OAI22_X1 inst1_U1008 ( .A1(inst1_n1093), .A2(inst1_n1185), .B1(inst1_n915),
        .B2(inst1_n1145), .ZN(inst1_n1036) );
  OAI211_X1 inst1_U1007 ( .C1(inst1_n957), .C2(inst1_n1035), .A(inst1_n1034),
        .B(inst1_n1033), .ZN(inst1_KeyArray_S01reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst1_U1006 ( .A1(inst1_n1032), .A2(inst1_n137), .ZN(inst1_n1033)
         );
  AOI22_X1 inst1_U1005 ( .A1(inst1_n1031), .A2(inst1_n1271), .B1(key1[113]),
        .B2(inst1_n1228), .ZN(inst1_n1034) );
  OAI211_X1 inst1_U1004 ( .C1(inst1_n958), .C2(inst1_n1035), .A(inst1_n1030),
        .B(inst1_n1029), .ZN(inst1_KeyArray_S01reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst1_U1003 ( .A1(inst1_n1032), .A2(inst1_n136), .ZN(inst1_n1029)
         );
  AOI22_X1 inst1_U1002 ( .A1(inst1_n1031), .A2(inst1_n1270), .B1(key1[114]),
        .B2(inst1_n1228), .ZN(inst1_n1030) );
  OAI211_X1 inst1_U1001 ( .C1(inst1_n959), .C2(inst1_n1035), .A(inst1_n1028),
        .B(inst1_n1027), .ZN(inst1_KeyArray_S01reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst1_U1000 ( .A1(inst1_n1032), .A2(inst1_n135), .ZN(inst1_n1027)
         );
  AOI22_X1 inst1_U999 ( .A1(inst1_n1031), .A2(inst1_n1269), .B1(key1[115]),
        .B2(inst1_n1228), .ZN(inst1_n1028) );
  OAI211_X1 inst1_U998 ( .C1(inst1_n960), .C2(inst1_n1035), .A(inst1_n1026),
        .B(inst1_n1025), .ZN(inst1_KeyArray_S01reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst1_U997 ( .A1(inst1_n1032), .A2(inst1_n134), .ZN(inst1_n1025) );
  AOI22_X1 inst1_U996 ( .A1(inst1_n1031), .A2(inst1_n1268), .B1(key1[116]),
        .B2(inst1_n1228), .ZN(inst1_n1026) );
  OAI211_X1 inst1_U995 ( .C1(inst1_n961), .C2(inst1_n1035), .A(inst1_n1024),
        .B(inst1_n1023), .ZN(inst1_KeyArray_S01reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst1_U994 ( .A1(inst1_n1032), .A2(inst1_n133), .ZN(inst1_n1023) );
  AOI22_X1 inst1_U993 ( .A1(inst1_n1031), .A2(inst1_n1267), .B1(key1[117]),
        .B2(inst1_n1228), .ZN(inst1_n1024) );
  OAI211_X1 inst1_U992 ( .C1(inst1_n962), .C2(inst1_n1035), .A(inst1_n1022),
        .B(inst1_n1021), .ZN(inst1_KeyArray_S01reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst1_U991 ( .A1(inst1_n1032), .A2(inst1_n132), .ZN(inst1_n1021) );
  AOI22_X1 inst1_U990 ( .A1(inst1_n1031), .A2(inst1_n1266), .B1(key1[118]),
        .B2(inst1_n1228), .ZN(inst1_n1022) );
  OAI211_X1 inst1_U989 ( .C1(inst1_n963), .C2(inst1_n1035), .A(inst1_n1020),
        .B(inst1_n1019), .ZN(inst1_KeyArray_S01reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst1_U988 ( .A1(inst1_n1018), .A2(inst1_n131), .ZN(inst1_n1019) );
  AOI22_X1 inst1_U987 ( .A1(inst1_n1031), .A2(inst1_n1265), .B1(key1[119]),
        .B2(inst1_n1228), .ZN(inst1_n1020) );
  OAI21_X1 inst1_U986 ( .B1(inst1_n740), .B2(inst1_n1297), .A(inst1_n1017),
        .ZN(inst1_KeyArray_S02reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst1_U985 ( .B1(key1[104]), .B2(inst1_n1133), .A(inst1_n1016),
        .ZN(inst1_n1017) );
  OAI22_X1 inst1_U984 ( .A1(inst1_n964), .A2(inst1_n1015), .B1(inst1_n956),
        .B2(inst1_n1222), .ZN(inst1_n1016) );
  OAI21_X1 inst1_U983 ( .B1(inst1_n849), .B2(inst1_n1296), .A(inst1_n1014),
        .ZN(inst1_KeyArray_S02reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst1_U982 ( .B1(key1[105]), .B2(inst1_n1133), .A(inst1_n1013),
        .ZN(inst1_n1014) );
  OAI22_X1 inst1_U981 ( .A1(inst1_n965), .A2(inst1_n1015), .B1(inst1_n957),
        .B2(inst1_n1222), .ZN(inst1_n1013) );
  OAI21_X1 inst1_U980 ( .B1(inst1_n686), .B2(inst1_n1295), .A(inst1_n1012),
        .ZN(inst1_KeyArray_S02reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst1_U979 ( .B1(key1[106]), .B2(inst1_n1133), .A(inst1_n1011),
        .ZN(inst1_n1012) );
  OAI22_X1 inst1_U978 ( .A1(inst1_n966), .A2(inst1_n1203), .B1(inst1_n958),
        .B2(inst1_n1222), .ZN(inst1_n1011) );
  OAI21_X1 inst1_U977 ( .B1(inst1_n849), .B2(inst1_n1294), .A(inst1_n1010),
        .ZN(inst1_KeyArray_S02reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst1_U976 ( .B1(key1[107]), .B2(inst1_n1133), .A(inst1_n1009),
        .ZN(inst1_n1010) );
  OAI22_X1 inst1_U975 ( .A1(inst1_n967), .A2(inst1_n1035), .B1(inst1_n959),
        .B2(inst1_n1222), .ZN(inst1_n1009) );
  OAI21_X1 inst1_U974 ( .B1(inst1_n740), .B2(inst1_n1293), .A(inst1_n1008),
        .ZN(inst1_KeyArray_S02reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst1_U973 ( .B1(key1[108]), .B2(inst1_n1133), .A(inst1_n1007),
        .ZN(inst1_n1008) );
  OAI22_X1 inst1_U972 ( .A1(inst1_n968), .A2(inst1_n1203), .B1(inst1_n960),
        .B2(inst1_n1006), .ZN(inst1_n1007) );
  OAI21_X1 inst1_U971 ( .B1(inst1_n740), .B2(inst1_n1292), .A(inst1_n1005),
        .ZN(inst1_KeyArray_S02reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst1_U970 ( .B1(key1[109]), .B2(inst1_n1133), .A(inst1_n1004),
        .ZN(inst1_n1005) );
  OAI22_X1 inst1_U969 ( .A1(inst1_n969), .A2(inst1_n1203), .B1(inst1_n961),
        .B2(inst1_n1222), .ZN(inst1_n1004) );
  OAI21_X1 inst1_U968 ( .B1(inst1_n686), .B2(inst1_n1291), .A(inst1_n1003),
        .ZN(inst1_KeyArray_S02reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst1_U967 ( .B1(key1[110]), .B2(inst1_n1133), .A(inst1_n1002),
        .ZN(inst1_n1003) );
  OAI22_X1 inst1_U966 ( .A1(inst1_n970), .A2(inst1_n1203), .B1(inst1_n962),
        .B2(inst1_n1006), .ZN(inst1_n1002) );
  OAI21_X1 inst1_U965 ( .B1(inst1_n849), .B2(inst1_n1290), .A(inst1_n1001),
        .ZN(inst1_KeyArray_S02reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst1_U964 ( .B1(key1[111]), .B2(inst1_n1133), .A(inst1_n1000),
        .ZN(inst1_n1001) );
  OAI22_X1 inst1_U963 ( .A1(inst1_n971), .A2(inst1_n1203), .B1(inst1_n963),
        .B2(inst1_n1006), .ZN(inst1_n1000) );
  OAI21_X1 inst1_U962 ( .B1(inst1_n849), .B2(inst1_n1287), .A(inst1_n999),
        .ZN(inst1_KeyArray_S03reg_gff_1_SFF_0_n5) );
  AOI21_X1 inst1_U961 ( .B1(key1[96]), .B2(inst1_n710), .A(inst1_n998), .ZN(
        inst1_n999) );
  OAI22_X1 inst1_U960 ( .A1(inst1_n972), .A2(inst1_n1035), .B1(inst1_n964),
        .B2(inst1_n997), .ZN(inst1_n998) );
  OAI21_X1 inst1_U959 ( .B1(inst1_n740), .B2(inst1_n1286), .A(inst1_n996),
        .ZN(inst1_KeyArray_S03reg_gff_1_SFF_1_n5) );
  AOI21_X1 inst1_U958 ( .B1(key1[97]), .B2(inst1_n522), .A(inst1_n995), .ZN(
        inst1_n996) );
  OAI22_X1 inst1_U957 ( .A1(inst1_n973), .A2(inst1_n1035), .B1(inst1_n965),
        .B2(inst1_n997), .ZN(inst1_n995) );
  OAI21_X1 inst1_U956 ( .B1(inst1_n849), .B2(inst1_n1285), .A(inst1_n994),
        .ZN(inst1_KeyArray_S03reg_gff_1_SFF_2_n5) );
  AOI21_X1 inst1_U955 ( .B1(key1[98]), .B2(inst1_n596), .A(inst1_n993), .ZN(
        inst1_n994) );
  OAI22_X1 inst1_U954 ( .A1(inst1_n974), .A2(inst1_n1035), .B1(inst1_n966),
        .B2(inst1_n997), .ZN(inst1_n993) );
  OAI21_X1 inst1_U953 ( .B1(inst1_n686), .B2(inst1_n1284), .A(inst1_n992),
        .ZN(inst1_KeyArray_S03reg_gff_1_SFF_3_n5) );
  AOI21_X1 inst1_U952 ( .B1(key1[99]), .B2(inst1_n494), .A(inst1_n991), .ZN(
        inst1_n992) );
  OAI22_X1 inst1_U951 ( .A1(inst1_n975), .A2(inst1_n1203), .B1(inst1_n967),
        .B2(inst1_n997), .ZN(inst1_n991) );
  OAI21_X1 inst1_U950 ( .B1(inst1_n740), .B2(inst1_n1283), .A(inst1_n990),
        .ZN(inst1_KeyArray_S03reg_gff_1_SFF_4_n5) );
  AOI21_X1 inst1_U949 ( .B1(key1[100]), .B2(inst1_n1156), .A(inst1_n989), .ZN(
        inst1_n990) );
  OAI22_X1 inst1_U948 ( .A1(inst1_n976), .A2(inst1_n1203), .B1(inst1_n968),
        .B2(inst1_n997), .ZN(inst1_n989) );
  OAI21_X1 inst1_U947 ( .B1(inst1_n740), .B2(inst1_n1282), .A(inst1_n988),
        .ZN(inst1_KeyArray_S03reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst1_U946 ( .B1(key1[101]), .B2(inst1_n710), .A(inst1_n987), .ZN(
        inst1_n988) );
  OAI22_X1 inst1_U945 ( .A1(inst1_n977), .A2(inst1_n1035), .B1(inst1_n969),
        .B2(inst1_n997), .ZN(inst1_n987) );
  OAI21_X1 inst1_U944 ( .B1(inst1_n849), .B2(inst1_n1281), .A(inst1_n986),
        .ZN(inst1_KeyArray_S03reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst1_U943 ( .B1(key1[102]), .B2(inst1_n494), .A(inst1_n985), .ZN(
        inst1_n986) );
  OAI22_X1 inst1_U942 ( .A1(inst1_n978), .A2(inst1_n1203), .B1(inst1_n970),
        .B2(inst1_n997), .ZN(inst1_n985) );
  OAI21_X1 inst1_U941 ( .B1(inst1_n740), .B2(inst1_n1280), .A(inst1_n984),
        .ZN(inst1_KeyArray_S03reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst1_U940 ( .B1(key1[103]), .B2(inst1_n494), .A(inst1_n983), .ZN(
        inst1_n984) );
  OAI22_X1 inst1_U939 ( .A1(inst1_n979), .A2(inst1_n1035), .B1(inst1_n971),
        .B2(inst1_n997), .ZN(inst1_n983) );
  OAI21_X1 inst1_U938 ( .B1(inst1_n686), .B2(inst1_n1289), .A(inst1_n982),
        .ZN(inst1_KeyArray_S10reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst1_U937 ( .B1(key1[88]), .B2(inst1_n899), .A(inst1_n981), .ZN(
        inst1_n982) );
  OAI22_X1 inst1_U936 ( .A1(inst1_n972), .A2(inst1_n1006), .B1(inst1_n980),
        .B2(inst1_n1203), .ZN(inst1_n981) );
  OAI211_X1 inst1_U935 ( .C1(inst1_n973), .C2(inst1_n1222), .A(inst1_n931),
        .B(inst1_n930), .ZN(inst1_KeyArray_S10reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst1_U934 ( .A1(inst1_n1018), .A2(inst1_n121), .ZN(inst1_n930) );
  AOI22_X1 inst1_U933 ( .A1(inst1_n137), .A2(inst1_n929), .B1(key1[89]), .B2(
        inst1_n1228), .ZN(inst1_n931) );
  OAI211_X1 inst1_U932 ( .C1(inst1_n974), .C2(inst1_n1222), .A(inst1_n928),
        .B(inst1_n927), .ZN(inst1_KeyArray_S10reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst1_U931 ( .A1(inst1_n1018), .A2(inst1_n120), .ZN(inst1_n927) );
  AOI22_X1 inst1_U930 ( .A1(inst1_n136), .A2(inst1_n926), .B1(key1[90]), .B2(
        inst1_n1228), .ZN(inst1_n928) );
  OAI211_X1 inst1_U929 ( .C1(inst1_n975), .C2(inst1_n1222), .A(inst1_n925),
        .B(inst1_n924), .ZN(inst1_KeyArray_S10reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst1_U928 ( .A1(inst1_n1032), .A2(inst1_n119), .ZN(inst1_n924) );
  AOI22_X1 inst1_U927 ( .A1(inst1_n135), .A2(inst1_n926), .B1(key1[91]), .B2(
        inst1_n1228), .ZN(inst1_n925) );
  OAI211_X1 inst1_U926 ( .C1(inst1_n976), .C2(inst1_n1222), .A(inst1_n907),
        .B(inst1_n906), .ZN(inst1_KeyArray_S10reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst1_U925 ( .A1(inst1_n1032), .A2(inst1_n118), .ZN(inst1_n906) );
  AOI22_X1 inst1_U924 ( .A1(inst1_n134), .A2(inst1_n926), .B1(key1[92]), .B2(
        inst1_n1228), .ZN(inst1_n907) );
  OAI211_X1 inst1_U923 ( .C1(inst1_n977), .C2(inst1_n1222), .A(inst1_n905),
        .B(inst1_n904), .ZN(inst1_KeyArray_S10reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst1_U922 ( .A1(inst1_n1018), .A2(inst1_n117), .ZN(inst1_n904) );
  AOI22_X1 inst1_U921 ( .A1(inst1_n133), .A2(inst1_n926), .B1(key1[93]), .B2(
        inst1_n1228), .ZN(inst1_n905) );
  OAI211_X1 inst1_U920 ( .C1(inst1_n978), .C2(inst1_n1222), .A(inst1_n903),
        .B(inst1_n902), .ZN(inst1_KeyArray_S10reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst1_U919 ( .A1(inst1_n1032), .A2(inst1_n116), .ZN(inst1_n902) );
  AOI22_X1 inst1_U918 ( .A1(inst1_n132), .A2(inst1_n926), .B1(key1[94]), .B2(
        inst1_n1228), .ZN(inst1_n903) );
  OAI211_X1 inst1_U917 ( .C1(inst1_n979), .C2(inst1_n1222), .A(inst1_n901),
        .B(inst1_n900), .ZN(inst1_KeyArray_S10reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst1_U916 ( .A1(inst1_n1032), .A2(inst1_n115), .ZN(inst1_n900) );
  AOI22_X1 inst1_U915 ( .A1(inst1_n131), .A2(inst1_n926), .B1(key1[95]), .B2(
        inst1_n899), .ZN(inst1_n901) );
  OAI211_X1 inst1_U914 ( .C1(inst1_n980), .C2(inst1_n1222), .A(inst1_n898),
        .B(inst1_n897), .ZN(inst1_KeyArray_S11reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst1_U913 ( .A1(inst1_n1032), .A2(inst1_n114), .ZN(inst1_n897) );
  AOI22_X1 inst1_U912 ( .A1(inst1_n130), .A2(inst1_n926), .B1(key1[80]), .B2(
        inst1_n899), .ZN(inst1_n898) );
  NAND2_X1 inst1_U911 ( .A1(inst1_n896), .A2(inst1_n895), .ZN(
        inst1_KeyArray_S11reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U910 ( .A1(inst1_n1031), .A2(inst1_n137), .B1(inst1_n1032),
        .B2(inst1_n113), .ZN(inst1_n895) );
  AOI22_X1 inst1_U909 ( .A1(inst1_n129), .A2(inst1_n894), .B1(key1[81]), .B2(
        inst1_n899), .ZN(inst1_n896) );
  NAND2_X1 inst1_U908 ( .A1(inst1_n893), .A2(inst1_n892), .ZN(
        inst1_KeyArray_S11reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U907 ( .A1(inst1_n1031), .A2(inst1_n136), .B1(inst1_n1032),
        .B2(inst1_n112), .ZN(inst1_n892) );
  AOI22_X1 inst1_U906 ( .A1(inst1_n128), .A2(inst1_n894), .B1(key1[82]), .B2(
        inst1_n899), .ZN(inst1_n893) );
  NAND2_X1 inst1_U905 ( .A1(inst1_n867), .A2(inst1_n866), .ZN(
        inst1_KeyArray_S11reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U904 ( .A1(inst1_n1031), .A2(inst1_n135), .B1(inst1_n1018),
        .B2(inst1_n111), .ZN(inst1_n866) );
  AOI22_X1 inst1_U903 ( .A1(inst1_n127), .A2(inst1_n894), .B1(key1[83]), .B2(
        inst1_n899), .ZN(inst1_n867) );
  NAND2_X1 inst1_U902 ( .A1(inst1_n865), .A2(inst1_n864), .ZN(
        inst1_KeyArray_S11reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U901 ( .A1(inst1_n1031), .A2(inst1_n134), .B1(inst1_n1032),
        .B2(inst1_n110), .ZN(inst1_n864) );
  AOI22_X1 inst1_U900 ( .A1(inst1_n126), .A2(inst1_n894), .B1(key1[84]), .B2(
        inst1_n899), .ZN(inst1_n865) );
  NAND2_X1 inst1_U899 ( .A1(inst1_n863), .A2(inst1_n862), .ZN(
        inst1_KeyArray_S11reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst1_U898 ( .A1(inst1_n1031), .A2(inst1_n133), .B1(inst1_n1032),
        .B2(inst1_n109), .ZN(inst1_n862) );
  INV_X1 inst1_U897 ( .A(inst1_n997), .ZN(inst1_n1031) );
  AOI22_X1 inst1_U896 ( .A1(inst1_n125), .A2(inst1_n894), .B1(key1[85]), .B2(
        inst1_n899), .ZN(inst1_n863) );
  NAND2_X1 inst1_U895 ( .A1(inst1_n861), .A2(inst1_n860), .ZN(
        inst1_KeyArray_S11reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst1_U894 ( .A1(inst1_n859), .A2(inst1_n132), .B1(inst1_n1032),
        .B2(inst1_n108), .ZN(inst1_n860) );
  AOI22_X1 inst1_U893 ( .A1(inst1_n124), .A2(inst1_n894), .B1(key1[86]), .B2(
        inst1_n899), .ZN(inst1_n861) );
  NAND2_X1 inst1_U892 ( .A1(inst1_n858), .A2(inst1_n857), .ZN(
        inst1_KeyArray_S11reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst1_U891 ( .A1(inst1_n859), .A2(inst1_n131), .B1(inst1_n1018),
        .B2(inst1_n107), .ZN(inst1_n857) );
  AOI22_X1 inst1_U890 ( .A1(inst1_n123), .A2(inst1_n894), .B1(key1[87]), .B2(
        inst1_n899), .ZN(inst1_n858) );
  OAI21_X1 inst1_U889 ( .B1(inst1_n956), .B2(inst1_n740), .A(inst1_n856), .ZN(
        inst1_KeyArray_S32reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst1_U888 ( .B1(key1[8]), .B2(inst1_n830), .A(inst1_n855), .ZN(
        inst1_n856) );
  OAI22_X1 inst1_U887 ( .A1(inst1_n1052), .A2(inst1_n1035), .B1(inst1_n1044),
        .B2(inst1_n1222), .ZN(inst1_n855) );
  OAI21_X1 inst1_U886 ( .B1(inst1_n958), .B2(inst1_n686), .A(inst1_n854), .ZN(
        inst1_KeyArray_S32reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst1_U885 ( .B1(key1[10]), .B2(inst1_n732), .A(inst1_n853), .ZN(
        inst1_n854) );
  OAI22_X1 inst1_U884 ( .A1(inst1_n1054), .A2(inst1_n1203), .B1(inst1_n1046),
        .B2(inst1_n1222), .ZN(inst1_n853) );
  OAI21_X1 inst1_U883 ( .B1(inst1_n959), .B2(inst1_n740), .A(inst1_n852), .ZN(
        inst1_KeyArray_S32reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst1_U882 ( .B1(key1[11]), .B2(inst1_n507), .A(inst1_n850), .ZN(
        inst1_n852) );
  OAI22_X1 inst1_U881 ( .A1(inst1_n1055), .A2(inst1_n1203), .B1(inst1_n1047),
        .B2(inst1_n997), .ZN(inst1_n850) );
  OAI21_X1 inst1_U880 ( .B1(inst1_n960), .B2(inst1_n849), .A(inst1_n848), .ZN(
        inst1_KeyArray_S32reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst1_U879 ( .B1(key1[12]), .B2(inst1_n1156), .A(inst1_n847), .ZN(
        inst1_n848) );
  OAI22_X1 inst1_U878 ( .A1(inst1_n1056), .A2(inst1_n1203), .B1(inst1_n1048),
        .B2(inst1_n1006), .ZN(inst1_n847) );
  OAI21_X1 inst1_U877 ( .B1(inst1_n961), .B2(inst1_n849), .A(inst1_n846), .ZN(
        inst1_KeyArray_S32reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst1_U876 ( .B1(key1[13]), .B2(inst1_n522), .A(inst1_n845), .ZN(
        inst1_n846) );
  OAI22_X1 inst1_U875 ( .A1(inst1_n1057), .A2(inst1_n1035), .B1(inst1_n1049),
        .B2(inst1_n1222), .ZN(inst1_n845) );
  OAI21_X1 inst1_U874 ( .B1(inst1_n962), .B2(inst1_n740), .A(inst1_n844), .ZN(
        inst1_KeyArray_S32reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst1_U873 ( .B1(key1[14]), .B2(inst1_n522), .A(inst1_n843), .ZN(
        inst1_n844) );
  OAI22_X1 inst1_U872 ( .A1(inst1_n1058), .A2(inst1_n1035), .B1(inst1_n1050),
        .B2(inst1_n997), .ZN(inst1_n843) );
  OAI21_X1 inst1_U871 ( .B1(inst1_n963), .B2(inst1_n686), .A(inst1_n842), .ZN(
        inst1_KeyArray_S32reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst1_U870 ( .B1(key1[15]), .B2(inst1_n596), .A(inst1_n841), .ZN(
        inst1_n842) );
  OAI22_X1 inst1_U869 ( .A1(inst1_n1059), .A2(inst1_n1035), .B1(inst1_n1051),
        .B2(inst1_n997), .ZN(inst1_n841) );
  OAI21_X1 inst1_U868 ( .B1(inst1_n980), .B2(inst1_n849), .A(inst1_n840), .ZN(
        inst1_KeyArray_S01reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst1_U867 ( .B1(key1[112]), .B2(inst1_n830), .A(inst1_n839), .ZN(
        inst1_n840) );
  OAI22_X1 inst1_U866 ( .A1(inst1_n948), .A2(inst1_n1006), .B1(inst1_n956),
        .B2(inst1_n1203), .ZN(inst1_n839) );
  NAND2_X1 inst1_U865 ( .A1(inst1_n838), .A2(inst1_n837), .ZN(
        inst1_KeyArray_S12reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst1_U864 ( .A1(inst1_n859), .A2(inst1_n130), .B1(inst1_n1032),
        .B2(inst1_n98), .ZN(inst1_n837) );
  AOI22_X1 inst1_U863 ( .A1(inst1_n22), .A2(inst1_n894), .B1(key1[72]), .B2(
        inst1_n899), .ZN(inst1_n838) );
  NAND2_X1 inst1_U862 ( .A1(inst1_n836), .A2(inst1_n835), .ZN(
        inst1_KeyArray_S12reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U861 ( .A1(inst1_n859), .A2(inst1_n129), .B1(inst1_n1018),
        .B2(inst1_n97), .ZN(inst1_n835) );
  AOI22_X1 inst1_U860 ( .A1(inst1_n17), .A2(inst1_n894), .B1(key1[73]), .B2(
        inst1_n899), .ZN(inst1_n836) );
  NAND2_X1 inst1_U859 ( .A1(inst1_n834), .A2(inst1_n833), .ZN(
        inst1_KeyArray_S12reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U858 ( .A1(inst1_n859), .A2(inst1_n128), .B1(inst1_n1032),
        .B2(inst1_n96), .ZN(inst1_n833) );
  AOI22_X1 inst1_U857 ( .A1(inst1_n14), .A2(inst1_n894), .B1(key1[74]), .B2(
        inst1_n899), .ZN(inst1_n834) );
  INV_X1 inst1_U856 ( .A(inst1_n6), .ZN(inst1_n899) );
  NAND2_X1 inst1_U855 ( .A1(inst1_n832), .A2(inst1_n831), .ZN(
        inst1_KeyArray_S12reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U854 ( .A1(inst1_n859), .A2(inst1_n127), .B1(inst1_n1032),
        .B2(inst1_n95), .ZN(inst1_n831) );
  AOI22_X1 inst1_U853 ( .A1(inst1_n12), .A2(inst1_n894), .B1(key1[75]), .B2(
        inst1_n830), .ZN(inst1_n832) );
  NAND2_X1 inst1_U852 ( .A1(inst1_n829), .A2(inst1_n828), .ZN(
        inst1_KeyArray_S12reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U851 ( .A1(inst1_n827), .A2(inst1_n126), .B1(inst1_n1032),
        .B2(inst1_n94), .ZN(inst1_n828) );
  AOI22_X1 inst1_U850 ( .A1(inst1_n11), .A2(inst1_n894), .B1(key1[76]), .B2(
        inst1_n830), .ZN(inst1_n829) );
  NAND2_X1 inst1_U849 ( .A1(inst1_n826), .A2(inst1_n825), .ZN(
        inst1_KeyArray_S12reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst1_U848 ( .A1(inst1_n827), .A2(inst1_n125), .B1(inst1_n1032),
        .B2(inst1_n93), .ZN(inst1_n825) );
  AOI22_X1 inst1_U847 ( .A1(inst1_n10), .A2(inst1_n894), .B1(key1[77]), .B2(
        inst1_n830), .ZN(inst1_n826) );
  NAND2_X1 inst1_U846 ( .A1(inst1_n824), .A2(inst1_n823), .ZN(
        inst1_KeyArray_S12reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst1_U845 ( .A1(inst1_n859), .A2(inst1_n124), .B1(inst1_n1032),
        .B2(inst1_n92), .ZN(inst1_n823) );
  AOI22_X1 inst1_U844 ( .A1(inst1_n24), .A2(inst1_n822), .B1(key1[78]), .B2(
        inst1_n830), .ZN(inst1_n824) );
  NAND2_X1 inst1_U843 ( .A1(inst1_n821), .A2(inst1_n820), .ZN(
        inst1_KeyArray_S12reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst1_U842 ( .A1(inst1_n819), .A2(inst1_n123), .B1(inst1_n1032),
        .B2(inst1_n91), .ZN(inst1_n820) );
  AOI22_X1 inst1_U841 ( .A1(inst1_n9), .A2(inst1_n926), .B1(key1[79]), .B2(
        inst1_n830), .ZN(inst1_n821) );
  NAND2_X1 inst1_U840 ( .A1(inst1_n818), .A2(inst1_n817), .ZN(
        inst1_KeyArray_S13reg_gff_1_SFF_0_n5) );
  AOI22_X1 inst1_U839 ( .A1(inst1_n1031), .A2(inst1_n22), .B1(inst1_n1018),
        .B2(inst1_n90), .ZN(inst1_n817) );
  AOI22_X1 inst1_U838 ( .A1(inst1_n122), .A2(inst1_n929), .B1(key1[64]), .B2(
        inst1_n830), .ZN(inst1_n818) );
  NAND2_X1 inst1_U837 ( .A1(inst1_n816), .A2(inst1_n815), .ZN(
        inst1_KeyArray_S13reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst1_U836 ( .A1(inst1_n819), .A2(inst1_n17), .B1(inst1_n1018),
        .B2(inst1_n89), .ZN(inst1_n815) );
  AOI22_X1 inst1_U835 ( .A1(inst1_n121), .A2(inst1_n822), .B1(key1[65]), .B2(
        inst1_n830), .ZN(inst1_n816) );
  NAND2_X1 inst1_U834 ( .A1(inst1_n814), .A2(inst1_n813), .ZN(
        inst1_KeyArray_S13reg_gff_1_SFF_2_n5) );
  AOI22_X1 inst1_U833 ( .A1(inst1_n859), .A2(inst1_n14), .B1(inst1_n1032),
        .B2(inst1_n88), .ZN(inst1_n813) );
  AOI22_X1 inst1_U832 ( .A1(inst1_n120), .A2(inst1_n822), .B1(key1[66]), .B2(
        inst1_n830), .ZN(inst1_n814) );
  NAND2_X1 inst1_U831 ( .A1(inst1_n812), .A2(inst1_n811), .ZN(
        inst1_KeyArray_S13reg_gff_1_SFF_3_n5) );
  AOI22_X1 inst1_U830 ( .A1(inst1_n819), .A2(inst1_n12), .B1(inst1_n1032),
        .B2(inst1_n87), .ZN(inst1_n811) );
  AOI22_X1 inst1_U829 ( .A1(inst1_n119), .A2(inst1_n822), .B1(key1[67]), .B2(
        inst1_n830), .ZN(inst1_n812) );
  NAND2_X1 inst1_U828 ( .A1(inst1_n810), .A2(inst1_n809), .ZN(
        inst1_KeyArray_S13reg_gff_1_SFF_4_n5) );
  AOI22_X1 inst1_U827 ( .A1(inst1_n859), .A2(inst1_n11), .B1(inst1_n1032),
        .B2(inst1_n86), .ZN(inst1_n809) );
  AOI22_X1 inst1_U826 ( .A1(inst1_n118), .A2(inst1_n926), .B1(key1[68]), .B2(
        inst1_n830), .ZN(inst1_n810) );
  NAND2_X1 inst1_U825 ( .A1(inst1_n808), .A2(inst1_n807), .ZN(
        inst1_KeyArray_S13reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst1_U824 ( .A1(inst1_n819), .A2(inst1_n10), .B1(inst1_n1032),
        .B2(inst1_n85), .ZN(inst1_n807) );
  AOI22_X1 inst1_U823 ( .A1(inst1_n117), .A2(inst1_n929), .B1(key1[69]), .B2(
        inst1_n830), .ZN(inst1_n808) );
  NAND2_X1 inst1_U822 ( .A1(inst1_n806), .A2(inst1_n805), .ZN(
        inst1_KeyArray_S13reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst1_U821 ( .A1(inst1_n819), .A2(inst1_n24), .B1(inst1_n1018),
        .B2(inst1_n84), .ZN(inst1_n805) );
  AOI22_X1 inst1_U820 ( .A1(inst1_n116), .A2(inst1_n926), .B1(key1[70]), .B2(
        inst1_n732), .ZN(inst1_n806) );
  NAND2_X1 inst1_U819 ( .A1(inst1_n804), .A2(inst1_n803), .ZN(
        inst1_KeyArray_S13reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst1_U818 ( .A1(inst1_n859), .A2(inst1_n9), .B1(inst1_n1032), .B2(
        inst1_n83), .ZN(inst1_n803) );
  AOI22_X1 inst1_U817 ( .A1(inst1_n115), .A2(inst1_n926), .B1(key1[71]), .B2(
        inst1_n899), .ZN(inst1_n804) );
  NAND2_X1 inst1_U816 ( .A1(inst1_n802), .A2(inst1_n801), .ZN(
        inst1_KeyArray_S20reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst1_U815 ( .A1(inst1_n819), .A2(inst1_n122), .B1(inst1_n1032),
        .B2(inst1_n82), .ZN(inst1_n801) );
  AOI22_X1 inst1_U814 ( .A1(inst1_n114), .A2(inst1_n929), .B1(key1[56]), .B2(
        inst1_n494), .ZN(inst1_n802) );
  NAND2_X1 inst1_U813 ( .A1(inst1_n800), .A2(inst1_n799), .ZN(
        inst1_KeyArray_S20reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U812 ( .A1(inst1_n827), .A2(inst1_n121), .B1(inst1_n1018),
        .B2(inst1_n81), .ZN(inst1_n799) );
  AOI22_X1 inst1_U811 ( .A1(inst1_n113), .A2(inst1_n929), .B1(key1[57]), .B2(
        inst1_n507), .ZN(inst1_n800) );
  NAND2_X1 inst1_U810 ( .A1(inst1_n798), .A2(inst1_n797), .ZN(
        inst1_KeyArray_S20reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U809 ( .A1(inst1_n859), .A2(inst1_n120), .B1(inst1_n1032),
        .B2(inst1_n80), .ZN(inst1_n797) );
  AOI22_X1 inst1_U808 ( .A1(inst1_n112), .A2(inst1_n929), .B1(key1[58]), .B2(
        inst1_n1156), .ZN(inst1_n798) );
  NAND2_X1 inst1_U807 ( .A1(inst1_n796), .A2(inst1_n795), .ZN(
        inst1_KeyArray_S20reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U806 ( .A1(inst1_n859), .A2(inst1_n119), .B1(inst1_n1032),
        .B2(inst1_n79), .ZN(inst1_n795) );
  AOI22_X1 inst1_U805 ( .A1(inst1_n111), .A2(inst1_n929), .B1(key1[59]), .B2(
        inst1_n710), .ZN(inst1_n796) );
  NAND2_X1 inst1_U804 ( .A1(inst1_n794), .A2(inst1_n793), .ZN(
        inst1_KeyArray_S20reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U803 ( .A1(inst1_n1031), .A2(inst1_n118), .B1(inst1_n78),
        .B2(inst1_n1018), .ZN(inst1_n793) );
  AOI22_X1 inst1_U802 ( .A1(inst1_n110), .A2(inst1_n929), .B1(key1[60]), .B2(
        inst1_n596), .ZN(inst1_n794) );
  NAND2_X1 inst1_U801 ( .A1(inst1_n792), .A2(inst1_n791), .ZN(
        inst1_KeyArray_S20reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst1_U800 ( .A1(inst1_n819), .A2(inst1_n117), .B1(inst1_n1032),
        .B2(inst1_n77), .ZN(inst1_n791) );
  AOI22_X1 inst1_U799 ( .A1(inst1_n109), .A2(inst1_n929), .B1(key1[61]), .B2(
        inst1_n522), .ZN(inst1_n792) );
  NAND2_X1 inst1_U798 ( .A1(inst1_n790), .A2(inst1_n789), .ZN(
        inst1_KeyArray_S20reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst1_U797 ( .A1(inst1_n819), .A2(inst1_n116), .B1(inst1_n1032),
        .B2(inst1_n76), .ZN(inst1_n789) );
  AOI22_X1 inst1_U796 ( .A1(inst1_n108), .A2(inst1_n929), .B1(key1[62]), .B2(
        inst1_n596), .ZN(inst1_n790) );
  NAND2_X1 inst1_U795 ( .A1(inst1_n788), .A2(inst1_n787), .ZN(
        inst1_KeyArray_S20reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst1_U794 ( .A1(inst1_n819), .A2(inst1_n115), .B1(inst1_n1018),
        .B2(inst1_n75), .ZN(inst1_n787) );
  AOI22_X1 inst1_U793 ( .A1(inst1_n107), .A2(inst1_n929), .B1(key1[63]), .B2(
        inst1_n830), .ZN(inst1_n788) );
  NAND2_X1 inst1_U792 ( .A1(inst1_n786), .A2(inst1_n785), .ZN(
        inst1_KeyArray_S21reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst1_U791 ( .A1(inst1_n819), .A2(inst1_n114), .B1(inst1_n1032),
        .B2(inst1_n74), .ZN(inst1_n785) );
  AOI22_X1 inst1_U790 ( .A1(inst1_n98), .A2(inst1_n929), .B1(key1[48]), .B2(
        inst1_n732), .ZN(inst1_n786) );
  NAND2_X1 inst1_U789 ( .A1(inst1_n784), .A2(inst1_n783), .ZN(
        inst1_KeyArray_S21reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U788 ( .A1(inst1_n1031), .A2(inst1_n113), .B1(inst1_n1032),
        .B2(inst1_n73), .ZN(inst1_n783) );
  AOI22_X1 inst1_U787 ( .A1(inst1_n97), .A2(inst1_n929), .B1(key1[49]), .B2(
        inst1_n1156), .ZN(inst1_n784) );
  NAND2_X1 inst1_U786 ( .A1(inst1_n782), .A2(inst1_n781), .ZN(
        inst1_KeyArray_S21reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U785 ( .A1(inst1_n827), .A2(inst1_n112), .B1(inst1_n1018),
        .B2(inst1_n72), .ZN(inst1_n781) );
  AOI22_X1 inst1_U784 ( .A1(inst1_n96), .A2(inst1_n929), .B1(key1[50]), .B2(
        inst1_n899), .ZN(inst1_n782) );
  NAND2_X1 inst1_U783 ( .A1(inst1_n780), .A2(inst1_n779), .ZN(
        inst1_KeyArray_S21reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U782 ( .A1(inst1_n827), .A2(inst1_n111), .B1(inst1_n1032),
        .B2(inst1_n71), .ZN(inst1_n779) );
  AOI22_X1 inst1_U781 ( .A1(inst1_n95), .A2(inst1_n929), .B1(key1[51]), .B2(
        inst1_n830), .ZN(inst1_n780) );
  NAND2_X1 inst1_U780 ( .A1(inst1_n778), .A2(inst1_n777), .ZN(
        inst1_KeyArray_S21reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U779 ( .A1(inst1_n1031), .A2(inst1_n110), .B1(inst1_n70),
        .B2(inst1_n1032), .ZN(inst1_n777) );
  AOI22_X1 inst1_U778 ( .A1(inst1_n94), .A2(inst1_n929), .B1(key1[52]), .B2(
        inst1_n732), .ZN(inst1_n778) );
  NAND2_X1 inst1_U777 ( .A1(inst1_n776), .A2(inst1_n775), .ZN(
        inst1_KeyArray_S21reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst1_U776 ( .A1(inst1_n819), .A2(inst1_n109), .B1(inst1_n1032),
        .B2(inst1_n69), .ZN(inst1_n775) );
  AOI22_X1 inst1_U775 ( .A1(inst1_n93), .A2(inst1_n929), .B1(key1[53]), .B2(
        inst1_n899), .ZN(inst1_n776) );
  NAND2_X1 inst1_U774 ( .A1(inst1_n774), .A2(inst1_n773), .ZN(
        inst1_KeyArray_S21reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst1_U773 ( .A1(inst1_n1031), .A2(inst1_n108), .B1(inst1_n1032),
        .B2(inst1_n68), .ZN(inst1_n773) );
  AOI22_X1 inst1_U772 ( .A1(inst1_n92), .A2(inst1_n822), .B1(key1[54]), .B2(
        inst1_n507), .ZN(inst1_n774) );
  NAND2_X1 inst1_U771 ( .A1(inst1_n772), .A2(inst1_n771), .ZN(
        inst1_KeyArray_S21reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst1_U770 ( .A1(inst1_n827), .A2(inst1_n107), .B1(inst1_n1032),
        .B2(inst1_n67), .ZN(inst1_n771) );
  AOI22_X1 inst1_U769 ( .A1(inst1_n91), .A2(inst1_n926), .B1(key1[55]), .B2(
        inst1_n494), .ZN(inst1_n772) );
  OAI211_X1 inst1_U768 ( .C1(inst1_n1044), .C2(inst1_n849), .A(inst1_n770),
        .B(inst1_n769), .ZN(inst1_KeyArray_S22reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst1_U767 ( .A1(inst1_n1031), .A2(inst1_n98), .ZN(inst1_n769) );
  AOI22_X1 inst1_U766 ( .A1(inst1_n90), .A2(inst1_n929), .B1(key1[40]), .B2(
        inst1_n494), .ZN(inst1_n770) );
  NAND2_X1 inst1_U765 ( .A1(inst1_n768), .A2(inst1_n767), .ZN(
        inst1_KeyArray_S22reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U764 ( .A1(inst1_n819), .A2(inst1_n97), .B1(inst1_n1032),
        .B2(inst1_n65), .ZN(inst1_n767) );
  AOI22_X1 inst1_U763 ( .A1(inst1_n89), .A2(inst1_n929), .B1(key1[41]), .B2(
        inst1_n710), .ZN(inst1_n768) );
  OAI211_X1 inst1_U762 ( .C1(inst1_n1046), .C2(inst1_n686), .A(inst1_n766),
        .B(inst1_n765), .ZN(inst1_KeyArray_S22reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst1_U761 ( .A1(inst1_n1031), .A2(inst1_n96), .ZN(inst1_n765) );
  AOI22_X1 inst1_U760 ( .A1(inst1_n88), .A2(inst1_n926), .B1(key1[42]), .B2(
        inst1_n522), .ZN(inst1_n766) );
  OAI211_X1 inst1_U759 ( .C1(inst1_n1047), .C2(inst1_n849), .A(inst1_n764),
        .B(inst1_n763), .ZN(inst1_KeyArray_S22reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst1_U758 ( .A1(inst1_n859), .A2(inst1_n95), .ZN(inst1_n763) );
  AOI22_X1 inst1_U757 ( .A1(inst1_n87), .A2(inst1_n929), .B1(key1[43]), .B2(
        inst1_n522), .ZN(inst1_n764) );
  OAI211_X1 inst1_U756 ( .C1(inst1_n1048), .C2(inst1_n686), .A(inst1_n762),
        .B(inst1_n761), .ZN(inst1_KeyArray_S22reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst1_U755 ( .A1(inst1_n819), .A2(inst1_n94), .ZN(inst1_n761) );
  AOI22_X1 inst1_U754 ( .A1(inst1_n86), .A2(inst1_n822), .B1(key1[44]), .B2(
        inst1_n732), .ZN(inst1_n762) );
  OAI211_X1 inst1_U753 ( .C1(inst1_n1049), .C2(inst1_n849), .A(inst1_n760),
        .B(inst1_n759), .ZN(inst1_KeyArray_S22reg_gff_1_SFF_5_n5) );
  NAND2_X1 inst1_U752 ( .A1(inst1_n827), .A2(inst1_n93), .ZN(inst1_n759) );
  AOI22_X1 inst1_U751 ( .A1(inst1_n85), .A2(inst1_n822), .B1(key1[45]), .B2(
        inst1_n596), .ZN(inst1_n760) );
  OAI211_X1 inst1_U750 ( .C1(inst1_n1050), .C2(inst1_n686), .A(inst1_n758),
        .B(inst1_n757), .ZN(inst1_KeyArray_S22reg_gff_1_SFF_6_n5) );
  NAND2_X1 inst1_U749 ( .A1(inst1_n859), .A2(inst1_n92), .ZN(inst1_n757) );
  AOI22_X1 inst1_U748 ( .A1(inst1_n84), .A2(inst1_n926), .B1(key1[46]), .B2(
        inst1_n494), .ZN(inst1_n758) );
  OAI211_X1 inst1_U747 ( .C1(inst1_n1051), .C2(inst1_n849), .A(inst1_n756),
        .B(inst1_n755), .ZN(inst1_KeyArray_S22reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst1_U746 ( .A1(inst1_n1031), .A2(inst1_n91), .ZN(inst1_n755) );
  AOI22_X1 inst1_U745 ( .A1(inst1_n83), .A2(inst1_n822), .B1(key1[47]), .B2(
        inst1_n899), .ZN(inst1_n756) );
  OAI211_X1 inst1_U744 ( .C1(inst1_n1052), .C2(inst1_n740), .A(inst1_n754),
        .B(inst1_n753), .ZN(inst1_KeyArray_S23reg_gff_1_SFF_0_n5) );
  NAND2_X1 inst1_U743 ( .A1(inst1_n819), .A2(inst1_n90), .ZN(inst1_n753) );
  AOI22_X1 inst1_U742 ( .A1(inst1_n82), .A2(inst1_n926), .B1(key1[32]), .B2(
        inst1_n899), .ZN(inst1_n754) );
  NAND2_X1 inst1_U741 ( .A1(inst1_n752), .A2(inst1_n751), .ZN(
        inst1_KeyArray_S23reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst1_U740 ( .A1(inst1_n827), .A2(inst1_n89), .B1(inst1_n1018),
        .B2(inst1_n57), .ZN(inst1_n751) );
  AOI22_X1 inst1_U739 ( .A1(inst1_n81), .A2(inst1_n929), .B1(key1[33]), .B2(
        inst1_n1156), .ZN(inst1_n752) );
  OAI211_X1 inst1_U738 ( .C1(inst1_n1054), .C2(inst1_n686), .A(inst1_n750),
        .B(inst1_n749), .ZN(inst1_KeyArray_S23reg_gff_1_SFF_2_n5) );
  NAND2_X1 inst1_U737 ( .A1(inst1_n827), .A2(inst1_n88), .ZN(inst1_n749) );
  AOI22_X1 inst1_U736 ( .A1(inst1_n80), .A2(inst1_n822), .B1(key1[34]), .B2(
        inst1_n507), .ZN(inst1_n750) );
  OAI211_X1 inst1_U735 ( .C1(inst1_n1055), .C2(inst1_n740), .A(inst1_n748),
        .B(inst1_n747), .ZN(inst1_KeyArray_S23reg_gff_1_SFF_3_n5) );
  NAND2_X1 inst1_U734 ( .A1(inst1_n859), .A2(inst1_n87), .ZN(inst1_n747) );
  AOI22_X1 inst1_U733 ( .A1(inst1_n79), .A2(inst1_n822), .B1(key1[35]), .B2(
        inst1_n710), .ZN(inst1_n748) );
  OAI211_X1 inst1_U732 ( .C1(inst1_n1056), .C2(inst1_n849), .A(inst1_n746),
        .B(inst1_n745), .ZN(inst1_KeyArray_S23reg_gff_1_SFF_4_n5) );
  NAND2_X1 inst1_U731 ( .A1(inst1_n1031), .A2(inst1_n86), .ZN(inst1_n745) );
  AOI22_X1 inst1_U730 ( .A1(inst1_n926), .A2(inst1_n78), .B1(key1[36]), .B2(
        inst1_n596), .ZN(inst1_n746) );
  OAI211_X1 inst1_U729 ( .C1(inst1_n1057), .C2(inst1_n686), .A(inst1_n744),
        .B(inst1_n743), .ZN(inst1_KeyArray_S23reg_gff_1_SFF_5_n5) );
  NAND2_X1 inst1_U728 ( .A1(inst1_n819), .A2(inst1_n85), .ZN(inst1_n743) );
  AOI22_X1 inst1_U727 ( .A1(inst1_n77), .A2(inst1_n926), .B1(key1[37]), .B2(
        inst1_n1156), .ZN(inst1_n744) );
  OAI211_X1 inst1_U726 ( .C1(inst1_n1058), .C2(inst1_n686), .A(inst1_n742),
        .B(inst1_n741), .ZN(inst1_KeyArray_S23reg_gff_1_SFF_6_n5) );
  NAND2_X1 inst1_U725 ( .A1(inst1_n859), .A2(inst1_n84), .ZN(inst1_n741) );
  AOI22_X1 inst1_U724 ( .A1(inst1_n76), .A2(inst1_n929), .B1(key1[38]), .B2(
        inst1_n522), .ZN(inst1_n742) );
  OAI211_X1 inst1_U723 ( .C1(inst1_n1059), .C2(inst1_n740), .A(inst1_n739),
        .B(inst1_n738), .ZN(inst1_KeyArray_S23reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst1_U722 ( .A1(inst1_n827), .A2(inst1_n83), .ZN(inst1_n738) );
  AOI22_X1 inst1_U721 ( .A1(inst1_n75), .A2(inst1_n822), .B1(key1[39]), .B2(
        inst1_n1156), .ZN(inst1_n739) );
  OAI21_X1 inst1_U720 ( .B1(inst1_n948), .B2(inst1_n849), .A(inst1_n737), .ZN(
        inst1_KeyArray_S31reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst1_U719 ( .B1(key1[16]), .B2(inst1_n732), .A(inst1_n736), .ZN(
        inst1_n737) );
  OAI22_X1 inst1_U718 ( .A1(inst1_n1044), .A2(inst1_n1203), .B1(inst1_n1222),
        .B2(inst1_n1239), .ZN(inst1_n736) );
  OAI211_X1 inst1_U717 ( .C1(inst1_n949), .C2(inst1_n740), .A(inst1_n735), .B(
        inst1_n734), .ZN(inst1_KeyArray_S31reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst1_U716 ( .A1(inst1_n1031), .A2(inst1_n73), .ZN(inst1_n734) );
  AOI22_X1 inst1_U715 ( .A1(inst1_n65), .A2(inst1_n929), .B1(key1[17]), .B2(
        inst1_n494), .ZN(inst1_n735) );
  INV_X1 inst1_U714 ( .A(inst1_n1015), .ZN(inst1_n929) );
  OAI21_X1 inst1_U713 ( .B1(inst1_n950), .B2(inst1_n849), .A(inst1_n733), .ZN(
        inst1_KeyArray_S31reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst1_U712 ( .B1(key1[18]), .B2(inst1_n732), .A(inst1_n731), .ZN(
        inst1_n733) );
  OAI22_X1 inst1_U711 ( .A1(inst1_n1046), .A2(inst1_n1203), .B1(inst1_n1222),
        .B2(inst1_n1238), .ZN(inst1_n731) );
  OAI21_X1 inst1_U710 ( .B1(inst1_n951), .B2(inst1_n849), .A(inst1_n730), .ZN(
        inst1_KeyArray_S31reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst1_U709 ( .B1(key1[19]), .B2(inst1_n899), .A(inst1_n729), .ZN(
        inst1_n730) );
  OAI22_X1 inst1_U708 ( .A1(inst1_n1047), .A2(inst1_n1203), .B1(inst1_n1222),
        .B2(inst1_n1262), .ZN(inst1_n729) );
  OAI21_X1 inst1_U707 ( .B1(inst1_n952), .B2(inst1_n849), .A(inst1_n728), .ZN(
        inst1_KeyArray_S31reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst1_U706 ( .B1(key1[20]), .B2(inst1_n732), .A(inst1_n727), .ZN(
        inst1_n728) );
  OAI22_X1 inst1_U705 ( .A1(inst1_n1048), .A2(inst1_n1035), .B1(inst1_n1222),
        .B2(inst1_n1237), .ZN(inst1_n727) );
  OAI21_X1 inst1_U704 ( .B1(inst1_n953), .B2(inst1_n849), .A(inst1_n726), .ZN(
        inst1_KeyArray_S31reg_gff_1_SFF_5_n6) );
  AOI21_X1 inst1_U703 ( .B1(key1[21]), .B2(inst1_n507), .A(inst1_n725), .ZN(
        inst1_n726) );
  OAI22_X1 inst1_U702 ( .A1(inst1_n1049), .A2(inst1_n1035), .B1(inst1_n997),
        .B2(inst1_n1261), .ZN(inst1_n725) );
  OAI21_X1 inst1_U701 ( .B1(inst1_n954), .B2(inst1_n849), .A(inst1_n724), .ZN(
        inst1_KeyArray_S31reg_gff_1_SFF_6_n6) );
  AOI21_X1 inst1_U700 ( .B1(key1[22]), .B2(inst1_n732), .A(inst1_n723), .ZN(
        inst1_n724) );
  OAI22_X1 inst1_U699 ( .A1(inst1_n1050), .A2(inst1_n1035), .B1(inst1_n1222),
        .B2(inst1_n1260), .ZN(inst1_n723) );
  OAI21_X1 inst1_U698 ( .B1(inst1_n955), .B2(inst1_n849), .A(inst1_n722), .ZN(
        inst1_KeyArray_S31reg_gff_1_SFF_7_n6) );
  AOI21_X1 inst1_U697 ( .B1(key1[23]), .B2(inst1_n596), .A(inst1_n721), .ZN(
        inst1_n722) );
  OAI22_X1 inst1_U696 ( .A1(inst1_n1051), .A2(inst1_n1035), .B1(inst1_n1222),
        .B2(inst1_n1259), .ZN(inst1_n721) );
  INV_X1 inst1_U695 ( .A(inst1_n720), .ZN(inst1_n1222) );
  OAI211_X1 inst1_U694 ( .C1(inst1_n957), .C2(inst1_n740), .A(inst1_n719), .B(
        inst1_n718), .ZN(inst1_KeyArray_S32reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst1_U693 ( .A1(inst1_n827), .A2(inst1_n65), .ZN(inst1_n718) );
  AOI22_X1 inst1_U692 ( .A1(inst1_n57), .A2(inst1_n926), .B1(key1[9]), .B2(
        inst1_n1156), .ZN(inst1_n719) );
  OAI21_X1 inst1_U691 ( .B1(inst1_n876), .B2(inst1_n717), .A(inst1_n716), .ZN(
        inst1_stateArray_S10reg_gff_1_SFF_0_n5) );
  AOI22_X1 inst1_U690 ( .A1(inst1_n385), .A2(ciphertext1[88]), .B1(
        plaintext1[88]), .B2(inst1_n899), .ZN(inst1_n716) );
  OAI21_X1 inst1_U689 ( .B1(inst1_n877), .B2(inst1_n717), .A(inst1_n715), .ZN(
        inst1_stateArray_S10reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst1_U688 ( .A1(inst1_n385), .A2(ciphertext1[89]), .B1(
        plaintext1[89]), .B2(inst1_n507), .ZN(inst1_n715) );
  OAI21_X1 inst1_U687 ( .B1(inst1_n878), .B2(inst1_n717), .A(inst1_n714), .ZN(
        inst1_stateArray_S10reg_gff_1_SFF_2_n5) );
  AOI22_X1 inst1_U686 ( .A1(inst1_n385), .A2(ciphertext1[90]), .B1(
        plaintext1[90]), .B2(inst1_n710), .ZN(inst1_n714) );
  OAI21_X1 inst1_U685 ( .B1(inst1_n879), .B2(inst1_n717), .A(inst1_n713), .ZN(
        inst1_stateArray_S10reg_gff_1_SFF_3_n5) );
  AOI22_X1 inst1_U684 ( .A1(inst1_n677), .A2(ciphertext1[91]), .B1(
        plaintext1[91]), .B2(inst1_n830), .ZN(inst1_n713) );
  INV_X1 inst1_U683 ( .A(inst1_n6), .ZN(inst1_n830) );
  OAI21_X1 inst1_U682 ( .B1(inst1_n880), .B2(inst1_n717), .A(inst1_n712), .ZN(
        inst1_stateArray_S10reg_gff_1_SFF_4_n5) );
  AOI22_X1 inst1_U681 ( .A1(done1), .A2(ciphertext1[92]), .B1(plaintext1[92]),
        .B2(inst1_n732), .ZN(inst1_n712) );
  OAI21_X1 inst1_U680 ( .B1(inst1_n881), .B2(inst1_n717), .A(inst1_n711), .ZN(
        inst1_stateArray_S10reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst1_U679 ( .A1(inst1_n385), .A2(ciphertext1[93]), .B1(
        plaintext1[93]), .B2(inst1_n710), .ZN(inst1_n711) );
  OAI21_X1 inst1_U678 ( .B1(inst1_n882), .B2(inst1_n717), .A(inst1_n709), .ZN(
        inst1_stateArray_S10reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst1_U677 ( .A1(inst1_n385), .A2(ciphertext1[94]), .B1(
        plaintext1[94]), .B2(inst1_n710), .ZN(inst1_n709) );
  OAI21_X1 inst1_U676 ( .B1(inst1_n883), .B2(inst1_n717), .A(inst1_n708), .ZN(
        inst1_stateArray_S10reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst1_U675 ( .A1(inst1_n385), .A2(ciphertext1[95]), .B1(
        plaintext1[95]), .B2(inst1_n710), .ZN(inst1_n708) );
  INV_X1 inst1_U674 ( .A(inst1_n707), .ZN(inst1_n717) );
  OAI21_X1 inst1_U673 ( .B1(inst1_n876), .B2(inst1_n1145), .A(inst1_n706),
        .ZN(inst1_stateArray_S11reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst1_U672 ( .A1(inst1_n707), .A2(ciphertext1[72]), .B1(
        plaintext1[80]), .B2(inst1_n710), .ZN(inst1_n706) );
  OAI21_X1 inst1_U671 ( .B1(inst1_n877), .B2(inst1_n1135), .A(inst1_n705),
        .ZN(inst1_stateArray_S11reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U670 ( .A1(inst1_n707), .A2(ciphertext1[73]), .B1(
        plaintext1[81]), .B2(inst1_n710), .ZN(inst1_n705) );
  OAI21_X1 inst1_U669 ( .B1(inst1_n878), .B2(inst1_n1145), .A(inst1_n704),
        .ZN(inst1_stateArray_S11reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U668 ( .A1(inst1_n707), .A2(ciphertext1[74]), .B1(
        plaintext1[82]), .B2(inst1_n710), .ZN(inst1_n704) );
  OAI21_X1 inst1_U667 ( .B1(inst1_n879), .B2(inst1_n1135), .A(inst1_n703),
        .ZN(inst1_stateArray_S11reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U666 ( .A1(inst1_n707), .A2(ciphertext1[75]), .B1(
        plaintext1[83]), .B2(inst1_n732), .ZN(inst1_n703) );
  OAI21_X1 inst1_U665 ( .B1(inst1_n891), .B2(inst1_n1135), .A(inst1_n702),
        .ZN(inst1_stateArray_S12reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst1_U664 ( .A1(inst1_n707), .A2(ciphertext1[71]), .B1(
        plaintext1[79]), .B2(inst1_n732), .ZN(inst1_n702) );
  OAI21_X1 inst1_U663 ( .B1(inst1_n880), .B2(inst1_n1135), .A(inst1_n701),
        .ZN(inst1_stateArray_S11reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U662 ( .A1(inst1_n707), .A2(ciphertext1[76]), .B1(
        plaintext1[84]), .B2(inst1_n732), .ZN(inst1_n701) );
  OAI21_X1 inst1_U661 ( .B1(inst1_n881), .B2(inst1_n1135), .A(inst1_n700),
        .ZN(inst1_stateArray_S11reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst1_U660 ( .A1(inst1_n707), .A2(ciphertext1[77]), .B1(
        plaintext1[85]), .B2(inst1_n710), .ZN(inst1_n700) );
  OAI21_X1 inst1_U659 ( .B1(inst1_n882), .B2(inst1_n1135), .A(inst1_n699),
        .ZN(inst1_stateArray_S11reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst1_U658 ( .A1(inst1_n707), .A2(ciphertext1[78]), .B1(
        plaintext1[86]), .B2(inst1_n732), .ZN(inst1_n699) );
  OAI21_X1 inst1_U657 ( .B1(inst1_n883), .B2(inst1_n1135), .A(inst1_n698),
        .ZN(inst1_stateArray_S11reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst1_U656 ( .A1(inst1_n707), .A2(ciphertext1[79]), .B1(
        plaintext1[87]), .B2(inst1_n732), .ZN(inst1_n698) );
  OAI21_X1 inst1_U655 ( .B1(inst1_n884), .B2(inst1_n1135), .A(inst1_n697),
        .ZN(inst1_stateArray_S12reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst1_U654 ( .A1(inst1_n707), .A2(ciphertext1[64]), .B1(
        plaintext1[72]), .B2(inst1_n710), .ZN(inst1_n697) );
  OAI21_X1 inst1_U653 ( .B1(inst1_n885), .B2(inst1_n1135), .A(inst1_n696),
        .ZN(inst1_stateArray_S12reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U652 ( .A1(inst1_n707), .A2(ciphertext1[65]), .B1(
        plaintext1[73]), .B2(inst1_n710), .ZN(inst1_n696) );
  OAI21_X1 inst1_U651 ( .B1(inst1_n886), .B2(inst1_n1135), .A(inst1_n695),
        .ZN(inst1_stateArray_S12reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U650 ( .A1(inst1_n707), .A2(ciphertext1[66]), .B1(
        plaintext1[74]), .B2(inst1_n732), .ZN(inst1_n695) );
  OAI21_X1 inst1_U649 ( .B1(inst1_n887), .B2(inst1_n1135), .A(inst1_n694),
        .ZN(inst1_stateArray_S12reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U648 ( .A1(inst1_n707), .A2(ciphertext1[67]), .B1(
        plaintext1[75]), .B2(inst1_n710), .ZN(inst1_n694) );
  OAI21_X1 inst1_U647 ( .B1(inst1_n888), .B2(inst1_n1135), .A(inst1_n693),
        .ZN(inst1_stateArray_S12reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U646 ( .A1(inst1_n707), .A2(ciphertext1[68]), .B1(
        plaintext1[76]), .B2(inst1_n732), .ZN(inst1_n693) );
  OAI21_X1 inst1_U645 ( .B1(inst1_n889), .B2(inst1_n1135), .A(inst1_n692),
        .ZN(inst1_stateArray_S12reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst1_U644 ( .A1(inst1_n707), .A2(ciphertext1[69]), .B1(
        plaintext1[77]), .B2(inst1_n710), .ZN(inst1_n692) );
  OAI21_X1 inst1_U643 ( .B1(inst1_n890), .B2(inst1_n1135), .A(inst1_n691),
        .ZN(inst1_stateArray_S12reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst1_U642 ( .A1(inst1_n707), .A2(ciphertext1[70]), .B1(
        plaintext1[78]), .B2(inst1_n732), .ZN(inst1_n691) );
  INV_X1 inst1_U641 ( .A(inst1_n6), .ZN(inst1_n732) );
  NOR2_X2 inst1_U640 ( .A1(inst1_n677), .A2(inst1_n1156), .ZN(inst1_n707) );
  OAI211_X1 inst1_U639 ( .C1(inst1_n965), .C2(inst1_n740), .A(inst1_n690), .B(
        inst1_n689), .ZN(inst1_KeyArray_S33reg_gff_1_SFF_1_n5) );
  NAND2_X1 inst1_U638 ( .A1(inst1_n1031), .A2(inst1_n57), .ZN(inst1_n689) );
  AOI22_X1 inst1_U637 ( .A1(inst1_n926), .A2(inst1_n1241), .B1(key1[1]), .B2(
        inst1_n710), .ZN(inst1_n690) );
  INV_X1 inst1_U636 ( .A(inst1_n6), .ZN(inst1_n710) );
  OAI21_X1 inst1_U635 ( .B1(inst1_n966), .B2(inst1_n849), .A(inst1_n688), .ZN(
        inst1_KeyArray_S33reg_gff_1_SFF_2_n5) );
  AOI21_X1 inst1_U634 ( .B1(key1[2]), .B2(inst1_n899), .A(inst1_n687), .ZN(
        inst1_n688) );
  OAI22_X1 inst1_U633 ( .A1(inst1_n1087), .A2(inst1_n1035), .B1(inst1_n1054),
        .B2(inst1_n997), .ZN(inst1_n687) );
  OAI21_X1 inst1_U632 ( .B1(inst1_n967), .B2(inst1_n686), .A(inst1_n685), .ZN(
        inst1_KeyArray_S33reg_gff_1_SFF_3_n5) );
  AOI21_X1 inst1_U631 ( .B1(key1[3]), .B2(inst1_n494), .A(inst1_n684), .ZN(
        inst1_n685) );
  OAI22_X1 inst1_U630 ( .A1(inst1_n1088), .A2(inst1_n1035), .B1(inst1_n1055),
        .B2(inst1_n997), .ZN(inst1_n684) );
  OAI211_X1 inst1_U629 ( .C1(inst1_n938), .C2(inst1_n1198), .A(inst1_n683),
        .B(inst1_n682), .ZN(inst1_stateArray_S31reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst1_U628 ( .A1(plaintext1[22]), .A2(inst1_n830), .ZN(inst1_n682)
         );
  AOI22_X1 inst1_U627 ( .A1(ciphertext1[22]), .A2(done1), .B1(inst1_n1217),
        .B2(ciphertext1[30]), .ZN(inst1_n683) );
  OAI211_X1 inst1_U626 ( .C1(inst1_n939), .C2(inst1_n1198), .A(inst1_n681),
        .B(inst1_n680), .ZN(inst1_stateArray_S31reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst1_U625 ( .A1(plaintext1[23]), .A2(inst1_n1156), .ZN(inst1_n680)
         );
  AOI22_X1 inst1_U624 ( .A1(done1), .A2(ciphertext1[23]), .B1(inst1_n1217),
        .B2(ciphertext1[31]), .ZN(inst1_n681) );
  OAI21_X1 inst1_U623 ( .B1(inst1_n921), .B2(inst1_n1198), .A(inst1_n679),
        .ZN(inst1_stateArray_S22reg_gff_1_SFF_5_n6) );
  AOI21_X1 inst1_U622 ( .B1(plaintext1[45]), .B2(inst1_n899), .A(inst1_n678),
        .ZN(inst1_n679) );
  OAI22_X1 inst1_U621 ( .A1(inst1_n913), .A2(inst1_n1145), .B1(inst1_n1182),
        .B2(inst1_n1249), .ZN(inst1_n678) );
  INV_X1 inst1_U620 ( .A(inst1_n677), .ZN(inst1_n1145) );
  INV_X1 inst1_U619 ( .A(inst1_n1135), .ZN(inst1_n677) );
  OAI21_X1 inst1_U618 ( .B1(inst1_n964), .B2(inst1_n849), .A(inst1_n676), .ZN(
        inst1_KeyArray_S33reg_gff_1_SFF_0_n5) );
  AOI21_X1 inst1_U617 ( .B1(key1[0]), .B2(inst1_n507), .A(inst1_n675), .ZN(
        inst1_n676) );
  OAI22_X1 inst1_U616 ( .A1(inst1_n1085), .A2(inst1_n1035), .B1(inst1_n1052),
        .B2(inst1_n997), .ZN(inst1_n675) );
  OAI21_X1 inst1_U615 ( .B1(inst1_n968), .B2(inst1_n849), .A(inst1_n674), .ZN(
        inst1_KeyArray_S33reg_gff_1_SFF_4_n5) );
  AOI21_X1 inst1_U614 ( .B1(key1[4]), .B2(inst1_n522), .A(inst1_n673), .ZN(
        inst1_n674) );
  OAI22_X1 inst1_U613 ( .A1(inst1_n1089), .A2(inst1_n1035), .B1(inst1_n1056),
        .B2(inst1_n997), .ZN(inst1_n673) );
  OAI21_X1 inst1_U612 ( .B1(inst1_n969), .B2(inst1_n686), .A(inst1_n672), .ZN(
        inst1_KeyArray_S33reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst1_U611 ( .B1(key1[5]), .B2(inst1_n494), .A(inst1_n671), .ZN(
        inst1_n672) );
  OAI22_X1 inst1_U610 ( .A1(inst1_n1084), .A2(inst1_n1035), .B1(inst1_n1057),
        .B2(inst1_n997), .ZN(inst1_n671) );
  OAI21_X1 inst1_U609 ( .B1(inst1_n970), .B2(inst1_n686), .A(inst1_n670), .ZN(
        inst1_KeyArray_S33reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst1_U608 ( .B1(key1[6]), .B2(inst1_n710), .A(inst1_n669), .ZN(
        inst1_n670) );
  OAI22_X1 inst1_U607 ( .A1(inst1_n1090), .A2(inst1_n1035), .B1(inst1_n1058),
        .B2(inst1_n997), .ZN(inst1_n669) );
  OAI21_X1 inst1_U606 ( .B1(inst1_n971), .B2(inst1_n686), .A(inst1_n668), .ZN(
        inst1_KeyArray_S33reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst1_U605 ( .B1(key1[7]), .B2(inst1_n507), .A(inst1_n667), .ZN(
        inst1_n668) );
  OAI22_X1 inst1_U604 ( .A1(inst1_n1091), .A2(inst1_n1035), .B1(inst1_n1059),
        .B2(inst1_n1222), .ZN(inst1_n667) );
  OAI211_X1 inst1_U603 ( .C1(inst1_n1102), .C2(inst1_n666), .A(inst1_n665),
        .B(inst1_n664), .ZN(inst1_stateArray_S03reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst1_U602 ( .A1(inst1_n926), .A2(ciphertext1[88]), .B1(inst1_n663),
        .B2(inst1_n662), .ZN(inst1_n664) );
  XNOR2_X1 inst1_U601 ( .A(inst1_n1209), .B(inst1_n661), .ZN(inst1_n662) );
  AOI22_X1 inst1_U600 ( .A1(inst1_n660), .A2(ciphertext1[88]), .B1(inst1_n1103), .B2(inst1_n659), .ZN(inst1_n661) );
  AOI22_X1 inst1_U599 ( .A1(inst1_n827), .A2(ciphertext1[96]), .B1(
        plaintext1[96]), .B2(inst1_n1228), .ZN(inst1_n665) );
  OAI211_X1 inst1_U598 ( .C1(inst1_n972), .C2(inst1_n740), .A(inst1_n658), .B(
        inst1_n657), .ZN(inst1_KeyArray_S00reg_gff_1_SFF_0_n6) );
  OAI21_X1 inst1_U597 ( .B1(inst1_n948), .B2(inst1_n656), .A(inst1_n655), .ZN(
        inst1_n657) );
  AOI21_X1 inst1_U596 ( .B1(inst1_n948), .B2(inst1_n656), .A(inst1_n1203),
        .ZN(inst1_n655) );
  NAND2_X1 inst1_U595 ( .A1(inst1_n654), .A2(inst1_n1248), .ZN(inst1_n656) );
  AOI22_X1 inst1_U594 ( .A1(inst1_n827), .A2(inst1_n1248), .B1(key1[120]),
        .B2(inst1_n1228), .ZN(inst1_n658) );
  OAI211_X1 inst1_U593 ( .C1(inst1_n973), .C2(inst1_n740), .A(inst1_n653), .B(
        inst1_n652), .ZN(inst1_KeyArray_S00reg_gff_1_SFF_1_n6) );
  OAI21_X1 inst1_U592 ( .B1(inst1_n949), .B2(inst1_n651), .A(inst1_n650), .ZN(
        inst1_n652) );
  AOI21_X1 inst1_U591 ( .B1(inst1_n949), .B2(inst1_n651), .A(inst1_n1203),
        .ZN(inst1_n650) );
  NAND2_X1 inst1_U590 ( .A1(inst1_n654), .A2(inst1_n1241), .ZN(inst1_n651) );
  AOI22_X1 inst1_U589 ( .A1(inst1_n827), .A2(inst1_n1241), .B1(key1[121]),
        .B2(inst1_n1228), .ZN(inst1_n653) );
  OAI211_X1 inst1_U588 ( .C1(inst1_n974), .C2(inst1_n740), .A(inst1_n649), .B(
        inst1_n648), .ZN(inst1_KeyArray_S00reg_gff_1_SFF_2_n6) );
  OAI21_X1 inst1_U587 ( .B1(inst1_n950), .B2(inst1_n647), .A(inst1_n646), .ZN(
        inst1_n648) );
  AOI21_X1 inst1_U586 ( .B1(inst1_n950), .B2(inst1_n647), .A(inst1_n1015),
        .ZN(inst1_n646) );
  NAND2_X1 inst1_U585 ( .A1(inst1_n654), .A2(inst1_n1242), .ZN(inst1_n647) );
  AOI22_X1 inst1_U584 ( .A1(inst1_n827), .A2(inst1_n1242), .B1(key1[122]),
        .B2(inst1_n1228), .ZN(inst1_n649) );
  OAI211_X1 inst1_U583 ( .C1(inst1_n975), .C2(inst1_n740), .A(inst1_n645), .B(
        inst1_n644), .ZN(inst1_KeyArray_S00reg_gff_1_SFF_3_n6) );
  OAI21_X1 inst1_U582 ( .B1(inst1_n951), .B2(inst1_n643), .A(inst1_n642), .ZN(
        inst1_n644) );
  AOI21_X1 inst1_U581 ( .B1(inst1_n951), .B2(inst1_n643), .A(inst1_n1015),
        .ZN(inst1_n642) );
  NAND2_X1 inst1_U580 ( .A1(inst1_n654), .A2(inst1_n1247), .ZN(inst1_n643) );
  AOI22_X1 inst1_U579 ( .A1(inst1_n827), .A2(inst1_n1247), .B1(key1[123]),
        .B2(inst1_n1228), .ZN(inst1_n645) );
  OAI211_X1 inst1_U578 ( .C1(inst1_n976), .C2(inst1_n740), .A(inst1_n641), .B(
        inst1_n640), .ZN(inst1_KeyArray_S00reg_gff_1_SFF_4_n6) );
  OAI21_X1 inst1_U577 ( .B1(inst1_n952), .B2(inst1_n639), .A(inst1_n638), .ZN(
        inst1_n640) );
  AOI21_X1 inst1_U576 ( .B1(inst1_n952), .B2(inst1_n639), .A(inst1_n1203),
        .ZN(inst1_n638) );
  NAND2_X1 inst1_U575 ( .A1(inst1_n654), .A2(inst1_n1246), .ZN(inst1_n639) );
  AOI22_X1 inst1_U574 ( .A1(inst1_n827), .A2(inst1_n1246), .B1(key1[124]),
        .B2(inst1_n1228), .ZN(inst1_n641) );
  OAI211_X1 inst1_U573 ( .C1(inst1_n977), .C2(inst1_n740), .A(inst1_n637), .B(
        inst1_n636), .ZN(inst1_KeyArray_S00reg_gff_1_SFF_5_n6) );
  OAI21_X1 inst1_U572 ( .B1(inst1_n953), .B2(inst1_n635), .A(inst1_n634), .ZN(
        inst1_n636) );
  AOI21_X1 inst1_U571 ( .B1(inst1_n953), .B2(inst1_n635), .A(inst1_n1015),
        .ZN(inst1_n634) );
  NAND2_X1 inst1_U570 ( .A1(inst1_n654), .A2(inst1_n1245), .ZN(inst1_n635) );
  AOI22_X1 inst1_U569 ( .A1(inst1_n827), .A2(inst1_n1245), .B1(key1[125]),
        .B2(inst1_n1228), .ZN(inst1_n637) );
  OAI211_X1 inst1_U568 ( .C1(inst1_n978), .C2(inst1_n740), .A(inst1_n633), .B(
        inst1_n632), .ZN(inst1_KeyArray_S00reg_gff_1_SFF_6_n6) );
  OAI21_X1 inst1_U567 ( .B1(inst1_n954), .B2(inst1_n631), .A(inst1_n630), .ZN(
        inst1_n632) );
  AOI21_X1 inst1_U566 ( .B1(inst1_n954), .B2(inst1_n631), .A(inst1_n1203),
        .ZN(inst1_n630) );
  NAND2_X1 inst1_U565 ( .A1(inst1_n654), .A2(inst1_n1244), .ZN(inst1_n631) );
  AOI22_X1 inst1_U564 ( .A1(inst1_n827), .A2(inst1_n1244), .B1(key1[126]),
        .B2(inst1_n1228), .ZN(inst1_n633) );
  OAI211_X1 inst1_U563 ( .C1(inst1_n979), .C2(inst1_n740), .A(inst1_n629), .B(
        inst1_n628), .ZN(inst1_KeyArray_S00reg_gff_1_SFF_7_n6) );
  OAI21_X1 inst1_U562 ( .B1(inst1_n955), .B2(inst1_n627), .A(inst1_n626), .ZN(
        inst1_n628) );
  AOI21_X1 inst1_U561 ( .B1(inst1_n955), .B2(inst1_n627), .A(inst1_n1015),
        .ZN(inst1_n626) );
  NAND2_X1 inst1_U560 ( .A1(inst1_n654), .A2(inst1_n1243), .ZN(inst1_n627) );
  AOI22_X1 inst1_U559 ( .A1(inst1_n625), .A2(inst1_n624), .B1(inst1_n1077),
        .B2(inst1_n1236), .ZN(inst1_n654) );
  AND4_X1 inst1_U558 ( .A1(inst1_n1226), .A2(inst1_n1240), .A3(inst1_n1264),
        .A4(inst1_n1071), .ZN(inst1_n624) );
  AND4_X1 inst1_U557 ( .A1(inst1_n1263), .A2(inst1_n1074), .A3(inst1_n1060),
        .A4(inst1_n1061), .ZN(inst1_n625) );
  AOI22_X1 inst1_U556 ( .A1(inst1_n827), .A2(inst1_n1243), .B1(key1[127]),
        .B2(inst1_n1228), .ZN(inst1_n629) );
  OAI211_X1 inst1_U555 ( .C1(inst1_n935), .C2(inst1_n1198), .A(inst1_n623),
        .B(inst1_n622), .ZN(inst1_stateArray_S31reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst1_U554 ( .A1(plaintext1[19]), .A2(inst1_n1156), .ZN(inst1_n622)
         );
  AOI22_X1 inst1_U553 ( .A1(inst1_n677), .A2(ciphertext1[19]), .B1(inst1_n1217), .B2(ciphertext1[27]), .ZN(inst1_n623) );
  OAI211_X1 inst1_U552 ( .C1(inst1_n1114), .C2(inst1_n666), .A(inst1_n621),
        .B(inst1_n620), .ZN(inst1_stateArray_S03reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U551 ( .A1(inst1_n926), .A2(ciphertext1[89]), .B1(inst1_n663),
        .B2(inst1_n619), .ZN(inst1_n620) );
  XNOR2_X1 inst1_U550 ( .A(inst1_n618), .B(inst1_n617), .ZN(inst1_n619) );
  AOI22_X1 inst1_U549 ( .A1(inst1_n660), .A2(inst1_n1115), .B1(ciphertext1[89]), .B2(inst1_n659), .ZN(inst1_n617) );
  XNOR2_X1 inst1_U548 ( .A(inst1_n616), .B(inst1_n1202), .ZN(inst1_n618) );
  AOI22_X1 inst1_U547 ( .A1(inst1_n827), .A2(ciphertext1[97]), .B1(
        plaintext1[97]), .B2(inst1_n1228), .ZN(inst1_n621) );
  INV_X1 inst1_U546 ( .A(inst1_n997), .ZN(inst1_n827) );
  OAI211_X1 inst1_U545 ( .C1(inst1_n1110), .C2(inst1_n666), .A(inst1_n615),
        .B(inst1_n614), .ZN(inst1_stateArray_S03reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U544 ( .A1(ciphertext1[91]), .A2(inst1_n926), .B1(inst1_n663),
        .B2(inst1_n613), .ZN(inst1_n614) );
  XNOR2_X1 inst1_U543 ( .A(ciphertext1[91]), .B(inst1_n612), .ZN(inst1_n613)
         );
  XNOR2_X1 inst1_U542 ( .A(inst1_n611), .B(inst1_n610), .ZN(inst1_n612) );
  AOI22_X1 inst1_U541 ( .A1(inst1_n660), .A2(inst1_n1187), .B1(inst1_n1186),
        .B2(inst1_n659), .ZN(inst1_n610) );
  INV_X1 inst1_U540 ( .A(inst1_n1187), .ZN(inst1_n1186) );
  AOI22_X1 inst1_U539 ( .A1(ciphertext1[122]), .A2(inst1_n1118), .B1(
        ciphertext1[90]), .B2(inst1_n1227), .ZN(inst1_n611) );
  AOI22_X1 inst1_U538 ( .A1(inst1_n859), .A2(ciphertext1[99]), .B1(
        plaintext1[99]), .B2(inst1_n1228), .ZN(inst1_n615) );
  OAI211_X1 inst1_U537 ( .C1(inst1_n1096), .C2(inst1_n666), .A(inst1_n609),
        .B(inst1_n608), .ZN(inst1_stateArray_S03reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst1_U536 ( .A1(inst1_n926), .A2(ciphertext1[94]), .B1(inst1_n663),
        .B2(inst1_n607), .ZN(inst1_n608) );
  XNOR2_X1 inst1_U535 ( .A(inst1_n606), .B(inst1_n605), .ZN(inst1_n607) );
  AOI22_X1 inst1_U534 ( .A1(inst1_n1098), .A2(ciphertext1[30]), .B1(
        inst1_n1097), .B2(ciphertext1[125]), .ZN(inst1_n605) );
  AOI22_X1 inst1_U533 ( .A1(inst1_n604), .A2(inst1_n1122), .B1(ciphertext1[93]), .B2(inst1_n603), .ZN(inst1_n606) );
  INV_X1 inst1_U532 ( .A(inst1_n604), .ZN(inst1_n603) );
  INV_X1 inst1_U531 ( .A(inst1_n1015), .ZN(inst1_n926) );
  AOI22_X1 inst1_U530 ( .A1(inst1_n859), .A2(ciphertext1[102]), .B1(
        plaintext1[102]), .B2(inst1_n1228), .ZN(inst1_n609) );
  OAI211_X1 inst1_U529 ( .C1(inst1_n1227), .C2(inst1_n666), .A(inst1_n602),
        .B(inst1_n601), .ZN(inst1_stateArray_S03reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U528 ( .A1(inst1_n822), .A2(ciphertext1[90]), .B1(inst1_n663),
        .B2(inst1_n600), .ZN(inst1_n601) );
  XNOR2_X1 inst1_U527 ( .A(inst1_n599), .B(inst1_n598), .ZN(inst1_n600) );
  AOI22_X1 inst1_U526 ( .A1(inst1_n1109), .A2(inst1_n1210), .B1(inst1_n597),
        .B2(ciphertext1[26]), .ZN(inst1_n598) );
  INV_X1 inst1_U525 ( .A(inst1_n1210), .ZN(inst1_n597) );
  AOI22_X1 inst1_U524 ( .A1(inst1_n859), .A2(ciphertext1[98]), .B1(
        plaintext1[98]), .B2(inst1_n596), .ZN(inst1_n602) );
  OAI211_X1 inst1_U523 ( .C1(inst1_n1098), .C2(inst1_n666), .A(inst1_n595),
        .B(inst1_n594), .ZN(inst1_stateArray_S03reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst1_U522 ( .A1(inst1_n822), .A2(ciphertext1[93]), .B1(inst1_n663),
        .B2(inst1_n593), .ZN(inst1_n594) );
  XNOR2_X1 inst1_U521 ( .A(inst1_n592), .B(inst1_n591), .ZN(inst1_n593) );
  AOI22_X1 inst1_U520 ( .A1(ciphertext1[124]), .A2(inst1_n1229), .B1(
        ciphertext1[29]), .B2(inst1_n1225), .ZN(inst1_n591) );
  AOI22_X1 inst1_U519 ( .A1(inst1_n1100), .A2(inst1_n590), .B1(inst1_n589),
        .B2(ciphertext1[92]), .ZN(inst1_n592) );
  INV_X1 inst1_U518 ( .A(inst1_n590), .ZN(inst1_n589) );
  AOI22_X1 inst1_U517 ( .A1(inst1_n859), .A2(ciphertext1[101]), .B1(
        plaintext1[101]), .B2(inst1_n596), .ZN(inst1_n595) );
  OAI211_X1 inst1_U516 ( .C1(inst1_n1225), .C2(inst1_n666), .A(inst1_n588),
        .B(inst1_n587), .ZN(inst1_stateArray_S03reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U515 ( .A1(inst1_n822), .A2(ciphertext1[92]), .B1(inst1_n663),
        .B2(inst1_n586), .ZN(inst1_n587) );
  XNOR2_X1 inst1_U514 ( .A(inst1_n585), .B(inst1_n584), .ZN(inst1_n586) );
  AOI22_X1 inst1_U513 ( .A1(inst1_n1105), .A2(inst1_n583), .B1(inst1_n582),
        .B2(ciphertext1[28]), .ZN(inst1_n584) );
  INV_X1 inst1_U512 ( .A(inst1_n582), .ZN(inst1_n583) );
  AOI22_X1 inst1_U511 ( .A1(inst1_n581), .A2(inst1_n660), .B1(inst1_n659),
        .B2(inst1_n580), .ZN(inst1_n585) );
  AOI22_X1 inst1_U510 ( .A1(inst1_n859), .A2(ciphertext1[100]), .B1(
        plaintext1[100]), .B2(inst1_n596), .ZN(inst1_n588) );
  OAI211_X1 inst1_U509 ( .C1(inst1_n933), .C2(inst1_n1198), .A(inst1_n579),
        .B(inst1_n578), .ZN(inst1_stateArray_S31reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst1_U508 ( .A1(plaintext1[17]), .A2(inst1_n1156), .ZN(inst1_n578)
         );
  AOI22_X1 inst1_U507 ( .A1(done1), .A2(ciphertext1[17]), .B1(inst1_n1217),
        .B2(ciphertext1[25]), .ZN(inst1_n579) );
  OAI211_X1 inst1_U506 ( .C1(inst1_n932), .C2(inst1_n1198), .A(inst1_n577),
        .B(inst1_n576), .ZN(inst1_stateArray_S31reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst1_U505 ( .A1(plaintext1[16]), .A2(inst1_n1156), .ZN(inst1_n576)
         );
  AOI22_X1 inst1_U504 ( .A1(inst1_n677), .A2(ciphertext1[16]), .B1(inst1_n1217), .B2(ciphertext1[24]), .ZN(inst1_n577) );
  OAI211_X1 inst1_U503 ( .C1(inst1_n1094), .C2(inst1_n666), .A(inst1_n575),
        .B(inst1_n574), .ZN(inst1_stateArray_S03reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst1_U502 ( .A1(inst1_n822), .A2(ciphertext1[95]), .B1(inst1_n663),
        .B2(inst1_n573), .ZN(inst1_n574) );
  XNOR2_X1 inst1_U501 ( .A(inst1_n572), .B(inst1_n571), .ZN(inst1_n573) );
  AOI22_X1 inst1_U500 ( .A1(inst1_n1096), .A2(ciphertext1[94]), .B1(
        inst1_n1106), .B2(ciphertext1[126]), .ZN(inst1_n571) );
  AOI22_X1 inst1_U499 ( .A1(inst1_n1092), .A2(inst1_n1212), .B1(inst1_n1211),
        .B2(ciphertext1[95]), .ZN(inst1_n572) );
  AOI22_X1 inst1_U498 ( .A1(inst1_n859), .A2(ciphertext1[103]), .B1(
        plaintext1[103]), .B2(inst1_n596), .ZN(inst1_n575) );
  INV_X1 inst1_U497 ( .A(inst1_n997), .ZN(inst1_n859) );
  OAI211_X1 inst1_U496 ( .C1(inst1_n934), .C2(inst1_n1198), .A(inst1_n570),
        .B(inst1_n569), .ZN(inst1_stateArray_S31reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst1_U495 ( .A1(plaintext1[18]), .A2(inst1_n507), .ZN(inst1_n569)
         );
  AOI22_X1 inst1_U494 ( .A1(done1), .A2(ciphertext1[18]), .B1(inst1_n1217),
        .B2(ciphertext1[26]), .ZN(inst1_n570) );
  OAI211_X1 inst1_U493 ( .C1(inst1_n936), .C2(inst1_n1198), .A(inst1_n568),
        .B(inst1_n567), .ZN(inst1_stateArray_S31reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst1_U492 ( .A1(plaintext1[20]), .A2(inst1_n1156), .ZN(inst1_n567)
         );
  AOI22_X1 inst1_U491 ( .A1(inst1_n677), .A2(ciphertext1[20]), .B1(inst1_n1217), .B2(ciphertext1[28]), .ZN(inst1_n568) );
  OAI211_X1 inst1_U490 ( .C1(inst1_n1220), .C2(inst1_n566), .A(inst1_n565),
        .B(inst1_n564), .ZN(inst1_stateArray_S13reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst1_U489 ( .A1(inst1_n822), .A2(ciphertext1[56]), .B1(
        ciphertext1[88]), .B2(inst1_n563), .ZN(inst1_n564) );
  AOI22_X1 inst1_U488 ( .A1(inst1_n677), .A2(ciphertext1[64]), .B1(
        plaintext1[64]), .B2(inst1_n596), .ZN(inst1_n565) );
  XNOR2_X1 inst1_U487 ( .A(inst1_n1209), .B(inst1_n562), .ZN(inst1_n566) );
  AOI22_X1 inst1_U486 ( .A1(inst1_n1102), .A2(inst1_n561), .B1(inst1_n560),
        .B2(ciphertext1[120]), .ZN(inst1_n562) );
  AOI22_X1 inst1_U485 ( .A1(inst1_n1113), .A2(ciphertext1[56]), .B1(
        inst1_n1233), .B2(ciphertext1[24]), .ZN(inst1_n1209) );
  OAI211_X1 inst1_U484 ( .C1(inst1_n559), .C2(inst1_n1207), .A(inst1_n558),
        .B(inst1_n557), .ZN(inst1_stateArray_S13reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U483 ( .A1(inst1_n822), .A2(ciphertext1[57]), .B1(
        ciphertext1[89]), .B2(inst1_n563), .ZN(inst1_n557) );
  AOI22_X1 inst1_U482 ( .A1(done1), .A2(ciphertext1[65]), .B1(plaintext1[65]),
        .B2(inst1_n596), .ZN(inst1_n558) );
  XNOR2_X1 inst1_U481 ( .A(inst1_n556), .B(inst1_n555), .ZN(inst1_n559) );
  AOI22_X1 inst1_U480 ( .A1(inst1_n1103), .A2(inst1_n561), .B1(inst1_n560),
        .B2(ciphertext1[88]), .ZN(inst1_n555) );
  XNOR2_X1 inst1_U479 ( .A(inst1_n1202), .B(inst1_n554), .ZN(inst1_n556) );
  AOI22_X1 inst1_U478 ( .A1(inst1_n1114), .A2(ciphertext1[56]), .B1(
        inst1_n1233), .B2(ciphertext1[121]), .ZN(inst1_n554) );
  AOI22_X1 inst1_U477 ( .A1(inst1_n1121), .A2(ciphertext1[57]), .B1(
        inst1_n1235), .B2(ciphertext1[25]), .ZN(inst1_n1202) );
  OAI211_X1 inst1_U476 ( .C1(inst1_n553), .C2(inst1_n1207), .A(inst1_n552),
        .B(inst1_n551), .ZN(inst1_stateArray_S13reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U475 ( .A1(inst1_n822), .A2(ciphertext1[58]), .B1(
        ciphertext1[90]), .B2(inst1_n563), .ZN(inst1_n551) );
  AOI22_X1 inst1_U474 ( .A1(inst1_n677), .A2(ciphertext1[66]), .B1(
        plaintext1[66]), .B2(inst1_n596), .ZN(inst1_n552) );
  XNOR2_X1 inst1_U473 ( .A(inst1_n550), .B(inst1_n549), .ZN(inst1_n553) );
  AOI22_X1 inst1_U472 ( .A1(inst1_n1200), .A2(ciphertext1[58]), .B1(
        inst1_n1119), .B2(inst1_n1199), .ZN(inst1_n549) );
  INV_X1 inst1_U471 ( .A(inst1_n1200), .ZN(inst1_n1199) );
  AOI22_X1 inst1_U470 ( .A1(inst1_n1115), .A2(ciphertext1[57]), .B1(
        inst1_n1235), .B2(ciphertext1[89]), .ZN(inst1_n550) );
  OAI211_X1 inst1_U469 ( .C1(inst1_n1220), .C2(inst1_n548), .A(inst1_n547),
        .B(inst1_n546), .ZN(inst1_stateArray_S13reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U468 ( .A1(inst1_n822), .A2(ciphertext1[59]), .B1(
        ciphertext1[91]), .B2(inst1_n563), .ZN(inst1_n546) );
  AOI22_X1 inst1_U467 ( .A1(done1), .A2(ciphertext1[67]), .B1(plaintext1[67]),
        .B2(inst1_n596), .ZN(inst1_n547) );
  XNOR2_X1 inst1_U466 ( .A(inst1_n545), .B(inst1_n544), .ZN(inst1_n548) );
  AOI22_X1 inst1_U465 ( .A1(inst1_n1110), .A2(inst1_n560), .B1(inst1_n561),
        .B2(ciphertext1[123]), .ZN(inst1_n544) );
  INV_X1 inst1_U464 ( .A(inst1_n561), .ZN(inst1_n560) );
  XNOR2_X1 inst1_U463 ( .A(inst1_n599), .B(inst1_n1187), .ZN(inst1_n545) );
  AOI22_X1 inst1_U462 ( .A1(ciphertext1[27]), .A2(inst1_n1116), .B1(
        ciphertext1[59]), .B2(inst1_n1231), .ZN(inst1_n1187) );
  OAI211_X1 inst1_U461 ( .C1(inst1_n543), .C2(inst1_n1220), .A(inst1_n542),
        .B(inst1_n541), .ZN(inst1_stateArray_S13reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U460 ( .A1(inst1_n822), .A2(ciphertext1[60]), .B1(
        ciphertext1[92]), .B2(inst1_n563), .ZN(inst1_n541) );
  AOI22_X1 inst1_U459 ( .A1(done1), .A2(ciphertext1[68]), .B1(plaintext1[68]),
        .B2(inst1_n596), .ZN(inst1_n542) );
  XNOR2_X1 inst1_U458 ( .A(inst1_n540), .B(inst1_n539), .ZN(inst1_n543) );
  AOI22_X1 inst1_U457 ( .A1(inst1_n1111), .A2(inst1_n1191), .B1(inst1_n1190),
        .B2(ciphertext1[91]), .ZN(inst1_n539) );
  INV_X1 inst1_U456 ( .A(inst1_n1191), .ZN(inst1_n1190) );
  XNOR2_X1 inst1_U455 ( .A(inst1_n561), .B(inst1_n538), .ZN(inst1_n540) );
  AOI22_X1 inst1_U454 ( .A1(ciphertext1[60]), .A2(inst1_n1116), .B1(
        ciphertext1[59]), .B2(inst1_n1234), .ZN(inst1_n538) );
  AOI22_X1 inst1_U453 ( .A1(inst1_n1093), .A2(inst1_n1092), .B1(
        ciphertext1[95]), .B2(ciphertext1[63]), .ZN(inst1_n561) );
  OAI211_X1 inst1_U452 ( .C1(inst1_n1220), .C2(inst1_n537), .A(inst1_n536),
        .B(inst1_n535), .ZN(inst1_stateArray_S13reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst1_U451 ( .A1(inst1_n822), .A2(ciphertext1[61]), .B1(
        ciphertext1[93]), .B2(inst1_n563), .ZN(inst1_n535) );
  AOI22_X1 inst1_U450 ( .A1(done1), .A2(ciphertext1[69]), .B1(plaintext1[69]),
        .B2(inst1_n596), .ZN(inst1_n536) );
  XNOR2_X1 inst1_U449 ( .A(inst1_n582), .B(inst1_n534), .ZN(inst1_n537) );
  AOI22_X1 inst1_U448 ( .A1(inst1_n533), .A2(ciphertext1[61]), .B1(inst1_n1249), .B2(inst1_n532), .ZN(inst1_n534) );
  OAI211_X1 inst1_U447 ( .C1(inst1_n531), .C2(inst1_n1220), .A(inst1_n530),
        .B(inst1_n529), .ZN(inst1_stateArray_S13reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst1_U446 ( .A1(inst1_n822), .A2(ciphertext1[62]), .B1(
        ciphertext1[94]), .B2(inst1_n563), .ZN(inst1_n529) );
  AOI22_X1 inst1_U445 ( .A1(inst1_n677), .A2(ciphertext1[70]), .B1(
        plaintext1[70]), .B2(inst1_n596), .ZN(inst1_n530) );
  XNOR2_X1 inst1_U444 ( .A(inst1_n590), .B(inst1_n528), .ZN(inst1_n531) );
  AOI22_X1 inst1_U443 ( .A1(ciphertext1[62]), .A2(inst1_n527), .B1(inst1_n526),
        .B2(inst1_n1232), .ZN(inst1_n528) );
  OAI211_X1 inst1_U442 ( .C1(inst1_n525), .C2(inst1_n1220), .A(inst1_n524),
        .B(inst1_n523), .ZN(inst1_stateArray_S13reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst1_U441 ( .A1(inst1_n822), .A2(ciphertext1[63]), .B1(
        ciphertext1[95]), .B2(inst1_n563), .ZN(inst1_n523) );
  NAND2_X1 inst1_U440 ( .A1(inst1_n1215), .A2(inst1_n1185), .ZN(inst1_n563) );
  INV_X1 inst1_U439 ( .A(inst1_n1015), .ZN(inst1_n822) );
  AOI22_X1 inst1_U438 ( .A1(done1), .A2(ciphertext1[71]), .B1(plaintext1[71]),
        .B2(inst1_n522), .ZN(inst1_n524) );
  XNOR2_X1 inst1_U437 ( .A(inst1_n604), .B(inst1_n521), .ZN(inst1_n525) );
  AOI22_X1 inst1_U436 ( .A1(inst1_n1094), .A2(inst1_n1211), .B1(inst1_n1212),
        .B2(ciphertext1[127]), .ZN(inst1_n521) );
  OAI211_X1 inst1_U435 ( .C1(inst1_n1217), .C2(inst1_n1075), .A(inst1_n6), .B(
        inst1_n520), .ZN(inst1_calcRCon_n51) );
  NAND2_X1 inst1_U434 ( .A1(inst1_n1217), .A2(inst1_n1226), .ZN(inst1_n520) );
  OAI221_X1 inst1_U433 ( .B1(inst1_n1217), .B2(inst1_n1073), .C1(inst1_n1185),
        .C2(inst1_n1074), .A(inst1_n6), .ZN(inst1_calcRCon_n49) );
  OAI221_X1 inst1_U432 ( .B1(inst1_n1217), .B2(inst1_n1070), .C1(inst1_n1182),
        .C2(inst1_n1071), .A(inst1_n6), .ZN(inst1_calcRCon_n44) );
  OAI21_X1 inst1_U431 ( .B1(inst1_n1102), .B2(inst1_n1006), .A(inst1_n519),
        .ZN(inst1_stateArray_S00reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst1_U430 ( .A1(ciphertext1[112]), .A2(inst1_n191), .B1(
        plaintext1[120]), .B2(inst1_n522), .ZN(inst1_n519) );
  OAI21_X1 inst1_U429 ( .B1(inst1_n1114), .B2(inst1_n1006), .A(inst1_n518),
        .ZN(inst1_stateArray_S00reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U428 ( .A1(ciphertext1[113]), .A2(inst1_n191), .B1(
        plaintext1[121]), .B2(inst1_n522), .ZN(inst1_n518) );
  OAI21_X1 inst1_U427 ( .B1(inst1_n1006), .B2(inst1_n1227), .A(inst1_n517),
        .ZN(inst1_stateArray_S00reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U426 ( .A1(ciphertext1[114]), .A2(inst1_n191), .B1(
        plaintext1[122]), .B2(inst1_n522), .ZN(inst1_n517) );
  OAI21_X1 inst1_U425 ( .B1(inst1_n1110), .B2(inst1_n1006), .A(inst1_n516),
        .ZN(inst1_stateArray_S00reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U424 ( .A1(ciphertext1[115]), .A2(inst1_n191), .B1(
        plaintext1[123]), .B2(inst1_n522), .ZN(inst1_n516) );
  OAI21_X1 inst1_U423 ( .B1(inst1_n1006), .B2(inst1_n1225), .A(inst1_n515),
        .ZN(inst1_stateArray_S00reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U422 ( .A1(ciphertext1[116]), .A2(inst1_n191), .B1(
        plaintext1[124]), .B2(inst1_n522), .ZN(inst1_n515) );
  OAI21_X1 inst1_U421 ( .B1(inst1_n1098), .B2(inst1_n1006), .A(inst1_n514),
        .ZN(inst1_stateArray_S00reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst1_U420 ( .A1(ciphertext1[117]), .A2(inst1_n191), .B1(
        plaintext1[125]), .B2(inst1_n522), .ZN(inst1_n514) );
  OAI21_X1 inst1_U419 ( .B1(inst1_n1096), .B2(inst1_n1006), .A(inst1_n513),
        .ZN(inst1_stateArray_S00reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst1_U418 ( .A1(ciphertext1[118]), .A2(inst1_n191), .B1(
        plaintext1[126]), .B2(inst1_n522), .ZN(inst1_n513) );
  OAI21_X1 inst1_U417 ( .B1(inst1_n1094), .B2(inst1_n1006), .A(inst1_n512),
        .ZN(inst1_stateArray_S00reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst1_U416 ( .A1(ciphertext1[119]), .A2(inst1_n191), .B1(
        plaintext1[127]), .B2(inst1_n522), .ZN(inst1_n512) );
  OAI21_X1 inst1_U415 ( .B1(inst1_n1006), .B2(inst1_n1279), .A(inst1_n511),
        .ZN(inst1_stateArray_S01reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst1_U414 ( .A1(ciphertext1[104]), .A2(inst1_n191), .B1(
        plaintext1[112]), .B2(inst1_n522), .ZN(inst1_n511) );
  OAI21_X1 inst1_U413 ( .B1(inst1_n1006), .B2(inst1_n1278), .A(inst1_n510),
        .ZN(inst1_stateArray_S01reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U412 ( .A1(ciphertext1[105]), .A2(inst1_n191), .B1(
        plaintext1[113]), .B2(inst1_n522), .ZN(inst1_n510) );
  OAI21_X1 inst1_U411 ( .B1(inst1_n1006), .B2(inst1_n1277), .A(inst1_n509),
        .ZN(inst1_stateArray_S01reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U410 ( .A1(ciphertext1[106]), .A2(inst1_n191), .B1(
        plaintext1[114]), .B2(inst1_n522), .ZN(inst1_n509) );
  INV_X1 inst1_U409 ( .A(inst1_n6), .ZN(inst1_n522) );
  OAI21_X1 inst1_U408 ( .B1(inst1_n1006), .B2(inst1_n1276), .A(inst1_n508),
        .ZN(inst1_stateArray_S01reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U407 ( .A1(ciphertext1[107]), .A2(inst1_n191), .B1(
        plaintext1[115]), .B2(inst1_n507), .ZN(inst1_n508) );
  OAI21_X1 inst1_U406 ( .B1(inst1_n1006), .B2(inst1_n1275), .A(inst1_n506),
        .ZN(inst1_stateArray_S01reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U405 ( .A1(ciphertext1[108]), .A2(inst1_n191), .B1(
        plaintext1[116]), .B2(inst1_n507), .ZN(inst1_n506) );
  OAI21_X1 inst1_U404 ( .B1(inst1_n1006), .B2(inst1_n1274), .A(inst1_n505),
        .ZN(inst1_stateArray_S01reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst1_U403 ( .A1(ciphertext1[109]), .A2(inst1_n191), .B1(
        plaintext1[117]), .B2(inst1_n507), .ZN(inst1_n505) );
  OAI21_X1 inst1_U402 ( .B1(inst1_n997), .B2(inst1_n1273), .A(inst1_n504),
        .ZN(inst1_stateArray_S01reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst1_U401 ( .A1(ciphertext1[110]), .A2(inst1_n191), .B1(
        plaintext1[118]), .B2(inst1_n507), .ZN(inst1_n504) );
  OAI21_X1 inst1_U400 ( .B1(inst1_n997), .B2(inst1_n1272), .A(inst1_n503),
        .ZN(inst1_stateArray_S01reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst1_U399 ( .A1(ciphertext1[111]), .A2(inst1_n191), .B1(
        plaintext1[119]), .B2(inst1_n507), .ZN(inst1_n503) );
  INV_X1 inst1_U398 ( .A(inst1_n720), .ZN(inst1_n997) );
  OAI21_X1 inst1_U397 ( .B1(inst1_n868), .B2(inst1_n1198), .A(inst1_n502),
        .ZN(inst1_stateArray_S02reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst1_U396 ( .A1(ciphertext1[104]), .A2(inst1_n827), .B1(
        plaintext1[104]), .B2(inst1_n507), .ZN(inst1_n502) );
  OAI21_X1 inst1_U395 ( .B1(inst1_n869), .B2(inst1_n1198), .A(inst1_n501),
        .ZN(inst1_stateArray_S02reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst1_U394 ( .A1(ciphertext1[105]), .A2(inst1_n819), .B1(
        plaintext1[105]), .B2(inst1_n507), .ZN(inst1_n501) );
  OAI21_X1 inst1_U393 ( .B1(inst1_n870), .B2(inst1_n1198), .A(inst1_n500),
        .ZN(inst1_stateArray_S02reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst1_U392 ( .A1(ciphertext1[106]), .A2(inst1_n819), .B1(
        plaintext1[106]), .B2(inst1_n507), .ZN(inst1_n500) );
  OAI21_X1 inst1_U391 ( .B1(inst1_n871), .B2(inst1_n1198), .A(inst1_n499),
        .ZN(inst1_stateArray_S02reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst1_U390 ( .A1(ciphertext1[107]), .A2(inst1_n819), .B1(
        plaintext1[107]), .B2(inst1_n507), .ZN(inst1_n499) );
  OAI21_X1 inst1_U389 ( .B1(inst1_n872), .B2(inst1_n1198), .A(inst1_n498),
        .ZN(inst1_stateArray_S02reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst1_U388 ( .A1(ciphertext1[108]), .A2(inst1_n720), .B1(
        plaintext1[108]), .B2(inst1_n507), .ZN(inst1_n498) );
  OAI21_X1 inst1_U387 ( .B1(inst1_n873), .B2(inst1_n1198), .A(inst1_n497),
        .ZN(inst1_stateArray_S02reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst1_U386 ( .A1(ciphertext1[109]), .A2(inst1_n819), .B1(
        plaintext1[109]), .B2(inst1_n507), .ZN(inst1_n497) );
  OAI21_X1 inst1_U385 ( .B1(inst1_n874), .B2(inst1_n1198), .A(inst1_n496),
        .ZN(inst1_stateArray_S02reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst1_U384 ( .A1(ciphertext1[110]), .A2(inst1_n720), .B1(
        plaintext1[110]), .B2(inst1_n507), .ZN(inst1_n496) );
  INV_X1 inst1_U383 ( .A(inst1_n6), .ZN(inst1_n507) );
  OAI21_X1 inst1_U382 ( .B1(inst1_n875), .B2(inst1_n1198), .A(inst1_n495),
        .ZN(inst1_stateArray_S02reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst1_U381 ( .A1(ciphertext1[111]), .A2(inst1_n819), .B1(
        plaintext1[111]), .B2(inst1_n494), .ZN(inst1_n495) );
  OAI211_X1 inst1_U380 ( .C1(inst1_n1220), .C2(inst1_n493), .A(inst1_n492),
        .B(inst1_n491), .ZN(inst1_stateArray_S23reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst1_U379 ( .B1(inst1_n1217), .B2(ciphertext1[48]), .A(inst1_n490),
        .ZN(inst1_n491) );
  OAI22_X1 inst1_U378 ( .A1(inst1_n1113), .A2(inst1_n1015), .B1(inst1_n666),
        .B2(inst1_n1233), .ZN(inst1_n490) );
  AOI22_X1 inst1_U377 ( .A1(inst1_n677), .A2(ciphertext1[32]), .B1(
        plaintext1[32]), .B2(inst1_n596), .ZN(inst1_n492) );
  INV_X1 inst1_U376 ( .A(inst1_n6), .ZN(inst1_n596) );
  XNOR2_X1 inst1_U375 ( .A(inst1_n616), .B(inst1_n489), .ZN(inst1_n493) );
  AOI22_X1 inst1_U374 ( .A1(inst1_n1113), .A2(inst1_n1212), .B1(inst1_n1211),
        .B2(ciphertext1[24]), .ZN(inst1_n489) );
  INV_X1 inst1_U373 ( .A(inst1_n1212), .ZN(inst1_n1211) );
  OAI211_X1 inst1_U372 ( .C1(inst1_n488), .C2(inst1_n1220), .A(inst1_n487),
        .B(inst1_n486), .ZN(inst1_stateArray_S23reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst1_U371 ( .B1(inst1_n1217), .B2(ciphertext1[53]), .A(inst1_n485),
        .ZN(inst1_n486) );
  OAI22_X1 inst1_U370 ( .A1(inst1_n1035), .A2(inst1_n1229), .B1(inst1_n666),
        .B2(inst1_n1249), .ZN(inst1_n485) );
  AOI22_X1 inst1_U369 ( .A1(inst1_n677), .A2(ciphertext1[37]), .B1(
        plaintext1[37]), .B2(inst1_n494), .ZN(inst1_n487) );
  XNOR2_X1 inst1_U368 ( .A(inst1_n484), .B(inst1_n483), .ZN(inst1_n488) );
  AOI22_X1 inst1_U367 ( .A1(inst1_n533), .A2(ciphertext1[28]), .B1(inst1_n1105), .B2(inst1_n532), .ZN(inst1_n483) );
  INV_X1 inst1_U366 ( .A(inst1_n533), .ZN(inst1_n532) );
  AOI22_X1 inst1_U365 ( .A1(ciphertext1[60]), .A2(inst1_n1122), .B1(
        ciphertext1[93]), .B2(inst1_n1234), .ZN(inst1_n484) );
  OAI211_X1 inst1_U364 ( .C1(inst1_n482), .C2(inst1_n1207), .A(inst1_n481),
        .B(inst1_n480), .ZN(inst1_stateArray_S23reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst1_U363 ( .B1(inst1_n1217), .B2(ciphertext1[54]), .A(inst1_n479),
        .ZN(inst1_n480) );
  OAI22_X1 inst1_U362 ( .A1(inst1_n1097), .A2(inst1_n1035), .B1(inst1_n666),
        .B2(inst1_n1232), .ZN(inst1_n479) );
  AOI22_X1 inst1_U361 ( .A1(done1), .A2(ciphertext1[38]), .B1(plaintext1[38]),
        .B2(inst1_n494), .ZN(inst1_n481) );
  XNOR2_X1 inst1_U360 ( .A(inst1_n478), .B(inst1_n477), .ZN(inst1_n482) );
  AOI22_X1 inst1_U359 ( .A1(inst1_n1106), .A2(inst1_n1229), .B1(
        ciphertext1[29]), .B2(ciphertext1[94]), .ZN(inst1_n477) );
  AOI22_X1 inst1_U358 ( .A1(inst1_n526), .A2(ciphertext1[61]), .B1(inst1_n1249), .B2(inst1_n527), .ZN(inst1_n478) );
  INV_X1 inst1_U357 ( .A(inst1_n526), .ZN(inst1_n527) );
  OAI211_X1 inst1_U356 ( .C1(inst1_n476), .C2(inst1_n1220), .A(inst1_n475),
        .B(inst1_n474), .ZN(inst1_stateArray_S23reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst1_U355 ( .B1(inst1_n1217), .B2(ciphertext1[55]), .A(inst1_n473),
        .ZN(inst1_n474) );
  OAI22_X1 inst1_U354 ( .A1(inst1_n1093), .A2(inst1_n1215), .B1(inst1_n1035),
        .B2(inst1_n1230), .ZN(inst1_n473) );
  AOI22_X1 inst1_U353 ( .A1(done1), .A2(ciphertext1[39]), .B1(plaintext1[39]),
        .B2(inst1_n494), .ZN(inst1_n475) );
  XNOR2_X1 inst1_U352 ( .A(inst1_n472), .B(inst1_n471), .ZN(inst1_n476) );
  AOI22_X1 inst1_U351 ( .A1(inst1_n1097), .A2(inst1_n1232), .B1(
        ciphertext1[62]), .B2(ciphertext1[30]), .ZN(inst1_n471) );
  AOI22_X1 inst1_U350 ( .A1(ciphertext1[31]), .A2(inst1_n660), .B1(inst1_n659),
        .B2(inst1_n1230), .ZN(inst1_n472) );
  INV_X1 inst1_U349 ( .A(inst1_n660), .ZN(inst1_n659) );
  OAI211_X1 inst1_U348 ( .C1(inst1_n470), .C2(inst1_n1207), .A(inst1_n469),
        .B(inst1_n468), .ZN(inst1_stateArray_S23reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst1_U347 ( .B1(inst1_n1217), .B2(ciphertext1[51]), .A(inst1_n467),
        .ZN(inst1_n468) );
  OAI22_X1 inst1_U346 ( .A1(inst1_n1116), .A2(inst1_n1215), .B1(inst1_n1035),
        .B2(inst1_n1231), .ZN(inst1_n467) );
  AOI22_X1 inst1_U345 ( .A1(inst1_n677), .A2(ciphertext1[35]), .B1(
        plaintext1[35]), .B2(inst1_n494), .ZN(inst1_n469) );
  XNOR2_X1 inst1_U344 ( .A(inst1_n466), .B(inst1_n465), .ZN(inst1_n470) );
  AOI22_X1 inst1_U343 ( .A1(ciphertext1[27]), .A2(inst1_n581), .B1(inst1_n580),
        .B2(inst1_n1231), .ZN(inst1_n465) );
  INV_X1 inst1_U342 ( .A(inst1_n581), .ZN(inst1_n580) );
  XNOR2_X1 inst1_U341 ( .A(inst1_n1212), .B(inst1_n464), .ZN(inst1_n466) );
  AOI22_X1 inst1_U340 ( .A1(inst1_n1109), .A2(inst1_n1119), .B1(
        ciphertext1[58]), .B2(ciphertext1[26]), .ZN(inst1_n464) );
  AOI22_X1 inst1_U339 ( .A1(ciphertext1[31]), .A2(inst1_n1093), .B1(
        ciphertext1[63]), .B2(inst1_n1230), .ZN(inst1_n1212) );
  NAND2_X1 inst1_U338 ( .A1(inst1_n463), .A2(inst1_n462), .ZN(
        inst1_stateArray_S33reg_gff_1_SFF_0_n5) );
  AOI22_X1 inst1_U337 ( .A1(inst1_n461), .A2(inst1_n460), .B1(inst1_n459),
        .B2(inst1_n458), .ZN(inst1_n462) );
  AOI211_X1 inst1_U336 ( .C1(plaintext1[0]), .C2(inst1_n1228), .A(inst1_n457),
        .B(inst1_n456), .ZN(inst1_n463) );
  OAI22_X1 inst1_U335 ( .A1(inst1_n455), .A2(inst1_n1207), .B1(inst1_n940),
        .B2(inst1_n1142), .ZN(inst1_n456) );
  XNOR2_X1 inst1_U334 ( .A(inst1_n616), .B(inst1_n454), .ZN(inst1_n455) );
  AOI22_X1 inst1_U333 ( .A1(inst1_n453), .A2(inst1_n1233), .B1(ciphertext1[56]), .B2(inst1_n452), .ZN(inst1_n454) );
  AOI22_X1 inst1_U332 ( .A1(inst1_n1102), .A2(inst1_n1103), .B1(
        ciphertext1[88]), .B2(ciphertext1[120]), .ZN(inst1_n616) );
  OAI22_X1 inst1_U331 ( .A1(inst1_n1113), .A2(inst1_n1215), .B1(inst1_n932),
        .B2(inst1_n1182), .ZN(inst1_n457) );
  NAND2_X1 inst1_U330 ( .A1(inst1_n451), .A2(inst1_n450), .ZN(
        inst1_stateArray_S33reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst1_U329 ( .A1(inst1_n449), .A2(inst1_n460), .B1(inst1_n459),
        .B2(inst1_n448), .ZN(inst1_n450) );
  AOI211_X1 inst1_U328 ( .C1(plaintext1[1]), .C2(inst1_n1228), .A(inst1_n447),
        .B(inst1_n446), .ZN(inst1_n451) );
  OAI22_X1 inst1_U327 ( .A1(inst1_n445), .A2(inst1_n1207), .B1(inst1_n941),
        .B2(inst1_n1142), .ZN(inst1_n446) );
  XNOR2_X1 inst1_U326 ( .A(inst1_n444), .B(inst1_n443), .ZN(inst1_n445) );
  AOI22_X1 inst1_U325 ( .A1(inst1_n1102), .A2(inst1_n453), .B1(inst1_n452),
        .B2(ciphertext1[120]), .ZN(inst1_n443) );
  XNOR2_X1 inst1_U324 ( .A(inst1_n1210), .B(inst1_n442), .ZN(inst1_n444) );
  AOI22_X1 inst1_U323 ( .A1(inst1_n1113), .A2(ciphertext1[57]), .B1(
        inst1_n1235), .B2(ciphertext1[24]), .ZN(inst1_n442) );
  AOI22_X1 inst1_U322 ( .A1(inst1_n1114), .A2(inst1_n1115), .B1(
        ciphertext1[89]), .B2(ciphertext1[121]), .ZN(inst1_n1210) );
  OAI22_X1 inst1_U321 ( .A1(inst1_n1121), .A2(inst1_n1215), .B1(inst1_n933),
        .B2(inst1_n1182), .ZN(inst1_n447) );
  NAND2_X1 inst1_U320 ( .A1(inst1_n441), .A2(inst1_n440), .ZN(
        inst1_stateArray_S33reg_gff_1_SFF_2_n5) );
  AOI22_X1 inst1_U319 ( .A1(inst1_n439), .A2(inst1_n459), .B1(inst1_n460),
        .B2(inst1_n438), .ZN(inst1_n440) );
  AOI211_X1 inst1_U318 ( .C1(plaintext1[2]), .C2(inst1_n1228), .A(inst1_n437),
        .B(inst1_n436), .ZN(inst1_n441) );
  OAI22_X1 inst1_U317 ( .A1(inst1_n942), .A2(inst1_n1142), .B1(inst1_n1207),
        .B2(inst1_n435), .ZN(inst1_n436) );
  XNOR2_X1 inst1_U316 ( .A(inst1_n434), .B(inst1_n433), .ZN(inst1_n435) );
  AOI22_X1 inst1_U315 ( .A1(ciphertext1[122]), .A2(ciphertext1[121]), .B1(
        inst1_n1114), .B2(inst1_n1227), .ZN(inst1_n433) );
  XNOR2_X1 inst1_U314 ( .A(inst1_n1121), .B(inst1_n599), .ZN(inst1_n434) );
  AOI22_X1 inst1_U313 ( .A1(inst1_n1118), .A2(inst1_n1119), .B1(
        ciphertext1[58]), .B2(ciphertext1[90]), .ZN(inst1_n599) );
  OAI22_X1 inst1_U312 ( .A1(inst1_n1109), .A2(inst1_n1215), .B1(inst1_n934),
        .B2(inst1_n1182), .ZN(inst1_n437) );
  NAND2_X1 inst1_U311 ( .A1(inst1_n432), .A2(inst1_n431), .ZN(
        inst1_stateArray_S33reg_gff_1_SFF_3_n5) );
  AOI22_X1 inst1_U310 ( .A1(inst1_n430), .A2(inst1_n460), .B1(inst1_n429),
        .B2(inst1_n459), .ZN(inst1_n431) );
  AOI211_X1 inst1_U309 ( .C1(plaintext1[3]), .C2(inst1_n1228), .A(inst1_n428),
        .B(inst1_n427), .ZN(inst1_n432) );
  OAI22_X1 inst1_U308 ( .A1(inst1_n426), .A2(inst1_n1207), .B1(inst1_n943),
        .B2(inst1_n1142), .ZN(inst1_n427) );
  XNOR2_X1 inst1_U307 ( .A(inst1_n425), .B(inst1_n424), .ZN(inst1_n426) );
  AOI22_X1 inst1_U306 ( .A1(inst1_n453), .A2(inst1_n1116), .B1(ciphertext1[59]), .B2(inst1_n452), .ZN(inst1_n424) );
  INV_X1 inst1_U305 ( .A(inst1_n453), .ZN(inst1_n452) );
  XNOR2_X1 inst1_U304 ( .A(inst1_n1200), .B(inst1_n581), .ZN(inst1_n425) );
  AOI22_X1 inst1_U303 ( .A1(inst1_n1110), .A2(inst1_n1111), .B1(
        ciphertext1[91]), .B2(ciphertext1[123]), .ZN(inst1_n581) );
  AOI22_X1 inst1_U302 ( .A1(ciphertext1[122]), .A2(inst1_n1109), .B1(
        ciphertext1[26]), .B2(inst1_n1227), .ZN(inst1_n1200) );
  OAI22_X1 inst1_U301 ( .A1(inst1_n935), .A2(inst1_n1185), .B1(inst1_n1215),
        .B2(inst1_n1231), .ZN(inst1_n428) );
  NAND2_X1 inst1_U300 ( .A1(inst1_n423), .A2(inst1_n422), .ZN(
        inst1_stateArray_S33reg_gff_1_SFF_4_n5) );
  AOI22_X1 inst1_U299 ( .A1(inst1_n459), .A2(inst1_n421), .B1(inst1_n460),
        .B2(inst1_n420), .ZN(inst1_n422) );
  AOI211_X1 inst1_U298 ( .C1(plaintext1[4]), .C2(inst1_n1228), .A(inst1_n419),
        .B(inst1_n418), .ZN(inst1_n423) );
  OAI22_X1 inst1_U297 ( .A1(inst1_n417), .A2(inst1_n1207), .B1(inst1_n944),
        .B2(inst1_n1145), .ZN(inst1_n418) );
  XNOR2_X1 inst1_U296 ( .A(inst1_n416), .B(inst1_n415), .ZN(inst1_n417) );
  XNOR2_X1 inst1_U295 ( .A(inst1_n1110), .B(inst1_n582), .ZN(inst1_n415) );
  AOI22_X1 inst1_U294 ( .A1(inst1_n1100), .A2(ciphertext1[60]), .B1(
        inst1_n1234), .B2(ciphertext1[92]), .ZN(inst1_n582) );
  XOR2_X1 inst1_U293 ( .A(inst1_n414), .B(inst1_n453), .Z(inst1_n416) );
  AOI22_X1 inst1_U292 ( .A1(inst1_n1094), .A2(ciphertext1[31]), .B1(
        inst1_n1230), .B2(ciphertext1[127]), .ZN(inst1_n453) );
  AOI22_X1 inst1_U291 ( .A1(ciphertext1[124]), .A2(ciphertext1[27]), .B1(
        inst1_n1231), .B2(inst1_n1225), .ZN(inst1_n414) );
  OAI22_X1 inst1_U290 ( .A1(inst1_n1105), .A2(inst1_n1215), .B1(inst1_n936),
        .B2(inst1_n1182), .ZN(inst1_n419) );
  NAND2_X1 inst1_U289 ( .A1(inst1_n413), .A2(inst1_n412), .ZN(
        inst1_stateArray_S33reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst1_U288 ( .A1(inst1_n411), .A2(inst1_n460), .B1(inst1_n459),
        .B2(inst1_n410), .ZN(inst1_n412) );
  AOI211_X1 inst1_U287 ( .C1(plaintext1[5]), .C2(inst1_n1228), .A(inst1_n409),
        .B(inst1_n408), .ZN(inst1_n413) );
  OAI22_X1 inst1_U286 ( .A1(inst1_n407), .A2(inst1_n1207), .B1(inst1_n945),
        .B2(inst1_n1145), .ZN(inst1_n408) );
  XNOR2_X1 inst1_U285 ( .A(inst1_n406), .B(inst1_n590), .ZN(inst1_n407) );
  AOI22_X1 inst1_U284 ( .A1(ciphertext1[61]), .A2(inst1_n1122), .B1(
        ciphertext1[93]), .B2(inst1_n1249), .ZN(inst1_n590) );
  XNOR2_X1 inst1_U283 ( .A(inst1_n1098), .B(inst1_n1191), .ZN(inst1_n406) );
  AOI22_X1 inst1_U282 ( .A1(ciphertext1[124]), .A2(inst1_n1105), .B1(
        ciphertext1[28]), .B2(inst1_n1225), .ZN(inst1_n1191) );
  OAI22_X1 inst1_U281 ( .A1(inst1_n937), .A2(inst1_n1185), .B1(inst1_n666),
        .B2(inst1_n1229), .ZN(inst1_n409) );
  NAND2_X1 inst1_U280 ( .A1(inst1_n405), .A2(inst1_n404), .ZN(
        inst1_stateArray_S33reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst1_U279 ( .A1(inst1_n403), .A2(inst1_n460), .B1(inst1_n459),
        .B2(inst1_n402), .ZN(inst1_n404) );
  AOI211_X1 inst1_U278 ( .C1(plaintext1[6]), .C2(inst1_n1228), .A(inst1_n401),
        .B(inst1_n400), .ZN(inst1_n405) );
  OAI22_X1 inst1_U277 ( .A1(inst1_n399), .A2(inst1_n1207), .B1(inst1_n946),
        .B2(inst1_n1145), .ZN(inst1_n400) );
  XNOR2_X1 inst1_U276 ( .A(inst1_n398), .B(inst1_n533), .ZN(inst1_n399) );
  AOI22_X1 inst1_U275 ( .A1(inst1_n1098), .A2(ciphertext1[29]), .B1(
        inst1_n1229), .B2(ciphertext1[125]), .ZN(inst1_n533) );
  XNOR2_X1 inst1_U274 ( .A(inst1_n1096), .B(inst1_n604), .ZN(inst1_n398) );
  AOI22_X1 inst1_U273 ( .A1(ciphertext1[62]), .A2(inst1_n1106), .B1(
        ciphertext1[94]), .B2(inst1_n1232), .ZN(inst1_n604) );
  OAI22_X1 inst1_U272 ( .A1(inst1_n1097), .A2(inst1_n1215), .B1(inst1_n938),
        .B2(inst1_n1182), .ZN(inst1_n401) );
  INV_X1 inst1_U271 ( .A(inst1_n1217), .ZN(inst1_n1182) );
  NAND2_X1 inst1_U270 ( .A1(inst1_n397), .A2(inst1_n396), .ZN(
        inst1_stateArray_S33reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst1_U269 ( .A1(inst1_n395), .A2(inst1_n460), .B1(inst1_n459),
        .B2(inst1_n394), .ZN(inst1_n396) );
  NOR2_X1 inst1_U268 ( .A1(inst1_n393), .A2(inst1_n1015), .ZN(inst1_n459) );
  NOR2_X1 inst1_U267 ( .A1(inst1_n1035), .A2(inst1_n392), .ZN(inst1_n460) );
  AOI211_X1 inst1_U266 ( .C1(plaintext1[7]), .C2(inst1_n1228), .A(inst1_n391),
        .B(inst1_n390), .ZN(inst1_n397) );
  OAI22_X1 inst1_U265 ( .A1(inst1_n389), .A2(inst1_n1207), .B1(inst1_n947),
        .B2(inst1_n1145), .ZN(inst1_n390) );
  INV_X1 inst1_U264 ( .A(inst1_n663), .ZN(inst1_n1207) );
  INV_X1 inst1_U263 ( .A(inst1_n1220), .ZN(inst1_n663) );
  NAND2_X1 inst1_U262 ( .A1(inst1_n1018), .A2(inst1_n392), .ZN(inst1_n1220) );
  INV_X1 inst1_U261 ( .A(inst1_n393), .ZN(inst1_n392) );
  XNOR2_X1 inst1_U260 ( .A(inst1_n388), .B(inst1_n526), .ZN(inst1_n389) );
  AOI22_X1 inst1_U259 ( .A1(inst1_n1096), .A2(inst1_n1097), .B1(
        ciphertext1[30]), .B2(ciphertext1[126]), .ZN(inst1_n526) );
  XNOR2_X1 inst1_U258 ( .A(inst1_n1093), .B(inst1_n660), .ZN(inst1_n388) );
  AOI22_X1 inst1_U257 ( .A1(inst1_n1094), .A2(inst1_n1092), .B1(
        ciphertext1[95]), .B2(ciphertext1[127]), .ZN(inst1_n660) );
  OAI22_X1 inst1_U256 ( .A1(inst1_n939), .A2(inst1_n1185), .B1(inst1_n1215),
        .B2(inst1_n1230), .ZN(inst1_n391) );
  INV_X1 inst1_U255 ( .A(inst1_n387), .ZN(inst1_n1215) );
  INV_X1 inst1_U254 ( .A(inst1_n666), .ZN(inst1_n387) );
  NAND2_X1 inst1_U253 ( .A1(inst1_n1032), .A2(inst1_n393), .ZN(inst1_n666) );
  INV_X2 inst1_U252 ( .A(inst1_n386), .ZN(inst1_n1032) );
  INV_X1 inst1_U251 ( .A(inst1_n1217), .ZN(inst1_n1185) );
  AND2_X2 inst1_U250 ( .A1(inst1_n859), .A2(inst1_n1142), .ZN(inst1_n1217) );
  INV_X1 inst1_U249 ( .A(inst1_n385), .ZN(inst1_n1142) );
  INV_X1 inst1_U248 ( .A(inst1_n1135), .ZN(inst1_n385) );
  OAI211_X1 inst1_U247 ( .C1(inst1_n1262), .C2(inst1_n1035), .A(inst1_n384),
        .B(inst1_n383), .ZN(inst1_KeyArray_S30reg_gff_1_SFF_3_n6) );
  OAI21_X1 inst1_U246 ( .B1(inst1_n1088), .B2(inst1_n382), .A(inst1_n381),
        .ZN(inst1_n383) );
  AOI21_X1 inst1_U245 ( .B1(inst1_n1088), .B2(inst1_n382), .A(inst1_n686),
        .ZN(inst1_n381) );
  XNOR2_X1 inst1_U244 ( .A(inst1_n429), .B(inst1_n380), .ZN(inst1_n382) );
  NOR2_X1 inst1_U243 ( .A1(inst1_n1076), .A2(inst1_n1072), .ZN(inst1_n380) );
  XNOR2_X1 inst1_U242 ( .A(inst1_n379), .B(inst1_n378), .ZN(inst1_n429) );
  XNOR2_X1 inst1_U241 ( .A(inst1_n377), .B(inst1_n376), .ZN(inst1_n379) );
  AOI22_X1 inst1_U240 ( .A1(inst1_n79), .A2(inst1_n819), .B1(key1[27]), .B2(
        inst1_n494), .ZN(inst1_n384) );
  OAI211_X1 inst1_U239 ( .C1(inst1_n1260), .C2(inst1_n1035), .A(inst1_n375),
        .B(inst1_n374), .ZN(inst1_KeyArray_S30reg_gff_1_SFF_6_n6) );
  OAI21_X1 inst1_U238 ( .B1(inst1_n1090), .B2(inst1_n373), .A(inst1_n372),
        .ZN(inst1_n374) );
  AOI21_X1 inst1_U237 ( .B1(inst1_n1090), .B2(inst1_n373), .A(inst1_n686),
        .ZN(inst1_n372) );
  XNOR2_X1 inst1_U236 ( .A(inst1_n371), .B(inst1_n402), .ZN(inst1_n373) );
  XNOR2_X1 inst1_U235 ( .A(inst1_n370), .B(inst1_n369), .ZN(inst1_n402) );
  XNOR2_X1 inst1_U234 ( .A(inst1_n368), .B(inst1_n367), .ZN(inst1_n370) );
  NOR2_X1 inst1_U233 ( .A1(inst1_n1071), .A2(inst1_n1076), .ZN(inst1_n371) );
  AOI22_X1 inst1_U232 ( .A1(inst1_n76), .A2(inst1_n720), .B1(key1[30]), .B2(
        inst1_n494), .ZN(inst1_n375) );
  OAI211_X1 inst1_U231 ( .C1(inst1_n1288), .C2(inst1_n1035), .A(inst1_n366),
        .B(inst1_n365), .ZN(inst1_KeyArray_S30reg_gff_1_SFF_1_n6) );
  OAI21_X1 inst1_U230 ( .B1(inst1_n1086), .B2(inst1_n364), .A(inst1_n363),
        .ZN(inst1_n365) );
  AOI21_X1 inst1_U229 ( .B1(inst1_n1086), .B2(inst1_n364), .A(inst1_n686),
        .ZN(inst1_n363) );
  XNOR2_X1 inst1_U228 ( .A(inst1_n362), .B(inst1_n448), .ZN(inst1_n364) );
  XNOR2_X1 inst1_U227 ( .A(inst1_n368), .B(inst1_n361), .ZN(inst1_n448) );
  XNOR2_X1 inst1_U226 ( .A(inst1_n360), .B(inst1_n359), .ZN(inst1_n361) );
  XOR2_X1 inst1_U225 ( .A(inst1_n378), .B(inst1_n358), .Z(inst1_n359) );
  XOR2_X1 inst1_U224 ( .A(inst1_n357), .B(inst1_n356), .Z(inst1_n378) );
  NOR2_X1 inst1_U223 ( .A1(inst1_n1074), .A2(inst1_n1076), .ZN(inst1_n362) );
  AOI22_X1 inst1_U222 ( .A1(inst1_n81), .A2(inst1_n819), .B1(key1[25]), .B2(
        inst1_n494), .ZN(inst1_n366) );
  OAI211_X1 inst1_U221 ( .C1(inst1_n1238), .C2(inst1_n1035), .A(inst1_n355),
        .B(inst1_n354), .ZN(inst1_KeyArray_S30reg_gff_1_SFF_2_n6) );
  OAI21_X1 inst1_U220 ( .B1(inst1_n1087), .B2(inst1_n353), .A(inst1_n352),
        .ZN(inst1_n354) );
  AOI21_X1 inst1_U219 ( .B1(inst1_n1087), .B2(inst1_n353), .A(inst1_n686),
        .ZN(inst1_n352) );
  XNOR2_X1 inst1_U218 ( .A(inst1_n351), .B(inst1_n439), .ZN(inst1_n353) );
  XNOR2_X1 inst1_U217 ( .A(inst1_n350), .B(inst1_n349), .ZN(inst1_n439) );
  XNOR2_X1 inst1_U216 ( .A(inst1_n348), .B(inst1_n347), .ZN(inst1_n350) );
  XNOR2_X1 inst1_U215 ( .A(inst1_n346), .B(inst1_n345), .ZN(inst1_n348) );
  NOR2_X1 inst1_U214 ( .A1(inst1_n344), .A2(inst1_n343), .ZN(inst1_n345) );
  AOI21_X1 inst1_U213 ( .B1(inst1_n342), .B2(inst1_n341), .A(inst1_n340), .ZN(
        inst1_n343) );
  NOR2_X1 inst1_U212 ( .A1(inst1_n1073), .A2(inst1_n1076), .ZN(inst1_n351) );
  AOI22_X1 inst1_U211 ( .A1(inst1_n80), .A2(inst1_n720), .B1(key1[26]), .B2(
        inst1_n494), .ZN(inst1_n355) );
  OAI211_X1 inst1_U210 ( .C1(inst1_n1237), .C2(inst1_n1035), .A(inst1_n339),
        .B(inst1_n338), .ZN(inst1_KeyArray_S30reg_gff_1_SFF_4_n6) );
  OAI21_X1 inst1_U209 ( .B1(inst1_n1089), .B2(inst1_n337), .A(inst1_n336),
        .ZN(inst1_n338) );
  AOI21_X1 inst1_U208 ( .B1(inst1_n1089), .B2(inst1_n337), .A(inst1_n686),
        .ZN(inst1_n336) );
  XNOR2_X1 inst1_U207 ( .A(inst1_n335), .B(inst1_n421), .ZN(inst1_n337) );
  XNOR2_X1 inst1_U206 ( .A(inst1_n334), .B(inst1_n369), .ZN(inst1_n421) );
  XNOR2_X1 inst1_U205 ( .A(inst1_n333), .B(inst1_n377), .ZN(inst1_n369) );
  XNOR2_X1 inst1_U204 ( .A(inst1_n332), .B(inst1_n331), .ZN(inst1_n377) );
  NAND2_X1 inst1_U203 ( .A1(inst1_n330), .A2(inst1_n329), .ZN(inst1_n332) );
  NOR2_X1 inst1_U202 ( .A1(inst1_n1076), .A2(inst1_n1060), .ZN(inst1_n335) );
  AOI22_X1 inst1_U201 ( .A1(inst1_n78), .A2(inst1_n819), .B1(key1[28]), .B2(
        inst1_n494), .ZN(inst1_n339) );
  INV_X1 inst1_U200 ( .A(inst1_n1006), .ZN(inst1_n819) );
  INV_X1 inst1_U199 ( .A(inst1_n720), .ZN(inst1_n1006) );
  OAI211_X1 inst1_U198 ( .C1(inst1_n1259), .C2(inst1_n1035), .A(inst1_n328),
        .B(inst1_n327), .ZN(inst1_KeyArray_S30reg_gff_1_SFF_7_n6) );
  OAI21_X1 inst1_U197 ( .B1(inst1_n1091), .B2(inst1_n326), .A(inst1_n325),
        .ZN(inst1_n327) );
  AOI21_X1 inst1_U196 ( .B1(inst1_n1091), .B2(inst1_n326), .A(inst1_n686),
        .ZN(inst1_n325) );
  XNOR2_X1 inst1_U195 ( .A(inst1_n324), .B(inst1_n394), .ZN(inst1_n326) );
  XNOR2_X1 inst1_U194 ( .A(inst1_n323), .B(inst1_n346), .ZN(inst1_n394) );
  XOR2_X1 inst1_U193 ( .A(inst1_n334), .B(inst1_n368), .Z(inst1_n346) );
  AOI221_X1 inst1_U192 ( .B1(inst1_n322), .B2(inst1_n321), .C1(inst1_n320),
        .C2(inst1_n319), .A(inst1_n318), .ZN(inst1_n368) );
  INV_X1 inst1_U191 ( .A(inst1_n319), .ZN(inst1_n321) );
  XNOR2_X1 inst1_U190 ( .A(inst1_n357), .B(inst1_n317), .ZN(inst1_n334) );
  AND2_X1 inst1_U189 ( .A1(inst1_n316), .A2(inst1_n315), .ZN(inst1_n357) );
  XNOR2_X1 inst1_U188 ( .A(inst1_n331), .B(inst1_n367), .ZN(inst1_n323) );
  XNOR2_X1 inst1_U187 ( .A(inst1_n314), .B(inst1_n349), .ZN(inst1_n331) );
  XNOR2_X1 inst1_U186 ( .A(inst1_n313), .B(inst1_n312), .ZN(inst1_n349) );
  NAND2_X1 inst1_U185 ( .A1(inst1_n330), .A2(inst1_n311), .ZN(inst1_n313) );
  XNOR2_X1 inst1_U184 ( .A(inst1_n310), .B(inst1_n309), .ZN(inst1_n330) );
  XNOR2_X1 inst1_U183 ( .A(inst1_n308), .B(inst1_n307), .ZN(inst1_n310) );
  NOR2_X1 inst1_U182 ( .A1(inst1_n306), .A2(inst1_n305), .ZN(inst1_n314) );
  NOR2_X1 inst1_U181 ( .A1(inst1_n1070), .A2(inst1_n1076), .ZN(inst1_n324) );
  AOI22_X1 inst1_U180 ( .A1(inst1_n75), .A2(inst1_n720), .B1(key1[31]), .B2(
        inst1_n494), .ZN(inst1_n328) );
  OAI211_X1 inst1_U179 ( .C1(inst1_n1239), .C2(inst1_n1203), .A(inst1_n304),
        .B(inst1_n303), .ZN(inst1_KeyArray_S30reg_gff_1_SFF_0_n6) );
  OAI21_X1 inst1_U178 ( .B1(inst1_n1085), .B2(inst1_n302), .A(inst1_n301),
        .ZN(inst1_n303) );
  AOI21_X1 inst1_U177 ( .B1(inst1_n1085), .B2(inst1_n302), .A(inst1_n686),
        .ZN(inst1_n301) );
  XNOR2_X1 inst1_U176 ( .A(inst1_n300), .B(inst1_n458), .ZN(inst1_n302) );
  XNOR2_X1 inst1_U175 ( .A(inst1_n299), .B(inst1_n360), .ZN(inst1_n458) );
  XNOR2_X1 inst1_U174 ( .A(inst1_n312), .B(inst1_n298), .ZN(inst1_n360) );
  OAI211_X1 inst1_U173 ( .C1(inst1_n297), .C2(inst1_n296), .A(inst1_n315), .B(
        inst1_n295), .ZN(inst1_n298) );
  XNOR2_X1 inst1_U172 ( .A(inst1_n294), .B(inst1_n307), .ZN(inst1_n315) );
  XOR2_X1 inst1_U171 ( .A(inst1_n293), .B(inst1_n292), .Z(inst1_n307) );
  XNOR2_X1 inst1_U170 ( .A(inst1_n291), .B(inst1_n290), .ZN(inst1_n294) );
  XNOR2_X1 inst1_U169 ( .A(inst1_n289), .B(inst1_n288), .ZN(inst1_n312) );
  NOR2_X1 inst1_U168 ( .A1(inst1_n319), .A2(inst1_n318), .ZN(inst1_n288) );
  XNOR2_X1 inst1_U167 ( .A(inst1_n287), .B(inst1_n286), .ZN(inst1_n318) );
  XNOR2_X1 inst1_U166 ( .A(inst1_n285), .B(inst1_n284), .ZN(inst1_n287) );
  XNOR2_X1 inst1_U165 ( .A(inst1_n356), .B(inst1_n283), .ZN(inst1_n299) );
  XNOR2_X1 inst1_U164 ( .A(inst1_n282), .B(inst1_n281), .ZN(inst1_n283) );
  XNOR2_X1 inst1_U163 ( .A(inst1_n280), .B(inst1_n317), .ZN(inst1_n282) );
  NAND2_X1 inst1_U162 ( .A1(inst1_n279), .A2(inst1_n278), .ZN(inst1_n317) );
  NOR2_X1 inst1_U161 ( .A1(inst1_n277), .A2(inst1_n276), .ZN(inst1_n356) );
  NOR2_X1 inst1_U160 ( .A1(inst1_n1075), .A2(inst1_n1076), .ZN(inst1_n300) );
  AOI22_X1 inst1_U159 ( .A1(inst1_n82), .A2(inst1_n720), .B1(key1[24]), .B2(
        inst1_n494), .ZN(inst1_n304) );
  INV_X1 inst1_U158 ( .A(inst1_n6), .ZN(inst1_n494) );
  INV_X1 inst1_U157 ( .A(inst1_n894), .ZN(inst1_n1203) );
  OAI211_X1 inst1_U156 ( .C1(inst1_n1261), .C2(inst1_n1035), .A(inst1_n275),
        .B(inst1_n274), .ZN(inst1_KeyArray_S30reg_gff_1_SFF_5_n6) );
  OAI21_X1 inst1_U155 ( .B1(inst1_n1084), .B2(inst1_n273), .A(inst1_n272),
        .ZN(inst1_n274) );
  AOI21_X1 inst1_U154 ( .B1(inst1_n1084), .B2(inst1_n273), .A(inst1_n686),
        .ZN(inst1_n272) );
  INV_X1 inst1_U153 ( .A(inst1_n1018), .ZN(inst1_n686) );
  NAND2_X1 inst1_U152 ( .A1(inst1_n271), .A2(inst1_n1006), .ZN(inst1_n386) );
  XNOR2_X1 inst1_U151 ( .A(inst1_n270), .B(inst1_n410), .ZN(inst1_n273) );
  XNOR2_X1 inst1_U150 ( .A(inst1_n289), .B(inst1_n269), .ZN(inst1_n410) );
  XNOR2_X1 inst1_U149 ( .A(inst1_n268), .B(inst1_n267), .ZN(inst1_n269) );
  NOR2_X1 inst1_U148 ( .A1(inst1_n266), .A2(inst1_n265), .ZN(inst1_n267) );
  XNOR2_X1 inst1_U147 ( .A(inst1_n367), .B(inst1_n347), .ZN(inst1_n268) );
  XNOR2_X1 inst1_U146 ( .A(inst1_n264), .B(inst1_n263), .ZN(inst1_n347) );
  NOR2_X1 inst1_U145 ( .A1(inst1_n276), .A2(inst1_n262), .ZN(inst1_n263) );
  XNOR2_X1 inst1_U144 ( .A(inst1_n261), .B(inst1_n260), .ZN(inst1_n276) );
  XNOR2_X1 inst1_U143 ( .A(inst1_n280), .B(inst1_n358), .ZN(inst1_n264) );
  XNOR2_X1 inst1_U142 ( .A(inst1_n259), .B(inst1_n281), .ZN(inst1_n358) );
  NAND2_X1 inst1_U141 ( .A1(inst1_n258), .A2(inst1_n278), .ZN(inst1_n281) );
  XNOR2_X1 inst1_U140 ( .A(inst1_n257), .B(inst1_n256), .ZN(inst1_n278) );
  XNOR2_X1 inst1_U139 ( .A(inst1_n255), .B(inst1_n254), .ZN(inst1_n256) );
  XOR2_X1 inst1_U138 ( .A(inst1_n261), .B(inst1_n290), .Z(inst1_n257) );
  NOR2_X1 inst1_U137 ( .A1(inst1_n265), .A2(inst1_n253), .ZN(inst1_n259) );
  XNOR2_X1 inst1_U136 ( .A(inst1_n252), .B(inst1_n286), .ZN(inst1_n265) );
  XNOR2_X1 inst1_U135 ( .A(inst1_n290), .B(inst1_n251), .ZN(inst1_n286) );
  INV_X1 inst1_U134 ( .A(inst1_n309), .ZN(inst1_n251) );
  XNOR2_X1 inst1_U133 ( .A(inst1_n295), .B(inst1_n250), .ZN(inst1_n309) );
  NAND2_X1 inst1_U132 ( .A1(inst1_n249), .A2(inst1_n248), .ZN(inst1_n250) );
  MUX2_X1 inst1_U131 ( .A(inst1_n247), .B(inst1_n246), .S(inst1_n245), .Z(
        inst1_n290) );
  AND2_X1 inst1_U130 ( .A1(inst1_n244), .A2(inst1_n243), .ZN(inst1_n245) );
  AOI22_X1 inst1_U129 ( .A1(inst1_n308), .A2(inst1_n291), .B1(inst1_n242),
        .B2(inst1_n241), .ZN(inst1_n252) );
  INV_X1 inst1_U128 ( .A(inst1_n308), .ZN(inst1_n241) );
  INV_X1 inst1_U127 ( .A(inst1_n242), .ZN(inst1_n291) );
  XOR2_X1 inst1_U126 ( .A(inst1_n333), .B(inst1_n376), .Z(inst1_n280) );
  NOR2_X1 inst1_U125 ( .A1(inst1_n342), .A2(inst1_n344), .ZN(inst1_n376) );
  XNOR2_X1 inst1_U124 ( .A(inst1_n240), .B(inst1_n244), .ZN(inst1_n344) );
  NOR2_X1 inst1_U123 ( .A1(inst1_n239), .A2(inst1_n305), .ZN(inst1_n333) );
  OAI22_X1 inst1_U122 ( .A1(inst1_n249), .A2(inst1_n248), .B1(inst1_n238),
        .B2(inst1_n293), .ZN(inst1_n305) );
  INV_X1 inst1_U121 ( .A(inst1_n254), .ZN(inst1_n293) );
  AND2_X1 inst1_U120 ( .A1(inst1_n238), .A2(inst1_n237), .ZN(inst1_n248) );
  NOR2_X1 inst1_U119 ( .A1(inst1_n236), .A2(inst1_n235), .ZN(inst1_n367) );
  NOR2_X1 inst1_U118 ( .A1(inst1_n234), .A2(inst1_n235), .ZN(inst1_n289) );
  XNOR2_X1 inst1_U117 ( .A(inst1_n233), .B(inst1_n232), .ZN(inst1_n235) );
  XOR2_X1 inst1_U116 ( .A(inst1_n284), .B(inst1_n231), .Z(inst1_n232) );
  NOR2_X1 inst1_U115 ( .A1(inst1_n308), .A2(inst1_n340), .ZN(inst1_n231) );
  XNOR2_X1 inst1_U114 ( .A(inst1_n230), .B(inst1_n240), .ZN(inst1_n284) );
  AOI21_X1 inst1_U113 ( .B1(inst1_n254), .B2(inst1_n237), .A(inst1_n229), .ZN(
        inst1_n240) );
  OAI21_X1 inst1_U112 ( .B1(inst1_n254), .B2(inst1_n237), .A(inst1_n238), .ZN(
        inst1_n229) );
  XOR2_X1 inst1_U111 ( .A(inst1_n228), .B(inst1_n295), .Z(inst1_n238) );
  NAND2_X1 inst1_U110 ( .A1(inst1_n297), .A2(inst1_n296), .ZN(inst1_n295) );
  XNOR2_X1 inst1_U109 ( .A(inst1_n308), .B(inst1_n292), .ZN(inst1_n228) );
  XNOR2_X1 inst1_U108 ( .A(inst1_n227), .B(inst1_n260), .ZN(inst1_n237) );
  XNOR2_X1 inst1_U107 ( .A(inst1_n226), .B(inst1_n340), .ZN(inst1_n260) );
  XNOR2_X1 inst1_U106 ( .A(inst1_n285), .B(inst1_n225), .ZN(inst1_n226) );
  XNOR2_X1 inst1_U105 ( .A(inst1_n224), .B(inst1_n261), .ZN(inst1_n230) );
  XNOR2_X1 inst1_U104 ( .A(inst1_n223), .B(inst1_n222), .ZN(inst1_n261) );
  OAI211_X1 inst1_U103 ( .C1(inst1_n244), .C2(inst1_n254), .A(inst1_n243), .B(
        inst1_n221), .ZN(inst1_n222) );
  NAND2_X1 inst1_U102 ( .A1(inst1_n244), .A2(inst1_n254), .ZN(inst1_n221) );
  XOR2_X1 inst1_U101 ( .A(inst1_n220), .B(inst1_n242), .Z(inst1_n243) );
  XOR2_X1 inst1_U100 ( .A(inst1_n340), .B(inst1_n320), .Z(inst1_n242) );
  NOR2_X1 inst1_U99 ( .A1(inst1_n342), .A2(inst1_n341), .ZN(inst1_n340) );
  XNOR2_X1 inst1_U98 ( .A(inst1_n285), .B(inst1_n219), .ZN(inst1_n341) );
  XOR2_X1 inst1_U97 ( .A(inst1_n247), .B(inst1_n292), .Z(inst1_n220) );
  XNOR2_X1 inst1_U96 ( .A(inst1_n218), .B(inst1_n217), .ZN(inst1_n292) );
  AOI21_X1 inst1_U95 ( .B1(inst1_n247), .B2(inst1_n246), .A(inst1_n216), .ZN(
        inst1_n254) );
  OAI21_X1 inst1_U94 ( .B1(inst1_n247), .B2(inst1_n246), .A(inst1_n249), .ZN(
        inst1_n216) );
  XNOR2_X1 inst1_U93 ( .A(inst1_n215), .B(inst1_n214), .ZN(inst1_n249) );
  NAND2_X1 inst1_U92 ( .A1(inst1_n316), .A2(inst1_n297), .ZN(inst1_n214) );
  INV_X1 inst1_U91 ( .A(inst1_n296), .ZN(inst1_n316) );
  XNOR2_X1 inst1_U90 ( .A(inst1_n285), .B(inst1_n213), .ZN(inst1_n296) );
  XNOR2_X1 inst1_U89 ( .A(inst1_n212), .B(inst1_n211), .ZN(inst1_n215) );
  XNOR2_X1 inst1_U88 ( .A(inst1_n210), .B(inst1_n209), .ZN(inst1_n211) );
  XNOR2_X1 inst1_U87 ( .A(inst1_n208), .B(inst1_n207), .ZN(inst1_n209) );
  XOR2_X1 inst1_U86 ( .A(inst1_n206), .B(inst1_n218), .Z(inst1_n210) );
  XNOR2_X1 inst1_U85 ( .A(inst1_n255), .B(inst1_n227), .ZN(inst1_n246) );
  INV_X1 inst1_U84 ( .A(inst1_n223), .ZN(inst1_n227) );
  XNOR2_X1 inst1_U83 ( .A(inst1_n205), .B(inst1_n204), .ZN(inst1_n255) );
  XNOR2_X1 inst1_U82 ( .A(inst1_n233), .B(inst1_n218), .ZN(inst1_n205) );
  NOR2_X1 inst1_U81 ( .A1(inst1_n322), .A2(inst1_n319), .ZN(inst1_n218) );
  XNOR2_X1 inst1_U80 ( .A(inst1_n208), .B(inst1_n203), .ZN(inst1_n319) );
  AND2_X1 inst1_U79 ( .A1(inst1_n329), .A2(inst1_n311), .ZN(inst1_n247) );
  XNOR2_X1 inst1_U78 ( .A(inst1_n262), .B(inst1_n202), .ZN(inst1_n311) );
  XOR2_X1 inst1_U77 ( .A(inst1_n342), .B(inst1_n239), .Z(inst1_n329) );
  XOR2_X1 inst1_U76 ( .A(inst1_n201), .B(inst1_n200), .Z(inst1_n244) );
  INV_X1 inst1_U75 ( .A(inst1_n225), .ZN(inst1_n200) );
  XOR2_X1 inst1_U74 ( .A(inst1_n204), .B(inst1_n217), .Z(inst1_n225) );
  NOR2_X1 inst1_U73 ( .A1(inst1_n253), .A2(inst1_n266), .ZN(inst1_n217) );
  XNOR2_X1 inst1_U72 ( .A(inst1_n208), .B(inst1_n233), .ZN(inst1_n266) );
  XNOR2_X1 inst1_U71 ( .A(inst1_n199), .B(inst1_n198), .ZN(inst1_n253) );
  XNOR2_X1 inst1_U70 ( .A(inst1_n197), .B(inst1_n322), .ZN(inst1_n199) );
  XNOR2_X1 inst1_U69 ( .A(inst1_n196), .B(inst1_n206), .ZN(inst1_n204) );
  NOR2_X1 inst1_U68 ( .A1(inst1_n234), .A2(inst1_n236), .ZN(inst1_n206) );
  XNOR2_X1 inst1_U67 ( .A(inst1_n195), .B(inst1_n194), .ZN(inst1_n236) );
  XNOR2_X1 inst1_U66 ( .A(inst1_n308), .B(inst1_n212), .ZN(inst1_n201) );
  XNOR2_X1 inst1_U65 ( .A(inst1_n322), .B(inst1_n224), .ZN(inst1_n212) );
  INV_X1 inst1_U64 ( .A(inst1_n320), .ZN(inst1_n322) );
  NOR2_X1 inst1_U63 ( .A1(inst1_n277), .A2(inst1_n262), .ZN(inst1_n308) );
  XNOR2_X1 inst1_U62 ( .A(inst1_n320), .B(inst1_n213), .ZN(inst1_n262) );
  XNOR2_X1 inst1_U61 ( .A(inst1_n285), .B(inst1_n233), .ZN(inst1_n320) );
  XNOR2_X1 inst1_U60 ( .A(inst1_n194), .B(inst1_n213), .ZN(inst1_n277) );
  XNOR2_X1 inst1_U59 ( .A(inst1_n195), .B(inst1_n342), .ZN(inst1_n213) );
  AOI22_X1 inst1_U58 ( .A1(inst1_n271), .A2(inst1_n22), .B1(inst1_n461), .B2(
        inst1_n1223), .ZN(inst1_n342) );
  AOI22_X1 inst1_U57 ( .A1(inst1_n1085), .A2(inst1_n1102), .B1(
        ciphertext1[120]), .B2(inst1_n1248), .ZN(inst1_n461) );
  INV_X1 inst1_U56 ( .A(inst1_n196), .ZN(inst1_n194) );
  XOR2_X1 inst1_U55 ( .A(inst1_n193), .B(inst1_n198), .Z(inst1_n223) );
  INV_X1 inst1_U54 ( .A(inst1_n219), .ZN(inst1_n198) );
  XOR2_X1 inst1_U53 ( .A(inst1_n203), .B(inst1_n195), .Z(inst1_n219) );
  AOI22_X1 inst1_U52 ( .A1(inst1_n271), .A2(inst1_n24), .B1(inst1_n403), .B2(
        inst1_n1223), .ZN(inst1_n195) );
  AOI22_X1 inst1_U51 ( .A1(inst1_n1090), .A2(inst1_n1096), .B1(
        ciphertext1[126]), .B2(inst1_n1244), .ZN(inst1_n403) );
  OR2_X1 inst1_U50 ( .A1(inst1_n306), .A2(inst1_n239), .ZN(inst1_n193) );
  XOR2_X1 inst1_U49 ( .A(inst1_n197), .B(inst1_n234), .Z(inst1_n239) );
  XOR2_X1 inst1_U48 ( .A(inst1_n234), .B(inst1_n202), .Z(inst1_n306) );
  XOR2_X1 inst1_U47 ( .A(inst1_n208), .B(inst1_n297), .Z(inst1_n202) );
  AND2_X1 inst1_U46 ( .A1(inst1_n279), .A2(inst1_n258), .ZN(inst1_n224) );
  XOR2_X1 inst1_U45 ( .A(inst1_n297), .B(inst1_n233), .Z(inst1_n258) );
  XNOR2_X1 inst1_U44 ( .A(inst1_n285), .B(inst1_n196), .ZN(inst1_n279) );
  XOR2_X1 inst1_U43 ( .A(inst1_n208), .B(inst1_n192), .Z(inst1_n196) );
  INV_X1 inst1_U42 ( .A(inst1_n197), .ZN(inst1_n192) );
  XOR2_X1 inst1_U41 ( .A(inst1_n207), .B(inst1_n297), .Z(inst1_n197) );
  AOI22_X1 inst1_U40 ( .A1(inst1_n271), .A2(inst1_n17), .B1(inst1_n449), .B2(
        inst1_n1223), .ZN(inst1_n297) );
  AOI22_X1 inst1_U39 ( .A1(inst1_n1114), .A2(inst1_n1086), .B1(inst1_n1241),
        .B2(ciphertext1[121]), .ZN(inst1_n449) );
  AOI22_X1 inst1_U38 ( .A1(inst1_n271), .A2(inst1_n12), .B1(inst1_n430), .B2(
        inst1_n1223), .ZN(inst1_n207) );
  AOI22_X1 inst1_U37 ( .A1(inst1_n1088), .A2(inst1_n1110), .B1(
        ciphertext1[123]), .B2(inst1_n1247), .ZN(inst1_n430) );
  AOI22_X1 inst1_U36 ( .A1(inst1_n271), .A2(inst1_n14), .B1(inst1_n438), .B2(
        inst1_n1223), .ZN(inst1_n208) );
  AOI22_X1 inst1_U35 ( .A1(ciphertext1[122]), .A2(inst1_n1242), .B1(
        inst1_n1087), .B2(inst1_n1227), .ZN(inst1_n438) );
  AOI22_X1 inst1_U34 ( .A1(inst1_n271), .A2(inst1_n10), .B1(inst1_n411), .B2(
        inst1_n1223), .ZN(inst1_n285) );
  AOI22_X1 inst1_U33 ( .A1(inst1_n1084), .A2(inst1_n1098), .B1(
        ciphertext1[125]), .B2(inst1_n1245), .ZN(inst1_n411) );
  XNOR2_X1 inst1_U32 ( .A(inst1_n233), .B(inst1_n203), .ZN(inst1_n234) );
  AOI22_X1 inst1_U31 ( .A1(inst1_n271), .A2(inst1_n11), .B1(inst1_n420), .B2(
        inst1_n1223), .ZN(inst1_n203) );
  AOI22_X1 inst1_U30 ( .A1(inst1_n1089), .A2(inst1_n1225), .B1(
        ciphertext1[124]), .B2(inst1_n1246), .ZN(inst1_n420) );
  AOI22_X1 inst1_U29 ( .A1(inst1_n271), .A2(inst1_n9), .B1(inst1_n395), .B2(
        inst1_n1223), .ZN(inst1_n233) );
  AOI22_X1 inst1_U28 ( .A1(inst1_n1091), .A2(inst1_n1094), .B1(
        ciphertext1[127]), .B2(inst1_n1243), .ZN(inst1_n395) );
  NOR2_X1 inst1_U27 ( .A1(inst1_n1061), .A2(inst1_n1076), .ZN(inst1_n270) );
  AOI22_X1 inst1_U26 ( .A1(inst1_n77), .A2(inst1_n720), .B1(key1[29]), .B2(
        inst1_n1156), .ZN(inst1_n275) );
  NAND2_X2 inst1_U25 ( .A1(inst1_n191), .A2(inst1_n1223), .ZN(inst1_n1035) );
  NAND2_X1 inst1_U24 ( .A1(inst1_n6), .A2(inst1_ctrl_n6), .ZN(inst1_n1223) );
  NAND2_X1 inst1_U23 ( .A1(inst1_n191), .A2(inst1_n1250), .ZN(
        inst1_ctrl_seq4_SFF_0_n5) );
  INV_X1 inst1_U22 ( .A(inst1_n189), .ZN(inst1_n190) );
  OAI221_X1 inst1_U21 ( .B1(inst1_n1080), .B2(inst1_n851), .C1(inst1_n188),
        .C2(inst1_n385), .A(inst1_n6), .ZN(inst1_ctrl_seq6_SFF_0_n5) );
  NAND2_X1 inst1_U20 ( .A1(inst1_n1080), .A2(inst1_n851), .ZN(inst1_n188) );
  NAND2_X1 inst1_U19 ( .A1(inst1_n6), .A2(inst1_n1081), .ZN(
        inst1_ctrl_seq6_SFF_4_n5) );
  NOR4_X1 inst1_U18 ( .A1(inst1_n1060), .A2(inst1_n1074), .A3(inst1_n1073),
        .A4(inst1_n1061), .ZN(inst1_n393) );
  NAND4_X1 inst1_U17 ( .A1(inst1_n1079), .A2(inst1_n1080), .A3(inst1_n851),
        .A4(inst1_n1081), .ZN(inst1_n189) );
  NAND2_X1 inst1_U16 ( .A1(inst1_n6), .A2(inst1_n1082), .ZN(
        inst1_ctrl_seq6_SFF_2_n5) );
  INV_X1 inst1_U15 ( .A(reset1), .ZN(inst1_n1189) );
  INV_X1 inst1_U14 ( .A(inst1_n1018), .ZN(inst1_n740) );
  INV_X1 inst1_U13 ( .A(inst1_n386), .ZN(inst1_n1018) );
  INV_X1 inst1_U12 ( .A(inst1_n1035), .ZN(inst1_n894) );
  INV_X1 inst1_U11 ( .A(inst1_n894), .ZN(inst1_n1015) );
  INV_X1 inst1_U10 ( .A(inst1_n1223), .ZN(inst1_n271) );
  NAND4_X1 inst1_U9 ( .A1(inst1_n720), .A2(inst1_n393), .A3(inst1_n143), .A4(
        inst1_n1077), .ZN(inst1_n1135) );
  INV_X1 inst1_U8 ( .A(inst1_n1032), .ZN(inst1_n849) );
  INV_X1 inst1_U7 ( .A(inst1_n6), .ZN(inst1_n1156) );
  INV_X1 inst1_U6 ( .A(inst1_n6), .ZN(inst1_n1133) );
  NOR2_X1 inst1_U5 ( .A1(inst1_ctrl_seq6_SFF_2_n5), .A2(inst1_n189), .ZN(
        inst1_n720) );
  AOI21_X4 inst1_U4 ( .B1(inst1_n1082), .B2(inst1_n190), .A(inst1_n1133), .ZN(
        inst1_n191) );
  INV_X4 inst1_U3 ( .A(inst1_n191), .ZN(inst1_n1198) );
  DFF_X2 inst1_nReset_reg_FF_FF ( .D(inst1_n1189), .CK(clk), .Q(inst1_n6),
        .QN(inst1_n1228) );
  DFF_X1 inst1_calcRCon_s_current_state_reg_7__FF_FF ( .D(inst1_calcRCon_n44),
        .CK(clk), .Q(inst1_n1226), .QN(inst1_n1070) );
  DFF_X1 inst1_calcRCon_s_current_state_reg_6__FF_FF ( .D(inst1_calcRCon_n45),
        .CK(clk), .QN(inst1_n1071) );
  DFF_X1 inst1_calcRCon_s_current_state_reg_5__FF_FF ( .D(inst1_calcRCon_n46),
        .CK(clk), .QN(inst1_n1061) );
  DFF_X1 inst1_calcRCon_s_current_state_reg_4__FF_FF ( .D(inst1_calcRCon_n47),
        .CK(clk), .QN(inst1_n1060) );
  DFF_X1 inst1_calcRCon_s_current_state_reg_3__FF_FF ( .D(inst1_calcRCon_n48),
        .CK(clk), .Q(inst1_n1240), .QN(inst1_n1072) );
  DFF_X1 inst1_calcRCon_s_current_state_reg_2__FF_FF ( .D(inst1_calcRCon_n49),
        .CK(clk), .Q(inst1_n1263), .QN(inst1_n1073) );
  DFF_X1 inst1_calcRCon_s_current_state_reg_1__FF_FF ( .D(inst1_calcRCon_n50),
        .CK(clk), .QN(inst1_n1074) );
  DFF_X1 inst1_calcRCon_s_current_state_reg_0__FF_FF ( .D(inst1_calcRCon_n51),
        .CK(clk), .Q(inst1_n1264), .QN(inst1_n1075) );
  DFF_X1 inst1_KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S33reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst1_n1059) );
  DFF_X1 inst1_KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S33reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst1_n1058) );
  DFF_X1 inst1_KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S33reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst1_n1057) );
  DFF_X1 inst1_KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S33reg_gff_1_SFF_4_n5), .CK(clk), .QN(inst1_n1056) );
  DFF_X1 inst1_KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S33reg_gff_1_SFF_3_n5), .CK(clk), .QN(inst1_n1055) );
  DFF_X1 inst1_KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S33reg_gff_1_SFF_2_n5), .CK(clk), .QN(inst1_n1054) );
  DFF_X1 inst1_KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S33reg_gff_1_SFF_1_n5), .CK(clk), .Q(inst1_n57) );
  DFF_X1 inst1_KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S33reg_gff_1_SFF_0_n5), .CK(clk), .QN(inst1_n1052) );
  DFF_X1 inst1_KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S32reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst1_n1051) );
  DFF_X1 inst1_KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S32reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst1_n1050) );
  DFF_X1 inst1_KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S32reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst1_n1049) );
  DFF_X1 inst1_KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S32reg_gff_1_SFF_4_n6), .CK(clk), .QN(inst1_n1048) );
  DFF_X1 inst1_KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S32reg_gff_1_SFF_3_n6), .CK(clk), .QN(inst1_n1047) );
  DFF_X1 inst1_KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S32reg_gff_1_SFF_2_n6), .CK(clk), .QN(inst1_n1046) );
  DFF_X1 inst1_KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S32reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst1_n65) );
  DFF_X1 inst1_KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S32reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst1_n1044) );
  DFF_X1 inst1_KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S31reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst1_n67), .QN(
        inst1_n1259) );
  DFF_X1 inst1_KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S31reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst1_n68), .QN(
        inst1_n1260) );
  DFF_X1 inst1_KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S31reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst1_n69), .QN(
        inst1_n1261) );
  DFF_X1 inst1_KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S31reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst1_n70), .QN(
        inst1_n1237) );
  DFF_X1 inst1_KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S31reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst1_n71), .QN(
        inst1_n1262) );
  DFF_X1 inst1_KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S31reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst1_n72), .QN(
        inst1_n1238) );
  DFF_X1 inst1_KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S31reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst1_n73), .QN(
        inst1_n1288) );
  DFF_X1 inst1_KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S31reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst1_n74), .QN(
        inst1_n1239) );
  DFF_X1 inst1_KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S30reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst1_n75) );
  DFF_X1 inst1_KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S30reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst1_n76) );
  DFF_X1 inst1_KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S30reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst1_n77) );
  DFF_X1 inst1_KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S30reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst1_n78) );
  DFF_X1 inst1_KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S30reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst1_n79) );
  DFF_X1 inst1_KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S30reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst1_n80) );
  DFF_X1 inst1_KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S30reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst1_n81) );
  DFF_X1 inst1_KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S30reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst1_n82) );
  DFF_X1 inst1_KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S23reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst1_n83) );
  DFF_X1 inst1_KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S23reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst1_n84) );
  DFF_X1 inst1_KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S23reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst1_n85) );
  DFF_X1 inst1_KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S23reg_gff_1_SFF_4_n5), .CK(clk), .Q(inst1_n86) );
  DFF_X1 inst1_KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S23reg_gff_1_SFF_3_n5), .CK(clk), .Q(inst1_n87) );
  DFF_X1 inst1_KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S23reg_gff_1_SFF_2_n5), .CK(clk), .Q(inst1_n88) );
  DFF_X1 inst1_KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S23reg_gff_1_SFF_1_n5), .CK(clk), .Q(inst1_n89) );
  DFF_X1 inst1_KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S23reg_gff_1_SFF_0_n5), .CK(clk), .Q(inst1_n90) );
  DFF_X1 inst1_KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S22reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst1_n91) );
  DFF_X1 inst1_KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S22reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst1_n92) );
  DFF_X1 inst1_KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S22reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst1_n93) );
  DFF_X1 inst1_KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S22reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst1_n94) );
  DFF_X1 inst1_KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S22reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst1_n95) );
  DFF_X1 inst1_KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S22reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst1_n96) );
  DFF_X1 inst1_KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S22reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst1_n97) );
  DFF_X1 inst1_KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S22reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst1_n98) );
  DFF_X1 inst1_KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S21reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst1_n107) );
  DFF_X1 inst1_KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S21reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst1_n108) );
  DFF_X1 inst1_KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S21reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst1_n109) );
  DFF_X1 inst1_KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S21reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst1_n110) );
  DFF_X1 inst1_KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S21reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst1_n111) );
  DFF_X1 inst1_KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S21reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst1_n112) );
  DFF_X1 inst1_KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S21reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst1_n113) );
  DFF_X1 inst1_KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S21reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst1_n114) );
  DFF_X1 inst1_KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S20reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst1_n115) );
  DFF_X1 inst1_KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S20reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst1_n116) );
  DFF_X1 inst1_KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S20reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst1_n117) );
  DFF_X1 inst1_KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S20reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst1_n118) );
  DFF_X1 inst1_KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S20reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst1_n119) );
  DFF_X1 inst1_KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S20reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst1_n120) );
  DFF_X1 inst1_KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S20reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst1_n121) );
  DFF_X1 inst1_KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S20reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst1_n122), .QN(
        inst1_n1289) );
  DFF_X1 inst1_KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S13reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst1_n9), .QN(
        inst1_n1280) );
  DFF_X1 inst1_KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S13reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst1_n24), .QN(
        inst1_n1281) );
  DFF_X1 inst1_KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S13reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst1_n10), .QN(
        inst1_n1282) );
  DFF_X1 inst1_KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S13reg_gff_1_SFF_4_n5), .CK(clk), .Q(inst1_n11), .QN(
        inst1_n1283) );
  DFF_X1 inst1_KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S13reg_gff_1_SFF_3_n5), .CK(clk), .Q(inst1_n12), .QN(
        inst1_n1284) );
  DFF_X1 inst1_KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S13reg_gff_1_SFF_2_n5), .CK(clk), .Q(inst1_n14), .QN(
        inst1_n1285) );
  DFF_X1 inst1_KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S13reg_gff_1_SFF_1_n5), .CK(clk), .Q(inst1_n17), .QN(
        inst1_n1286) );
  DFF_X1 inst1_KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S13reg_gff_1_SFF_0_n5), .CK(clk), .Q(inst1_n22), .QN(
        inst1_n1287) );
  DFF_X1 inst1_KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S12reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst1_n123), .QN(
        inst1_n1290) );
  DFF_X1 inst1_KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S12reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst1_n124), .QN(
        inst1_n1291) );
  DFF_X1 inst1_KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S12reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst1_n125), .QN(
        inst1_n1292) );
  DFF_X1 inst1_KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S12reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst1_n126), .QN(
        inst1_n1293) );
  DFF_X1 inst1_KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S12reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst1_n127), .QN(
        inst1_n1294) );
  DFF_X1 inst1_KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S12reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst1_n128), .QN(
        inst1_n1295) );
  DFF_X1 inst1_KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S12reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst1_n129), .QN(
        inst1_n1296) );
  DFF_X1 inst1_KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S12reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst1_n130), .QN(
        inst1_n1297) );
  DFF_X1 inst1_KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S11reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst1_n131) );
  DFF_X1 inst1_KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S11reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst1_n132) );
  DFF_X1 inst1_KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S11reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst1_n133) );
  DFF_X1 inst1_KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S11reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst1_n134) );
  DFF_X1 inst1_KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S11reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst1_n135) );
  DFF_X1 inst1_KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S11reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst1_n136) );
  DFF_X1 inst1_KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S11reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst1_n137) );
  DFF_X1 inst1_KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S11reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst1_n980) );
  DFF_X1 inst1_KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S10reg_gff_1_SFF_7_n6), .CK(clk), .QN(inst1_n979) );
  DFF_X1 inst1_KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S10reg_gff_1_SFF_6_n6), .CK(clk), .QN(inst1_n978) );
  DFF_X1 inst1_KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S10reg_gff_1_SFF_5_n6), .CK(clk), .QN(inst1_n977) );
  DFF_X1 inst1_KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S10reg_gff_1_SFF_4_n6), .CK(clk), .QN(inst1_n976) );
  DFF_X1 inst1_KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S10reg_gff_1_SFF_3_n6), .CK(clk), .QN(inst1_n975) );
  DFF_X1 inst1_KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S10reg_gff_1_SFF_2_n6), .CK(clk), .QN(inst1_n974) );
  DFF_X1 inst1_KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S10reg_gff_1_SFF_1_n6), .CK(clk), .QN(inst1_n973) );
  DFF_X1 inst1_KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S10reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst1_n972) );
  DFF_X1 inst1_KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S03reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst1_n971) );
  DFF_X1 inst1_KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S03reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst1_n970) );
  DFF_X1 inst1_KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S03reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst1_n969) );
  DFF_X1 inst1_KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S03reg_gff_1_SFF_4_n5), .CK(clk), .QN(inst1_n968) );
  DFF_X1 inst1_KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S03reg_gff_1_SFF_3_n5), .CK(clk), .QN(inst1_n967) );
  DFF_X1 inst1_KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S03reg_gff_1_SFF_2_n5), .CK(clk), .QN(inst1_n966) );
  DFF_X1 inst1_KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S03reg_gff_1_SFF_1_n5), .CK(clk), .QN(inst1_n965) );
  DFF_X1 inst1_KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S03reg_gff_1_SFF_0_n5), .CK(clk), .QN(inst1_n964) );
  DFF_X1 inst1_KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S02reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst1_n963) );
  DFF_X1 inst1_KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S02reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst1_n962) );
  DFF_X1 inst1_KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S02reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst1_n961) );
  DFF_X1 inst1_KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S02reg_gff_1_SFF_4_n6), .CK(clk), .QN(inst1_n960) );
  DFF_X1 inst1_KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S02reg_gff_1_SFF_3_n6), .CK(clk), .QN(inst1_n959) );
  DFF_X1 inst1_KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S02reg_gff_1_SFF_2_n6), .CK(clk), .QN(inst1_n958) );
  DFF_X1 inst1_KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S02reg_gff_1_SFF_1_n6), .CK(clk), .QN(inst1_n957) );
  DFF_X1 inst1_KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S02reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst1_n956) );
  DFF_X1 inst1_KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S01reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst1_n1265), .QN(
        inst1_n955) );
  DFF_X1 inst1_KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S01reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst1_n1266), .QN(
        inst1_n954) );
  DFF_X1 inst1_KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S01reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst1_n1267), .QN(
        inst1_n953) );
  DFF_X1 inst1_KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S01reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst1_n1268), .QN(
        inst1_n952) );
  DFF_X1 inst1_KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S01reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst1_n1269), .QN(
        inst1_n951) );
  DFF_X1 inst1_KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S01reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst1_n1270), .QN(
        inst1_n950) );
  DFF_X1 inst1_KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S01reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst1_n1271), .QN(
        inst1_n949) );
  DFF_X1 inst1_KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S01reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst1_n948) );
  DFF_X1 inst1_KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S00reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst1_n1243), .QN(
        inst1_n1091) );
  DFF_X1 inst1_KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S00reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst1_n1244), .QN(
        inst1_n1090) );
  DFF_X1 inst1_KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S00reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst1_n1245), .QN(
        inst1_n1084) );
  DFF_X1 inst1_KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S00reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst1_n1246), .QN(
        inst1_n1089) );
  DFF_X1 inst1_KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S00reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst1_n1247), .QN(
        inst1_n1088) );
  DFF_X1 inst1_KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S00reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst1_n1242), .QN(
        inst1_n1087) );
  DFF_X1 inst1_KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S00reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst1_n1241), .QN(
        inst1_n1086) );
  DFF_X1 inst1_KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_KeyArray_S00reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst1_n1248), .QN(
        inst1_n1085) );
  DFF_X1 inst1_stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S33reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext1[7]),
        .QN(inst1_n947) );
  DFF_X1 inst1_stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S33reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext1[6]),
        .QN(inst1_n946) );
  DFF_X1 inst1_stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S33reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext1[5]),
        .QN(inst1_n945) );
  DFF_X1 inst1_stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S33reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext1[4]),
        .QN(inst1_n944) );
  DFF_X1 inst1_stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S33reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext1[3]),
        .QN(inst1_n943) );
  DFF_X1 inst1_stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S33reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext1[2]),
        .QN(inst1_n942) );
  DFF_X1 inst1_stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S33reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext1[1]),
        .QN(inst1_n941) );
  DFF_X1 inst1_stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S33reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext1[0]),
        .QN(inst1_n940) );
  DFF_X1 inst1_stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S32reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext1[15]),
        .QN(inst1_n939) );
  DFF_X1 inst1_stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S32reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext1[14]),
        .QN(inst1_n938) );
  DFF_X1 inst1_stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S32reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext1[13]),
        .QN(inst1_n937) );
  DFF_X1 inst1_stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S32reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[12]),
        .QN(inst1_n936) );
  DFF_X1 inst1_stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S32reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[11]),
        .QN(inst1_n935) );
  DFF_X1 inst1_stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S32reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[10]),
        .QN(inst1_n934) );
  DFF_X1 inst1_stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S32reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[9]),
        .QN(inst1_n933) );
  DFF_X1 inst1_stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S32reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[8]),
        .QN(inst1_n932) );
  DFF_X1 inst1_stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S31reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext1[23]),
        .QN(inst1_n1252) );
  DFF_X1 inst1_stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S31reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext1[22]),
        .QN(inst1_n1251) );
  DFF_X1 inst1_stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S31reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext1[21]),
        .QN(inst1_n1253) );
  DFF_X1 inst1_stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S31reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[20]),
        .QN(inst1_n1254) );
  DFF_X1 inst1_stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S31reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[19]),
        .QN(inst1_n1255) );
  DFF_X1 inst1_stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S31reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[18]),
        .QN(inst1_n1256) );
  DFF_X1 inst1_stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S31reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[17]),
        .QN(inst1_n1257) );
  DFF_X1 inst1_stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S31reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[16]),
        .QN(inst1_n1258) );
  DFF_X1 inst1_stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S30reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext1[31]),
        .QN(inst1_n1230) );
  DFF_X1 inst1_stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S30reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext1[30]),
        .QN(inst1_n1097) );
  DFF_X1 inst1_stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S30reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext1[29]),
        .QN(inst1_n1229) );
  DFF_X1 inst1_stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S30reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext1[28]),
        .QN(inst1_n1105) );
  DFF_X1 inst1_stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S30reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext1[27]),
        .QN(inst1_n1231) );
  DFF_X1 inst1_stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S30reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext1[26]),
        .QN(inst1_n1109) );
  DFF_X1 inst1_stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S30reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext1[25]),
        .QN(inst1_n1121) );
  DFF_X1 inst1_stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S30reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext1[24]),
        .QN(inst1_n1113) );
  DFF_X1 inst1_stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S23reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext1[39]),
        .QN(inst1_n923) );
  DFF_X1 inst1_stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S23reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext1[38]),
        .QN(inst1_n922) );
  DFF_X1 inst1_stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S23reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext1[37]),
        .QN(inst1_n921) );
  DFF_X1 inst1_stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S23reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[36]),
        .QN(inst1_n920) );
  DFF_X1 inst1_stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S23reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[35]),
        .QN(inst1_n919) );
  DFF_X1 inst1_stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S23reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[34]),
        .QN(inst1_n918) );
  DFF_X1 inst1_stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S23reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[33]),
        .QN(inst1_n917) );
  DFF_X1 inst1_stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S23reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[32]),
        .QN(inst1_n916) );
  DFF_X1 inst1_stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S22reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext1[47]),
        .QN(inst1_n915) );
  DFF_X1 inst1_stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S22reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext1[46]),
        .QN(inst1_n914) );
  DFF_X1 inst1_stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S22reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext1[45]),
        .QN(inst1_n913) );
  DFF_X1 inst1_stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S22reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[44]),
        .QN(inst1_n912) );
  DFF_X1 inst1_stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S22reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[43]),
        .QN(inst1_n911) );
  DFF_X1 inst1_stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S22reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[42]),
        .QN(inst1_n910) );
  DFF_X1 inst1_stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S22reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[41]),
        .QN(inst1_n909) );
  DFF_X1 inst1_stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S22reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[40]),
        .QN(inst1_n908) );
  DFF_X1 inst1_stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S21reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext1[55])
         );
  DFF_X1 inst1_stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S21reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext1[54])
         );
  DFF_X1 inst1_stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S21reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext1[53])
         );
  DFF_X1 inst1_stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S21reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[52])
         );
  DFF_X1 inst1_stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S21reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[51])
         );
  DFF_X1 inst1_stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S21reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[50])
         );
  DFF_X1 inst1_stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S21reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[49])
         );
  DFF_X1 inst1_stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S21reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[48])
         );
  DFF_X1 inst1_stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S20reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext1[63]),
        .QN(inst1_n1093) );
  DFF_X1 inst1_stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S20reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext1[62]),
        .QN(inst1_n1232) );
  DFF_X1 inst1_stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S20reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext1[61]),
        .QN(inst1_n1249) );
  DFF_X1 inst1_stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S20reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext1[60]),
        .QN(inst1_n1234) );
  DFF_X1 inst1_stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S20reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext1[59]),
        .QN(inst1_n1116) );
  DFF_X1 inst1_stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S20reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext1[58]),
        .QN(inst1_n1119) );
  DFF_X1 inst1_stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S20reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext1[57]),
        .QN(inst1_n1235) );
  DFF_X1 inst1_stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S20reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext1[56]),
        .QN(inst1_n1233) );
  DFF_X1 inst1_stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S13reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext1[71])
         );
  DFF_X1 inst1_stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S13reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext1[70])
         );
  DFF_X1 inst1_stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S13reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext1[69])
         );
  DFF_X1 inst1_stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S13reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[68])
         );
  DFF_X1 inst1_stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S13reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[67])
         );
  DFF_X1 inst1_stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S13reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[66])
         );
  DFF_X1 inst1_stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S13reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[65])
         );
  DFF_X1 inst1_stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S13reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[64])
         );
  DFF_X1 inst1_stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S12reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext1[79]),
        .QN(inst1_n891) );
  DFF_X1 inst1_stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S12reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext1[78]),
        .QN(inst1_n890) );
  DFF_X1 inst1_stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S12reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext1[77]),
        .QN(inst1_n889) );
  DFF_X1 inst1_stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S12reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[76]),
        .QN(inst1_n888) );
  DFF_X1 inst1_stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S12reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[75]),
        .QN(inst1_n887) );
  DFF_X1 inst1_stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S12reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[74]),
        .QN(inst1_n886) );
  DFF_X1 inst1_stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S12reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[73]),
        .QN(inst1_n885) );
  DFF_X1 inst1_stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S12reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[72]),
        .QN(inst1_n884) );
  DFF_X1 inst1_stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S11reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext1[87]),
        .QN(inst1_n883) );
  DFF_X1 inst1_stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S11reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext1[86]),
        .QN(inst1_n882) );
  DFF_X1 inst1_stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S11reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext1[85]),
        .QN(inst1_n881) );
  DFF_X1 inst1_stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S11reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[84]),
        .QN(inst1_n880) );
  DFF_X1 inst1_stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S11reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[83]),
        .QN(inst1_n879) );
  DFF_X1 inst1_stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S11reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[82]),
        .QN(inst1_n878) );
  DFF_X1 inst1_stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S11reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[81]),
        .QN(inst1_n877) );
  DFF_X1 inst1_stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S11reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[80]),
        .QN(inst1_n876) );
  DFF_X1 inst1_stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S10reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext1[95]),
        .QN(inst1_n1092) );
  DFF_X1 inst1_stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S10reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext1[94]),
        .QN(inst1_n1106) );
  DFF_X1 inst1_stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S10reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext1[93]),
        .QN(inst1_n1122) );
  DFF_X1 inst1_stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S10reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext1[92]),
        .QN(inst1_n1100) );
  DFF_X1 inst1_stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S10reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext1[91]),
        .QN(inst1_n1111) );
  DFF_X1 inst1_stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S10reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext1[90]),
        .QN(inst1_n1118) );
  DFF_X1 inst1_stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S10reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext1[89]),
        .QN(inst1_n1115) );
  DFF_X1 inst1_stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S10reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext1[88]),
        .QN(inst1_n1103) );
  DFF_X1 inst1_stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S03reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext1[103]), .QN(inst1_n875) );
  DFF_X1 inst1_stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S03reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext1[102]), .QN(inst1_n874) );
  DFF_X1 inst1_stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S03reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext1[101]), .QN(inst1_n873) );
  DFF_X1 inst1_stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S03reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[100]), .QN(inst1_n872) );
  DFF_X1 inst1_stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S03reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[99]),
        .QN(inst1_n871) );
  DFF_X1 inst1_stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S03reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[98]),
        .QN(inst1_n870) );
  DFF_X1 inst1_stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S03reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[97]),
        .QN(inst1_n869) );
  DFF_X1 inst1_stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S03reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[96]),
        .QN(inst1_n868) );
  DFF_X1 inst1_stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S02reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext1[111]) );
  DFF_X1 inst1_stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S02reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext1[110]) );
  DFF_X1 inst1_stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S02reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext1[109]) );
  DFF_X1 inst1_stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S02reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[108]) );
  DFF_X1 inst1_stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S02reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[107]) );
  DFF_X1 inst1_stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S02reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[106]) );
  DFF_X1 inst1_stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S02reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[105]) );
  DFF_X1 inst1_stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S02reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[104]) );
  DFF_X1 inst1_stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S01reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext1[119]), .QN(inst1_n1272) );
  DFF_X1 inst1_stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S01reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext1[118]), .QN(inst1_n1273) );
  DFF_X1 inst1_stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S01reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext1[117]), .QN(inst1_n1274) );
  DFF_X1 inst1_stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S01reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[116]), .QN(inst1_n1275) );
  DFF_X1 inst1_stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S01reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[115]), .QN(inst1_n1276) );
  DFF_X1 inst1_stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S01reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[114]), .QN(inst1_n1277) );
  DFF_X1 inst1_stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S01reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[113]), .QN(inst1_n1278) );
  DFF_X1 inst1_stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S01reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[112]), .QN(inst1_n1279) );
  DFF_X1 inst1_stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst1_stateArray_S00reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext1[127]), .QN(inst1_n1094) );
  DFF_X1 inst1_stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst1_stateArray_S00reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext1[126]), .QN(inst1_n1096) );
  DFF_X1 inst1_stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst1_stateArray_S00reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext1[125]), .QN(inst1_n1098) );
  DFF_X1 inst1_stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst1_stateArray_S00reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext1[124]), .QN(inst1_n1225) );
  DFF_X1 inst1_stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst1_stateArray_S00reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext1[123]), .QN(inst1_n1110) );
  DFF_X1 inst1_stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst1_stateArray_S00reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext1[122]), .QN(inst1_n1227) );
  DFF_X1 inst1_stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst1_stateArray_S00reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext1[121]), .QN(inst1_n1114) );
  DFF_X1 inst1_stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst1_stateArray_S00reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext1[120]), .QN(inst1_n1102) );
  DFF_X1 inst1_ctrl_CSenRC_reg_FF_FF ( .D(inst1_n827), .CK(clk), .QN(
        inst1_n1076) );
  DFF_X1 inst1_ctrl_CSselMC_reg_FF_FF ( .D(inst1_n1188), .CK(clk), .Q(
        inst1_ctrl_n6) );
  DFF_X1 inst1_ctrl_seq4_SFF_1_Q_reg_FF_FF ( .D(inst1_ctrl_seq4_SFF_1_n5),
        .CK(clk), .Q(inst1_n1250), .QN(inst1_n1077) );
  DFF_X1 inst1_ctrl_seq4_SFF_0_Q_reg_FF_FF ( .D(inst1_ctrl_seq4_SFF_0_n5),
        .CK(clk), .Q(inst1_n143), .QN(inst1_n1236) );
  DFF_X1 inst1_ctrl_seq6_SFF_4_Q_reg_FF_FF ( .D(inst1_ctrl_seq6_SFF_4_n5),
        .CK(clk), .QN(inst1_n851) );
  DFF_X1 inst1_ctrl_seq6_SFF_3_Q_reg_FF_FF ( .D(inst1_ctrl_seq6_SFF_3_n5),
        .CK(clk), .QN(inst1_n1081) );
  DFF_X1 inst1_ctrl_seq6_SFF_2_Q_reg_FF_FF ( .D(inst1_ctrl_seq6_SFF_2_n5),
        .CK(clk), .QN(inst1_n1079) );
  DFF_X1 inst1_ctrl_seq6_SFF_1_Q_reg_FF_FF ( .D(inst1_ctrl_seq6_SFF_1_n5),
        .CK(clk), .QN(inst1_n1082) );
  DFF_X1 inst1_ctrl_seq6_SFF_0_Q_reg_FF_FF ( .D(inst1_ctrl_seq6_SFF_0_n5),
        .CK(clk), .QN(inst1_n1080) );
  OAI21_X1 inst2_U1161 ( .B1(inst2_n2798), .B2(inst2_n2797), .A(inst2_n2796),
        .ZN(inst2_n1088) );
  NOR2_X1 inst2_U1160 ( .A1(inst2_n143), .A2(inst2_n2826), .ZN(inst2_n2798) );
  OAI211_X1 inst2_U1159 ( .C1(inst2_n2795), .C2(inst2_n2794), .A(inst2_n2793),
        .B(inst2_n2792), .ZN(inst2_stateArray_S23reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst2_U1158 ( .B1(inst2_n2791), .B2(ciphertext2[49]), .A(
        inst2_n2790), .ZN(inst2_n2792) );
  OAI22_X1 inst2_U1157 ( .A1(inst2_n191), .A2(inst2_n2776), .B1(inst2_n2789),
        .B2(inst2_n2810), .ZN(inst2_n2790) );
  AOI22_X1 inst2_U1156 ( .A1(inst2_n2788), .A2(ciphertext2[33]), .B1(
        plaintext2[33]), .B2(inst2_n2803), .ZN(inst2_n2793) );
  XNOR2_X1 inst2_U1155 ( .A(inst2_n2787), .B(inst2_n2786), .ZN(inst2_n2795) );
  AOI22_X1 inst2_U1154 ( .A1(inst2_n191), .A2(inst2_n2785), .B1(inst2_n2784),
        .B2(ciphertext2[25]), .ZN(inst2_n2786) );
  XNOR2_X1 inst2_U1153 ( .A(inst2_n2783), .B(inst2_n2782), .ZN(inst2_n2787) );
  OAI211_X1 inst2_U1152 ( .C1(inst2_n2781), .C2(inst2_n2780), .A(inst2_n2779),
        .B(inst2_n2778), .ZN(inst2_stateArray_S23reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst2_U1151 ( .B1(inst2_n2791), .B2(ciphertext2[50]), .A(
        inst2_n2777), .ZN(inst2_n2778) );
  OAI22_X1 inst2_U1150 ( .A1(inst2_n203), .A2(inst2_n2776), .B1(inst2_n193),
        .B2(inst2_n2789), .ZN(inst2_n2777) );
  AOI22_X1 inst2_U1149 ( .A1(inst2_n2788), .A2(ciphertext2[34]), .B1(
        plaintext2[34]), .B2(inst2_n2803), .ZN(inst2_n2779) );
  XNOR2_X1 inst2_U1148 ( .A(inst2_n2775), .B(inst2_n2774), .ZN(inst2_n2781) );
  AOI22_X1 inst2_U1147 ( .A1(inst2_n203), .A2(inst2_n2773), .B1(inst2_n2772),
        .B2(ciphertext2[26]), .ZN(inst2_n2774) );
  NOR2_X1 inst2_U1146 ( .A1(inst2_n2771), .A2(inst2_n2811), .ZN(
        inst2_ctrl_seq4_SFF_1_n5) );
  NOR2_X1 inst2_U1145 ( .A1(inst2_n232), .A2(inst2_n2713), .ZN(
        inst2_ctrl_seq6_SFF_1_n5) );
  NOR2_X1 inst2_U1144 ( .A1(inst2_n233), .A2(inst2_n2582), .ZN(
        inst2_ctrl_seq6_SFF_3_n5) );
  OAI211_X1 inst2_U1143 ( .C1(inst2_n2794), .C2(inst2_n2770), .A(inst2_n2769),
        .B(inst2_n2768), .ZN(inst2_stateArray_S23reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst2_U1142 ( .B1(inst2_n2791), .B2(ciphertext2[52]), .A(
        inst2_n2767), .ZN(inst2_n2768) );
  OAI22_X1 inst2_U1141 ( .A1(inst2_n207), .A2(inst2_n2776), .B1(inst2_n2789),
        .B2(inst2_n2809), .ZN(inst2_n2767) );
  AOI22_X1 inst2_U1140 ( .A1(inst2_n2788), .A2(ciphertext2[36]), .B1(
        plaintext2[36]), .B2(inst2_n2803), .ZN(inst2_n2769) );
  XNOR2_X1 inst2_U1139 ( .A(inst2_n2766), .B(inst2_n2765), .ZN(inst2_n2770) );
  AOI22_X1 inst2_U1138 ( .A1(inst2_n212), .A2(inst2_n2764), .B1(inst2_n2763),
        .B2(ciphertext2[92]), .ZN(inst2_n2765) );
  AOI22_X1 inst2_U1137 ( .A1(inst2_n2785), .A2(inst2_n2762), .B1(inst2_n2761),
        .B2(inst2_n2784), .ZN(inst2_n2766) );
  OAI22_X1 inst2_U1136 ( .A1(inst2_n1080), .A2(inst2_n2760), .B1(inst2_n718),
        .B2(inst2_n2759), .ZN(inst2_calcRCon_n45) );
  OAI21_X1 inst2_U1135 ( .B1(inst2_n499), .B2(inst2_n2759), .A(inst2_n2758),
        .ZN(inst2_calcRCon_n50) );
  OAI221_X1 inst2_U1134 ( .B1(inst2_n1071), .B2(inst2_n444), .C1(inst2_n2801),
        .C2(inst2_n2837), .A(inst2_n2791), .ZN(inst2_n2758) );
  OAI22_X1 inst2_U1133 ( .A1(inst2_n1080), .A2(inst2_n2759), .B1(inst2_n1081),
        .B2(inst2_n2757), .ZN(inst2_calcRCon_n46) );
  OAI21_X1 inst2_U1132 ( .B1(inst2_n1081), .B2(inst2_n2759), .A(inst2_n2756),
        .ZN(inst2_calcRCon_n47) );
  OAI221_X1 inst2_U1131 ( .B1(inst2_n706), .B2(inst2_n1071), .C1(inst2_n2812),
        .C2(inst2_n2801), .A(inst2_n2791), .ZN(inst2_n2756) );
  NAND2_X1 inst2_U1130 ( .A1(inst2_n6), .A2(inst2_n2757), .ZN(inst2_n2759) );
  OAI211_X1 inst2_U1129 ( .C1(inst2_n1233), .C2(inst2_n2760), .A(inst2_n2755),
        .B(inst2_n2754), .ZN(inst2_stateArray_S20reg_gff_1_SFF_0_n5) );
  NAND2_X1 inst2_U1128 ( .A1(inst2_n1917), .A2(ciphertext2[48]), .ZN(
        inst2_n2754) );
  AOI22_X1 inst2_U1127 ( .A1(ciphertext2[56]), .A2(done2), .B1(plaintext2[56]),
        .B2(inst2_n2803), .ZN(inst2_n2755) );
  OAI211_X1 inst2_U1126 ( .C1(inst2_n1232), .C2(inst2_n2760), .A(inst2_n2753),
        .B(inst2_n2752), .ZN(inst2_stateArray_S20reg_gff_1_SFF_1_n5) );
  NAND2_X1 inst2_U1125 ( .A1(inst2_n1917), .A2(ciphertext2[49]), .ZN(
        inst2_n2752) );
  AOI22_X1 inst2_U1124 ( .A1(ciphertext2[57]), .A2(done2), .B1(plaintext2[57]),
        .B2(inst2_n2803), .ZN(inst2_n2753) );
  OAI211_X1 inst2_U1123 ( .C1(inst2_n1231), .C2(inst2_n2760), .A(inst2_n2751),
        .B(inst2_n2750), .ZN(inst2_stateArray_S20reg_gff_1_SFF_2_n5) );
  NAND2_X1 inst2_U1122 ( .A1(inst2_n1917), .A2(ciphertext2[50]), .ZN(
        inst2_n2750) );
  AOI22_X1 inst2_U1121 ( .A1(inst2_n2788), .A2(ciphertext2[58]), .B1(
        plaintext2[58]), .B2(inst2_n2803), .ZN(inst2_n2751) );
  OAI211_X1 inst2_U1120 ( .C1(inst2_n1230), .C2(inst2_n2760), .A(inst2_n2749),
        .B(inst2_n2748), .ZN(inst2_stateArray_S20reg_gff_1_SFF_3_n5) );
  NAND2_X1 inst2_U1119 ( .A1(inst2_n1917), .A2(ciphertext2[51]), .ZN(
        inst2_n2748) );
  AOI22_X1 inst2_U1118 ( .A1(inst2_n2788), .A2(ciphertext2[59]), .B1(
        plaintext2[59]), .B2(inst2_n2803), .ZN(inst2_n2749) );
  OAI211_X1 inst2_U1117 ( .C1(inst2_n1229), .C2(inst2_n2760), .A(inst2_n2747),
        .B(inst2_n2746), .ZN(inst2_stateArray_S20reg_gff_1_SFF_4_n5) );
  NAND2_X1 inst2_U1116 ( .A1(inst2_n1917), .A2(ciphertext2[52]), .ZN(
        inst2_n2746) );
  AOI22_X1 inst2_U1115 ( .A1(ciphertext2[60]), .A2(done2), .B1(plaintext2[60]),
        .B2(inst2_n2803), .ZN(inst2_n2747) );
  OAI211_X1 inst2_U1114 ( .C1(inst2_n1228), .C2(inst2_n2757), .A(inst2_n2745),
        .B(inst2_n2744), .ZN(inst2_stateArray_S20reg_gff_1_SFF_5_n5) );
  NAND2_X1 inst2_U1113 ( .A1(inst2_n1917), .A2(ciphertext2[53]), .ZN(
        inst2_n2744) );
  AOI22_X1 inst2_U1112 ( .A1(ciphertext2[61]), .A2(done2), .B1(plaintext2[61]),
        .B2(inst2_n2803), .ZN(inst2_n2745) );
  OAI211_X1 inst2_U1111 ( .C1(inst2_n1227), .C2(inst2_n2760), .A(inst2_n2743),
        .B(inst2_n2742), .ZN(inst2_stateArray_S20reg_gff_1_SFF_6_n5) );
  NAND2_X1 inst2_U1110 ( .A1(inst2_n1917), .A2(ciphertext2[54]), .ZN(
        inst2_n2742) );
  AOI22_X1 inst2_U1109 ( .A1(ciphertext2[62]), .A2(done2), .B1(plaintext2[62]),
        .B2(inst2_n2803), .ZN(inst2_n2743) );
  OAI211_X1 inst2_U1108 ( .C1(inst2_n1226), .C2(inst2_n2757), .A(inst2_n2741),
        .B(inst2_n2740), .ZN(inst2_stateArray_S20reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst2_U1107 ( .A1(inst2_n1917), .A2(ciphertext2[55]), .ZN(
        inst2_n2740) );
  AOI22_X1 inst2_U1106 ( .A1(inst2_n2788), .A2(ciphertext2[63]), .B1(
        plaintext2[63]), .B2(inst2_n2803), .ZN(inst2_n2741) );
  OAI211_X1 inst2_U1105 ( .C1(inst2_n1233), .C2(inst2_n2771), .A(inst2_n2739),
        .B(inst2_n2738), .ZN(inst2_stateArray_S21reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst2_U1104 ( .A1(plaintext2[48]), .A2(inst2_n2713), .ZN(
        inst2_n2738) );
  AOI22_X1 inst2_U1103 ( .A1(inst2_n2788), .A2(ciphertext2[48]), .B1(
        inst2_n2791), .B2(ciphertext2[32]), .ZN(inst2_n2739) );
  OAI211_X1 inst2_U1102 ( .C1(inst2_n1232), .C2(inst2_n2771), .A(inst2_n2737),
        .B(inst2_n2736), .ZN(inst2_stateArray_S21reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst2_U1101 ( .A1(plaintext2[49]), .A2(inst2_n2550), .ZN(
        inst2_n2736) );
  AOI22_X1 inst2_U1100 ( .A1(inst2_n2788), .A2(ciphertext2[49]), .B1(
        inst2_n2791), .B2(ciphertext2[33]), .ZN(inst2_n2737) );
  OAI211_X1 inst2_U1099 ( .C1(inst2_n1231), .C2(inst2_n2771), .A(inst2_n2735),
        .B(inst2_n2734), .ZN(inst2_stateArray_S21reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst2_U1098 ( .A1(plaintext2[50]), .A2(inst2_n2595), .ZN(
        inst2_n2734) );
  AOI22_X1 inst2_U1097 ( .A1(done2), .A2(ciphertext2[50]), .B1(inst2_n2791),
        .B2(ciphertext2[34]), .ZN(inst2_n2735) );
  OAI211_X1 inst2_U1096 ( .C1(inst2_n1230), .C2(inst2_n2771), .A(inst2_n2733),
        .B(inst2_n2732), .ZN(inst2_stateArray_S21reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst2_U1095 ( .A1(plaintext2[51]), .A2(inst2_n2722), .ZN(
        inst2_n2732) );
  AOI22_X1 inst2_U1094 ( .A1(done2), .A2(ciphertext2[51]), .B1(inst2_n2791),
        .B2(ciphertext2[35]), .ZN(inst2_n2733) );
  OAI211_X1 inst2_U1093 ( .C1(inst2_n1229), .C2(inst2_n2771), .A(inst2_n2731),
        .B(inst2_n2730), .ZN(inst2_stateArray_S21reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst2_U1092 ( .A1(plaintext2[52]), .A2(inst2_n2713), .ZN(
        inst2_n2730) );
  AOI22_X1 inst2_U1091 ( .A1(done2), .A2(ciphertext2[52]), .B1(inst2_n2791),
        .B2(ciphertext2[36]), .ZN(inst2_n2731) );
  OAI211_X1 inst2_U1090 ( .C1(inst2_n1228), .C2(inst2_n2771), .A(inst2_n2729),
        .B(inst2_n2728), .ZN(inst2_stateArray_S21reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst2_U1089 ( .A1(plaintext2[53]), .A2(inst2_n2484), .ZN(
        inst2_n2728) );
  AOI22_X1 inst2_U1088 ( .A1(done2), .A2(ciphertext2[53]), .B1(inst2_n2791),
        .B2(ciphertext2[37]), .ZN(inst2_n2729) );
  OAI211_X1 inst2_U1087 ( .C1(inst2_n1227), .C2(inst2_n2771), .A(inst2_n2727),
        .B(inst2_n2726), .ZN(inst2_stateArray_S21reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst2_U1086 ( .A1(plaintext2[54]), .A2(inst2_n2713), .ZN(
        inst2_n2726) );
  AOI22_X1 inst2_U1085 ( .A1(done2), .A2(ciphertext2[54]), .B1(inst2_n2791),
        .B2(ciphertext2[38]), .ZN(inst2_n2727) );
  OAI211_X1 inst2_U1084 ( .C1(inst2_n1226), .C2(inst2_n2771), .A(inst2_n2725),
        .B(inst2_n2724), .ZN(inst2_stateArray_S21reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst2_U1083 ( .A1(plaintext2[55]), .A2(inst2_n2657), .ZN(
        inst2_n2724) );
  AOI22_X1 inst2_U1082 ( .A1(done2), .A2(ciphertext2[55]), .B1(inst2_n2791),
        .B2(ciphertext2[39]), .ZN(inst2_n2725) );
  OAI21_X1 inst2_U1081 ( .B1(inst2_n1221), .B2(inst2_n2771), .A(inst2_n2723),
        .ZN(inst2_stateArray_S22reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst2_U1080 ( .B1(plaintext2[44]), .B2(inst2_n2722), .A(inst2_n2721), .ZN(inst2_n2723) );
  OAI22_X1 inst2_U1079 ( .A1(inst2_n1229), .A2(inst2_n2711), .B1(inst2_n2760),
        .B2(inst2_n2809), .ZN(inst2_n2721) );
  OAI21_X1 inst2_U1078 ( .B1(inst2_n2771), .B2(inst2_n2835), .A(inst2_n2720),
        .ZN(inst2_stateArray_S30reg_gff_1_SFF_0_n5) );
  AOI21_X1 inst2_U1077 ( .B1(plaintext2[24]), .B2(inst2_n2722), .A(inst2_n2719), .ZN(inst2_n2720) );
  OAI22_X1 inst2_U1076 ( .A1(inst2_n199), .A2(inst2_n2711), .B1(inst2_n1201),
        .B2(inst2_n2757), .ZN(inst2_n2719) );
  OAI21_X1 inst2_U1075 ( .B1(inst2_n2771), .B2(inst2_n2834), .A(inst2_n2718),
        .ZN(inst2_stateArray_S30reg_gff_1_SFF_1_n5) );
  AOI21_X1 inst2_U1074 ( .B1(plaintext2[25]), .B2(inst2_n2722), .A(inst2_n2717), .ZN(inst2_n2718) );
  OAI22_X1 inst2_U1073 ( .A1(inst2_n191), .A2(inst2_n2711), .B1(inst2_n1200),
        .B2(inst2_n2757), .ZN(inst2_n2717) );
  OAI21_X1 inst2_U1072 ( .B1(inst2_n2771), .B2(inst2_n2833), .A(inst2_n2716),
        .ZN(inst2_stateArray_S30reg_gff_1_SFF_2_n5) );
  AOI21_X1 inst2_U1071 ( .B1(plaintext2[26]), .B2(inst2_n2484), .A(inst2_n2715), .ZN(inst2_n2716) );
  OAI22_X1 inst2_U1070 ( .A1(inst2_n203), .A2(inst2_n2711), .B1(inst2_n1199),
        .B2(inst2_n2757), .ZN(inst2_n2715) );
  OAI21_X1 inst2_U1069 ( .B1(inst2_n2771), .B2(inst2_n2832), .A(inst2_n2714),
        .ZN(inst2_stateArray_S30reg_gff_1_SFF_3_n5) );
  AOI21_X1 inst2_U1068 ( .B1(plaintext2[27]), .B2(inst2_n2713), .A(inst2_n2712), .ZN(inst2_n2714) );
  OAI22_X1 inst2_U1067 ( .A1(inst2_n1198), .A2(inst2_n2760), .B1(inst2_n2711),
        .B2(inst2_n2806), .ZN(inst2_n2712) );
  OAI21_X1 inst2_U1066 ( .B1(inst2_n2771), .B2(inst2_n2831), .A(inst2_n2710),
        .ZN(inst2_stateArray_S30reg_gff_1_SFF_4_n5) );
  AOI21_X1 inst2_U1065 ( .B1(plaintext2[28]), .B2(inst2_n2722), .A(inst2_n2709), .ZN(inst2_n2710) );
  OAI22_X1 inst2_U1064 ( .A1(inst2_n207), .A2(inst2_n2711), .B1(inst2_n1197),
        .B2(inst2_n2757), .ZN(inst2_n2709) );
  OAI21_X1 inst2_U1063 ( .B1(inst2_n2771), .B2(inst2_n2830), .A(inst2_n2708),
        .ZN(inst2_stateArray_S30reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst2_U1062 ( .B1(plaintext2[29]), .B2(inst2_n2713), .A(inst2_n2707), .ZN(inst2_n2708) );
  OAI22_X1 inst2_U1061 ( .A1(inst2_n1196), .A2(inst2_n2760), .B1(inst2_n2711),
        .B2(inst2_n2804), .ZN(inst2_n2707) );
  OAI21_X1 inst2_U1060 ( .B1(inst2_n2771), .B2(inst2_n2827), .A(inst2_n2706),
        .ZN(inst2_stateArray_S30reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst2_U1059 ( .B1(plaintext2[30]), .B2(inst2_n2722), .A(inst2_n2705), .ZN(inst2_n2706) );
  OAI22_X1 inst2_U1058 ( .A1(inst2_n215), .A2(inst2_n2711), .B1(inst2_n1195),
        .B2(inst2_n2757), .ZN(inst2_n2705) );
  OAI21_X1 inst2_U1057 ( .B1(inst2_n2771), .B2(inst2_n2829), .A(inst2_n2704),
        .ZN(inst2_stateArray_S30reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst2_U1056 ( .B1(plaintext2[31]), .B2(inst2_n2713), .A(inst2_n2703), .ZN(inst2_n2704) );
  OAI22_X1 inst2_U1055 ( .A1(inst2_n1194), .A2(inst2_n2760), .B1(inst2_n2711),
        .B2(inst2_n2805), .ZN(inst2_n2703) );
  OAI21_X1 inst2_U1054 ( .B1(inst2_n1201), .B2(inst2_n2771), .A(inst2_n2702),
        .ZN(inst2_stateArray_S32reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst2_U1053 ( .B1(plaintext2[8]), .B2(inst2_n2722), .A(inst2_n2701),
        .ZN(inst2_n2702) );
  OAI22_X1 inst2_U1052 ( .A1(inst2_n1209), .A2(inst2_n2711), .B1(inst2_n2760),
        .B2(inst2_n2835), .ZN(inst2_n2701) );
  OAI21_X1 inst2_U1051 ( .B1(inst2_n1200), .B2(inst2_n2771), .A(inst2_n2700),
        .ZN(inst2_stateArray_S32reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst2_U1050 ( .B1(plaintext2[9]), .B2(inst2_n2713), .A(inst2_n2699),
        .ZN(inst2_n2700) );
  OAI22_X1 inst2_U1049 ( .A1(inst2_n1208), .A2(inst2_n2711), .B1(inst2_n2757),
        .B2(inst2_n2834), .ZN(inst2_n2699) );
  OAI21_X1 inst2_U1048 ( .B1(inst2_n1199), .B2(inst2_n2771), .A(inst2_n2698),
        .ZN(inst2_stateArray_S32reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst2_U1047 ( .B1(plaintext2[10]), .B2(inst2_n2722), .A(inst2_n2697), .ZN(inst2_n2698) );
  OAI22_X1 inst2_U1046 ( .A1(inst2_n1207), .A2(inst2_n2711), .B1(inst2_n2757),
        .B2(inst2_n2833), .ZN(inst2_n2697) );
  OAI21_X1 inst2_U1045 ( .B1(inst2_n1198), .B2(inst2_n2771), .A(inst2_n2696),
        .ZN(inst2_stateArray_S32reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst2_U1044 ( .B1(plaintext2[11]), .B2(inst2_n2713), .A(inst2_n2695), .ZN(inst2_n2696) );
  OAI22_X1 inst2_U1043 ( .A1(inst2_n1206), .A2(inst2_n2711), .B1(inst2_n2757),
        .B2(inst2_n2832), .ZN(inst2_n2695) );
  OAI21_X1 inst2_U1042 ( .B1(inst2_n1197), .B2(inst2_n2771), .A(inst2_n2694),
        .ZN(inst2_stateArray_S32reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst2_U1041 ( .B1(plaintext2[12]), .B2(inst2_n2713), .A(inst2_n2693), .ZN(inst2_n2694) );
  OAI22_X1 inst2_U1040 ( .A1(inst2_n1205), .A2(inst2_n2711), .B1(inst2_n2757),
        .B2(inst2_n2831), .ZN(inst2_n2693) );
  OAI21_X1 inst2_U1039 ( .B1(inst2_n1196), .B2(inst2_n2771), .A(inst2_n2692),
        .ZN(inst2_stateArray_S32reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst2_U1038 ( .B1(plaintext2[13]), .B2(inst2_n2713), .A(inst2_n2691), .ZN(inst2_n2692) );
  OAI22_X1 inst2_U1037 ( .A1(inst2_n1204), .A2(inst2_n2711), .B1(inst2_n2760),
        .B2(inst2_n2830), .ZN(inst2_n2691) );
  OAI21_X1 inst2_U1036 ( .B1(inst2_n1195), .B2(inst2_n2771), .A(inst2_n2690),
        .ZN(inst2_stateArray_S32reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst2_U1035 ( .B1(plaintext2[14]), .B2(inst2_n2713), .A(inst2_n2689), .ZN(inst2_n2690) );
  OAI22_X1 inst2_U1034 ( .A1(inst2_n1203), .A2(inst2_n2711), .B1(inst2_n2757),
        .B2(inst2_n2827), .ZN(inst2_n2689) );
  OAI21_X1 inst2_U1033 ( .B1(inst2_n1194), .B2(inst2_n2771), .A(inst2_n2688),
        .ZN(inst2_stateArray_S32reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst2_U1032 ( .B1(plaintext2[15]), .B2(inst2_n2713), .A(inst2_n2687), .ZN(inst2_n2688) );
  OAI22_X1 inst2_U1031 ( .A1(inst2_n1202), .A2(inst2_n2711), .B1(inst2_n2757),
        .B2(inst2_n2829), .ZN(inst2_n2687) );
  OAI211_X1 inst2_U1030 ( .C1(inst2_n706), .C2(inst2_n2791), .A(inst2_n6), .B(
        inst2_n2685), .ZN(inst2_calcRCon_n48) );
  OAI221_X1 inst2_U1029 ( .B1(inst2_n581), .B2(inst2_n1071), .C1(inst2_n2836),
        .C2(inst2_n2801), .A(inst2_n2791), .ZN(inst2_n2685) );
  OAI21_X1 inst2_U1028 ( .B1(inst2_n1225), .B2(inst2_n2771), .A(inst2_n2684),
        .ZN(inst2_stateArray_S22reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst2_U1027 ( .B1(plaintext2[40]), .B2(inst2_n2713), .A(inst2_n2683), .ZN(inst2_n2684) );
  OAI22_X1 inst2_U1026 ( .A1(inst2_n1233), .A2(inst2_n2711), .B1(inst2_n2757),
        .B2(inst2_n2808), .ZN(inst2_n2683) );
  OAI211_X1 inst2_U1025 ( .C1(inst2_n1204), .C2(inst2_n2771), .A(inst2_n2682),
        .B(inst2_n2681), .ZN(inst2_stateArray_S31reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst2_U1024 ( .A1(plaintext2[21]), .A2(inst2_n2713), .ZN(
        inst2_n2681) );
  AOI22_X1 inst2_U1023 ( .A1(inst2_n2788), .A2(ciphertext2[21]), .B1(
        inst2_n2791), .B2(ciphertext2[29]), .ZN(inst2_n2682) );
  OAI21_X1 inst2_U1022 ( .B1(inst2_n1224), .B2(inst2_n2771), .A(inst2_n2680),
        .ZN(inst2_stateArray_S22reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst2_U1021 ( .B1(plaintext2[41]), .B2(inst2_n2713), .A(inst2_n2679), .ZN(inst2_n2680) );
  OAI22_X1 inst2_U1020 ( .A1(inst2_n1232), .A2(inst2_n2711), .B1(inst2_n2760),
        .B2(inst2_n2810), .ZN(inst2_n2679) );
  OAI21_X1 inst2_U1019 ( .B1(inst2_n1223), .B2(inst2_n2771), .A(inst2_n2678),
        .ZN(inst2_stateArray_S22reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst2_U1018 ( .B1(plaintext2[42]), .B2(inst2_n2713), .A(inst2_n2677), .ZN(inst2_n2678) );
  OAI22_X1 inst2_U1017 ( .A1(inst2_n193), .A2(inst2_n2760), .B1(inst2_n1231),
        .B2(inst2_n2711), .ZN(inst2_n2677) );
  INV_X2 inst2_U1016 ( .A(inst2_n6), .ZN(inst2_n2713) );
  OAI21_X1 inst2_U1015 ( .B1(inst2_n1222), .B2(inst2_n2771), .A(inst2_n2676),
        .ZN(inst2_stateArray_S22reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst2_U1014 ( .B1(plaintext2[43]), .B2(inst2_n2550), .A(inst2_n2675), .ZN(inst2_n2676) );
  OAI22_X1 inst2_U1013 ( .A1(inst2_n196), .A2(inst2_n2760), .B1(inst2_n1230),
        .B2(inst2_n2711), .ZN(inst2_n2675) );
  OAI21_X1 inst2_U1012 ( .B1(inst2_n1219), .B2(inst2_n2771), .A(inst2_n2674),
        .ZN(inst2_stateArray_S22reg_gff_1_SFF_6_n6) );
  AOI21_X1 inst2_U1011 ( .B1(plaintext2[46]), .B2(inst2_n2595), .A(inst2_n2673), .ZN(inst2_n2674) );
  OAI22_X1 inst2_U1010 ( .A1(inst2_n1227), .A2(inst2_n2711), .B1(inst2_n2757),
        .B2(inst2_n2807), .ZN(inst2_n2673) );
  OAI21_X1 inst2_U1009 ( .B1(inst2_n1218), .B2(inst2_n2771), .A(inst2_n2672),
        .ZN(inst2_stateArray_S22reg_gff_1_SFF_7_n6) );
  AOI21_X1 inst2_U1008 ( .B1(plaintext2[47]), .B2(inst2_n2722), .A(inst2_n2671), .ZN(inst2_n2672) );
  OAI22_X1 inst2_U1007 ( .A1(inst2_n219), .A2(inst2_n2760), .B1(inst2_n1226),
        .B2(inst2_n2711), .ZN(inst2_n2671) );
  OAI211_X1 inst2_U1006 ( .C1(inst2_n1184), .C2(inst2_n2670), .A(inst2_n2669),
        .B(inst2_n2668), .ZN(inst2_KeyArray_S01reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst2_U1005 ( .A1(inst2_n2667), .A2(inst2_n137), .ZN(inst2_n2668)
         );
  AOI22_X1 inst2_U1004 ( .A1(inst2_n2666), .A2(inst2_n2839), .B1(key2[113]),
        .B2(inst2_n2803), .ZN(inst2_n2669) );
  OAI211_X1 inst2_U1003 ( .C1(inst2_n1183), .C2(inst2_n2670), .A(inst2_n2665),
        .B(inst2_n2664), .ZN(inst2_KeyArray_S01reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst2_U1002 ( .A1(inst2_n2667), .A2(inst2_n136), .ZN(inst2_n2664)
         );
  AOI22_X1 inst2_U1001 ( .A1(inst2_n2666), .A2(inst2_n2825), .B1(key2[114]),
        .B2(inst2_n2803), .ZN(inst2_n2665) );
  OAI211_X1 inst2_U1000 ( .C1(inst2_n1182), .C2(inst2_n2670), .A(inst2_n2663),
        .B(inst2_n2662), .ZN(inst2_KeyArray_S01reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst2_U999 ( .A1(inst2_n2667), .A2(inst2_n135), .ZN(inst2_n2662) );
  AOI22_X1 inst2_U998 ( .A1(inst2_n2666), .A2(inst2_n2824), .B1(key2[115]),
        .B2(inst2_n2803), .ZN(inst2_n2663) );
  OAI211_X1 inst2_U997 ( .C1(inst2_n1181), .C2(inst2_n2670), .A(inst2_n2661),
        .B(inst2_n2660), .ZN(inst2_KeyArray_S01reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst2_U996 ( .A1(inst2_n2667), .A2(inst2_n134), .ZN(inst2_n2660) );
  AOI22_X1 inst2_U995 ( .A1(inst2_n2666), .A2(inst2_n2838), .B1(key2[116]),
        .B2(inst2_n2803), .ZN(inst2_n2661) );
  OAI211_X1 inst2_U994 ( .C1(inst2_n1180), .C2(inst2_n2670), .A(inst2_n2659),
        .B(inst2_n2658), .ZN(inst2_KeyArray_S01reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst2_U993 ( .A1(inst2_n2667), .A2(inst2_n133), .ZN(inst2_n2658) );
  AOI22_X1 inst2_U992 ( .A1(inst2_n2666), .A2(inst2_n2823), .B1(key2[117]),
        .B2(inst2_n2657), .ZN(inst2_n2659) );
  OAI211_X1 inst2_U991 ( .C1(inst2_n1179), .C2(inst2_n2670), .A(inst2_n2656),
        .B(inst2_n2655), .ZN(inst2_KeyArray_S01reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst2_U990 ( .A1(inst2_n2667), .A2(inst2_n132), .ZN(inst2_n2655) );
  AOI22_X1 inst2_U989 ( .A1(inst2_n2666), .A2(inst2_n2822), .B1(key2[118]),
        .B2(inst2_n2657), .ZN(inst2_n2656) );
  OAI211_X1 inst2_U988 ( .C1(inst2_n1178), .C2(inst2_n2670), .A(inst2_n2654),
        .B(inst2_n2653), .ZN(inst2_KeyArray_S01reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst2_U987 ( .A1(inst2_n2667), .A2(inst2_n131), .ZN(inst2_n2653) );
  AOI22_X1 inst2_U986 ( .A1(inst2_n2666), .A2(inst2_n2821), .B1(key2[119]),
        .B2(inst2_n2657), .ZN(inst2_n2654) );
  OAI21_X1 inst2_U985 ( .B1(inst2_n2652), .B2(inst2_n2871), .A(inst2_n2651),
        .ZN(inst2_KeyArray_S02reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst2_U984 ( .B1(key2[104]), .B2(inst2_n2722), .A(inst2_n2650),
        .ZN(inst2_n2651) );
  OAI22_X1 inst2_U983 ( .A1(inst2_n1177), .A2(inst2_n2776), .B1(inst2_n1185),
        .B2(inst2_n2796), .ZN(inst2_n2650) );
  OAI21_X1 inst2_U982 ( .B1(inst2_n2115), .B2(inst2_n2870), .A(inst2_n2649),
        .ZN(inst2_KeyArray_S02reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst2_U981 ( .B1(key2[105]), .B2(inst2_n2484), .A(inst2_n2648),
        .ZN(inst2_n2649) );
  OAI22_X1 inst2_U980 ( .A1(inst2_n1176), .A2(inst2_n2776), .B1(inst2_n1184),
        .B2(inst2_n2647), .ZN(inst2_n2648) );
  OAI21_X1 inst2_U979 ( .B1(inst2_n2652), .B2(inst2_n2869), .A(inst2_n2646),
        .ZN(inst2_KeyArray_S02reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst2_U978 ( .B1(key2[106]), .B2(inst2_n2595), .A(inst2_n2645),
        .ZN(inst2_n2646) );
  OAI22_X1 inst2_U977 ( .A1(inst2_n1175), .A2(inst2_n2776), .B1(inst2_n1183),
        .B2(inst2_n2796), .ZN(inst2_n2645) );
  OAI21_X1 inst2_U976 ( .B1(inst2_n2652), .B2(inst2_n2868), .A(inst2_n2644),
        .ZN(inst2_KeyArray_S02reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst2_U975 ( .B1(key2[107]), .B2(inst2_n2722), .A(inst2_n2643),
        .ZN(inst2_n2644) );
  OAI22_X1 inst2_U974 ( .A1(inst2_n1174), .A2(inst2_n2776), .B1(inst2_n1182),
        .B2(inst2_n2647), .ZN(inst2_n2643) );
  OAI21_X1 inst2_U973 ( .B1(inst2_n2652), .B2(inst2_n2867), .A(inst2_n2642),
        .ZN(inst2_KeyArray_S02reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst2_U972 ( .B1(key2[108]), .B2(inst2_n2657), .A(inst2_n2641),
        .ZN(inst2_n2642) );
  OAI22_X1 inst2_U971 ( .A1(inst2_n1173), .A2(inst2_n2776), .B1(inst2_n1181),
        .B2(inst2_n2796), .ZN(inst2_n2641) );
  OAI21_X1 inst2_U970 ( .B1(inst2_n2652), .B2(inst2_n2866), .A(inst2_n2640),
        .ZN(inst2_KeyArray_S02reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst2_U969 ( .B1(key2[109]), .B2(inst2_n2657), .A(inst2_n2639),
        .ZN(inst2_n2640) );
  OAI22_X1 inst2_U968 ( .A1(inst2_n1172), .A2(inst2_n2776), .B1(inst2_n1180),
        .B2(inst2_n2647), .ZN(inst2_n2639) );
  OAI21_X1 inst2_U967 ( .B1(inst2_n2652), .B2(inst2_n2865), .A(inst2_n2638),
        .ZN(inst2_KeyArray_S02reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst2_U966 ( .B1(key2[110]), .B2(inst2_n2582), .A(inst2_n2637),
        .ZN(inst2_n2638) );
  OAI22_X1 inst2_U965 ( .A1(inst2_n1171), .A2(inst2_n2776), .B1(inst2_n1179),
        .B2(inst2_n2647), .ZN(inst2_n2637) );
  OAI21_X1 inst2_U964 ( .B1(inst2_n2115), .B2(inst2_n2864), .A(inst2_n2636),
        .ZN(inst2_KeyArray_S02reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst2_U963 ( .B1(key2[111]), .B2(inst2_n2713), .A(inst2_n2635),
        .ZN(inst2_n2636) );
  OAI22_X1 inst2_U962 ( .A1(inst2_n1170), .A2(inst2_n2776), .B1(inst2_n1178),
        .B2(inst2_n2647), .ZN(inst2_n2635) );
  OAI21_X1 inst2_U961 ( .B1(inst2_n2652), .B2(inst2_n2847), .A(inst2_n2634),
        .ZN(inst2_KeyArray_S03reg_gff_1_SFF_0_n5) );
  AOI21_X1 inst2_U960 ( .B1(key2[96]), .B2(inst2_n2657), .A(inst2_n2633), .ZN(
        inst2_n2634) );
  OAI22_X1 inst2_U959 ( .A1(inst2_n1169), .A2(inst2_n2776), .B1(inst2_n1177),
        .B2(inst2_n2796), .ZN(inst2_n2633) );
  OAI21_X1 inst2_U958 ( .B1(inst2_n2652), .B2(inst2_n2846), .A(inst2_n2632),
        .ZN(inst2_KeyArray_S03reg_gff_1_SFF_1_n5) );
  AOI21_X1 inst2_U957 ( .B1(key2[97]), .B2(inst2_n2484), .A(inst2_n2631), .ZN(
        inst2_n2632) );
  OAI22_X1 inst2_U956 ( .A1(inst2_n1168), .A2(inst2_n2670), .B1(inst2_n1176),
        .B2(inst2_n2796), .ZN(inst2_n2631) );
  OAI21_X1 inst2_U955 ( .B1(inst2_n2115), .B2(inst2_n2845), .A(inst2_n2630),
        .ZN(inst2_KeyArray_S03reg_gff_1_SFF_2_n5) );
  AOI21_X1 inst2_U954 ( .B1(key2[98]), .B2(inst2_n2713), .A(inst2_n2629), .ZN(
        inst2_n2630) );
  OAI22_X1 inst2_U953 ( .A1(inst2_n1167), .A2(inst2_n2776), .B1(inst2_n1175),
        .B2(inst2_n2796), .ZN(inst2_n2629) );
  OAI21_X1 inst2_U952 ( .B1(inst2_n2652), .B2(inst2_n2844), .A(inst2_n2628),
        .ZN(inst2_KeyArray_S03reg_gff_1_SFF_3_n5) );
  AOI21_X1 inst2_U951 ( .B1(key2[99]), .B2(inst2_n2713), .A(inst2_n2627), .ZN(
        inst2_n2628) );
  OAI22_X1 inst2_U950 ( .A1(inst2_n1166), .A2(inst2_n2463), .B1(inst2_n1174),
        .B2(inst2_n2796), .ZN(inst2_n2627) );
  OAI21_X1 inst2_U949 ( .B1(inst2_n2652), .B2(inst2_n2843), .A(inst2_n2626),
        .ZN(inst2_KeyArray_S03reg_gff_1_SFF_4_n5) );
  AOI21_X1 inst2_U948 ( .B1(key2[100]), .B2(inst2_n2713), .A(inst2_n2625),
        .ZN(inst2_n2626) );
  OAI22_X1 inst2_U947 ( .A1(inst2_n1165), .A2(inst2_n2463), .B1(inst2_n1173),
        .B2(inst2_n2796), .ZN(inst2_n2625) );
  OAI21_X1 inst2_U946 ( .B1(inst2_n2652), .B2(inst2_n2842), .A(inst2_n2624),
        .ZN(inst2_KeyArray_S03reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst2_U945 ( .B1(key2[101]), .B2(inst2_n2713), .A(inst2_n2623),
        .ZN(inst2_n2624) );
  OAI22_X1 inst2_U944 ( .A1(inst2_n1164), .A2(inst2_n2463), .B1(inst2_n1172),
        .B2(inst2_n2796), .ZN(inst2_n2623) );
  OAI21_X1 inst2_U943 ( .B1(inst2_n2652), .B2(inst2_n2841), .A(inst2_n2622),
        .ZN(inst2_KeyArray_S03reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst2_U942 ( .B1(key2[102]), .B2(inst2_n2713), .A(inst2_n2621),
        .ZN(inst2_n2622) );
  OAI22_X1 inst2_U941 ( .A1(inst2_n1163), .A2(inst2_n2463), .B1(inst2_n1171),
        .B2(inst2_n2647), .ZN(inst2_n2621) );
  OAI21_X1 inst2_U940 ( .B1(inst2_n2652), .B2(inst2_n2840), .A(inst2_n2620),
        .ZN(inst2_KeyArray_S03reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst2_U939 ( .B1(key2[103]), .B2(inst2_n2713), .A(inst2_n2619),
        .ZN(inst2_n2620) );
  OAI22_X1 inst2_U938 ( .A1(inst2_n1162), .A2(inst2_n2670), .B1(inst2_n1170),
        .B2(inst2_n2647), .ZN(inst2_n2619) );
  OAI21_X1 inst2_U937 ( .B1(inst2_n2652), .B2(inst2_n2863), .A(inst2_n2618),
        .ZN(inst2_KeyArray_S10reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst2_U936 ( .B1(key2[88]), .B2(inst2_n2713), .A(inst2_n2617), .ZN(
        inst2_n2618) );
  OAI22_X1 inst2_U935 ( .A1(inst2_n1169), .A2(inst2_n2647), .B1(inst2_n1161),
        .B2(inst2_n2776), .ZN(inst2_n2617) );
  OAI211_X1 inst2_U934 ( .C1(inst2_n1168), .C2(inst2_n2796), .A(inst2_n2616),
        .B(inst2_n2615), .ZN(inst2_KeyArray_S10reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst2_U933 ( .A1(inst2_n2667), .A2(inst2_n121), .ZN(inst2_n2615) );
  AOI22_X1 inst2_U932 ( .A1(inst2_n137), .A2(inst2_n2614), .B1(key2[89]), .B2(
        inst2_n2657), .ZN(inst2_n2616) );
  OAI211_X1 inst2_U931 ( .C1(inst2_n1167), .C2(inst2_n2565), .A(inst2_n2613),
        .B(inst2_n2612), .ZN(inst2_KeyArray_S10reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst2_U930 ( .A1(inst2_n2667), .A2(inst2_n120), .ZN(inst2_n2612) );
  AOI22_X1 inst2_U929 ( .A1(inst2_n136), .A2(inst2_n2568), .B1(key2[90]), .B2(
        inst2_n2657), .ZN(inst2_n2613) );
  OAI211_X1 inst2_U928 ( .C1(inst2_n1166), .C2(inst2_n2565), .A(inst2_n2611),
        .B(inst2_n2610), .ZN(inst2_KeyArray_S10reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst2_U927 ( .A1(inst2_n2667), .A2(inst2_n119), .ZN(inst2_n2610) );
  AOI22_X1 inst2_U926 ( .A1(inst2_n135), .A2(inst2_n2568), .B1(key2[91]), .B2(
        inst2_n2657), .ZN(inst2_n2611) );
  OAI211_X1 inst2_U925 ( .C1(inst2_n1165), .C2(inst2_n2796), .A(inst2_n2609),
        .B(inst2_n2608), .ZN(inst2_KeyArray_S10reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst2_U924 ( .A1(inst2_n2667), .A2(inst2_n118), .ZN(inst2_n2608) );
  AOI22_X1 inst2_U923 ( .A1(inst2_n134), .A2(inst2_n2122), .B1(key2[92]), .B2(
        inst2_n2657), .ZN(inst2_n2609) );
  OAI211_X1 inst2_U922 ( .C1(inst2_n1164), .C2(inst2_n2565), .A(inst2_n2607),
        .B(inst2_n2606), .ZN(inst2_KeyArray_S10reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst2_U921 ( .A1(inst2_n2667), .A2(inst2_n117), .ZN(inst2_n2606) );
  AOI22_X1 inst2_U920 ( .A1(inst2_n133), .A2(inst2_n2375), .B1(key2[93]), .B2(
        inst2_n2657), .ZN(inst2_n2607) );
  OAI211_X1 inst2_U919 ( .C1(inst2_n1163), .C2(inst2_n2565), .A(inst2_n2605),
        .B(inst2_n2604), .ZN(inst2_KeyArray_S10reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst2_U918 ( .A1(inst2_n2667), .A2(inst2_n116), .ZN(inst2_n2604) );
  AOI22_X1 inst2_U917 ( .A1(inst2_n132), .A2(inst2_n2568), .B1(key2[94]), .B2(
        inst2_n2657), .ZN(inst2_n2605) );
  OAI211_X1 inst2_U916 ( .C1(inst2_n1162), .C2(inst2_n2565), .A(inst2_n2603),
        .B(inst2_n2602), .ZN(inst2_KeyArray_S10reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst2_U915 ( .A1(inst2_n2667), .A2(inst2_n115), .ZN(inst2_n2602) );
  AOI22_X1 inst2_U914 ( .A1(inst2_n131), .A2(inst2_n2122), .B1(key2[95]), .B2(
        inst2_n2657), .ZN(inst2_n2603) );
  OAI211_X1 inst2_U913 ( .C1(inst2_n1161), .C2(inst2_n2565), .A(inst2_n2601),
        .B(inst2_n2600), .ZN(inst2_KeyArray_S11reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst2_U912 ( .A1(inst2_n2667), .A2(inst2_n114), .ZN(inst2_n2600) );
  AOI22_X1 inst2_U911 ( .A1(inst2_n130), .A2(inst2_n2568), .B1(key2[80]), .B2(
        inst2_n2657), .ZN(inst2_n2601) );
  NAND2_X1 inst2_U910 ( .A1(inst2_n2599), .A2(inst2_n2598), .ZN(
        inst2_KeyArray_S11reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U909 ( .A1(inst2_n2666), .A2(inst2_n137), .B1(inst2_n2667),
        .B2(inst2_n113), .ZN(inst2_n2598) );
  AOI22_X1 inst2_U908 ( .A1(inst2_n129), .A2(inst2_n2568), .B1(key2[81]), .B2(
        inst2_n2657), .ZN(inst2_n2599) );
  INV_X1 inst2_U907 ( .A(inst2_n6), .ZN(inst2_n2657) );
  NAND2_X1 inst2_U906 ( .A1(inst2_n2597), .A2(inst2_n2596), .ZN(
        inst2_KeyArray_S11reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U905 ( .A1(inst2_n2666), .A2(inst2_n136), .B1(inst2_n2667),
        .B2(inst2_n112), .ZN(inst2_n2596) );
  AOI22_X1 inst2_U904 ( .A1(inst2_n128), .A2(inst2_n2614), .B1(key2[82]), .B2(
        inst2_n2595), .ZN(inst2_n2597) );
  NAND2_X1 inst2_U903 ( .A1(inst2_n2594), .A2(inst2_n2593), .ZN(
        inst2_KeyArray_S11reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U902 ( .A1(inst2_n2666), .A2(inst2_n135), .B1(inst2_n2667),
        .B2(inst2_n111), .ZN(inst2_n2593) );
  AOI22_X1 inst2_U901 ( .A1(inst2_n127), .A2(inst2_n2122), .B1(key2[83]), .B2(
        inst2_n2595), .ZN(inst2_n2594) );
  NAND2_X1 inst2_U900 ( .A1(inst2_n2592), .A2(inst2_n2591), .ZN(
        inst2_KeyArray_S11reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U899 ( .A1(inst2_n2666), .A2(inst2_n134), .B1(inst2_n2667),
        .B2(inst2_n110), .ZN(inst2_n2591) );
  AOI22_X1 inst2_U898 ( .A1(inst2_n126), .A2(inst2_n2375), .B1(key2[84]), .B2(
        inst2_n2595), .ZN(inst2_n2592) );
  NAND2_X1 inst2_U897 ( .A1(inst2_n2590), .A2(inst2_n2589), .ZN(
        inst2_KeyArray_S11reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst2_U896 ( .A1(inst2_n2666), .A2(inst2_n133), .B1(inst2_n2667),
        .B2(inst2_n109), .ZN(inst2_n2589) );
  INV_X1 inst2_U895 ( .A(inst2_n2647), .ZN(inst2_n2666) );
  AOI22_X1 inst2_U894 ( .A1(inst2_n125), .A2(inst2_n2614), .B1(key2[85]), .B2(
        inst2_n2595), .ZN(inst2_n2590) );
  NAND2_X1 inst2_U893 ( .A1(inst2_n2588), .A2(inst2_n2587), .ZN(
        inst2_KeyArray_S11reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst2_U892 ( .A1(inst2_n2586), .A2(inst2_n132), .B1(inst2_n2667),
        .B2(inst2_n108), .ZN(inst2_n2587) );
  AOI22_X1 inst2_U891 ( .A1(inst2_n124), .A2(inst2_n2375), .B1(key2[86]), .B2(
        inst2_n2595), .ZN(inst2_n2588) );
  NAND2_X1 inst2_U890 ( .A1(inst2_n2585), .A2(inst2_n2584), .ZN(
        inst2_KeyArray_S11reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst2_U889 ( .A1(inst2_n2586), .A2(inst2_n131), .B1(inst2_n2667),
        .B2(inst2_n107), .ZN(inst2_n2584) );
  AOI22_X1 inst2_U888 ( .A1(inst2_n123), .A2(inst2_n2122), .B1(key2[87]), .B2(
        inst2_n2595), .ZN(inst2_n2585) );
  OAI21_X1 inst2_U887 ( .B1(inst2_n1185), .B2(inst2_n2115), .A(inst2_n2583),
        .ZN(inst2_KeyArray_S32reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst2_U886 ( .B1(key2[8]), .B2(inst2_n2582), .A(inst2_n2581), .ZN(
        inst2_n2583) );
  OAI22_X1 inst2_U885 ( .A1(inst2_n1089), .A2(inst2_n2776), .B1(inst2_n1097),
        .B2(inst2_n2647), .ZN(inst2_n2581) );
  OAI21_X1 inst2_U884 ( .B1(inst2_n1183), .B2(inst2_n2652), .A(inst2_n2580),
        .ZN(inst2_KeyArray_S32reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst2_U883 ( .B1(key2[10]), .B2(inst2_n2582), .A(inst2_n2579), .ZN(
        inst2_n2580) );
  OAI22_X1 inst2_U882 ( .A1(inst2_n1087), .A2(inst2_n2670), .B1(inst2_n1095),
        .B2(inst2_n2796), .ZN(inst2_n2579) );
  OAI21_X1 inst2_U881 ( .B1(inst2_n1182), .B2(inst2_n2115), .A(inst2_n2578),
        .ZN(inst2_KeyArray_S32reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst2_U880 ( .B1(key2[11]), .B2(inst2_n2582), .A(inst2_n2577), .ZN(
        inst2_n2578) );
  OAI22_X1 inst2_U879 ( .A1(inst2_n1086), .A2(inst2_n2776), .B1(inst2_n1094),
        .B2(inst2_n2796), .ZN(inst2_n2577) );
  OAI21_X1 inst2_U878 ( .B1(inst2_n1181), .B2(inst2_n2652), .A(inst2_n2576),
        .ZN(inst2_KeyArray_S32reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst2_U877 ( .B1(key2[12]), .B2(inst2_n2582), .A(inst2_n2575), .ZN(
        inst2_n2576) );
  OAI22_X1 inst2_U876 ( .A1(inst2_n1085), .A2(inst2_n2463), .B1(inst2_n1093),
        .B2(inst2_n2796), .ZN(inst2_n2575) );
  OAI21_X1 inst2_U875 ( .B1(inst2_n1180), .B2(inst2_n2115), .A(inst2_n2574),
        .ZN(inst2_KeyArray_S32reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst2_U874 ( .B1(key2[13]), .B2(inst2_n2582), .A(inst2_n2573), .ZN(
        inst2_n2574) );
  OAI22_X1 inst2_U873 ( .A1(inst2_n1084), .A2(inst2_n2776), .B1(inst2_n1092),
        .B2(inst2_n2647), .ZN(inst2_n2573) );
  OAI21_X1 inst2_U872 ( .B1(inst2_n1179), .B2(inst2_n2652), .A(inst2_n2572),
        .ZN(inst2_KeyArray_S32reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst2_U871 ( .B1(key2[14]), .B2(inst2_n2582), .A(inst2_n2571), .ZN(
        inst2_n2572) );
  OAI22_X1 inst2_U870 ( .A1(inst2_n1083), .A2(inst2_n2670), .B1(inst2_n1091),
        .B2(inst2_n2647), .ZN(inst2_n2571) );
  OAI21_X1 inst2_U869 ( .B1(inst2_n1178), .B2(inst2_n2115), .A(inst2_n2570),
        .ZN(inst2_KeyArray_S32reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst2_U868 ( .B1(key2[15]), .B2(inst2_n2582), .A(inst2_n2569), .ZN(
        inst2_n2570) );
  OAI22_X1 inst2_U867 ( .A1(inst2_n1082), .A2(inst2_n2776), .B1(inst2_n1090),
        .B2(inst2_n2647), .ZN(inst2_n2569) );
  INV_X1 inst2_U866 ( .A(inst2_n2670), .ZN(inst2_n2568) );
  OAI21_X1 inst2_U865 ( .B1(inst2_n1161), .B2(inst2_n2652), .A(inst2_n2567),
        .ZN(inst2_KeyArray_S01reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst2_U864 ( .B1(key2[112]), .B2(inst2_n2722), .A(inst2_n2566),
        .ZN(inst2_n2567) );
  OAI22_X1 inst2_U863 ( .A1(inst2_n1193), .A2(inst2_n2565), .B1(inst2_n1185),
        .B2(inst2_n2776), .ZN(inst2_n2566) );
  NAND2_X1 inst2_U862 ( .A1(inst2_n2564), .A2(inst2_n2563), .ZN(
        inst2_KeyArray_S12reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst2_U861 ( .A1(inst2_n2586), .A2(inst2_n130), .B1(inst2_n2667),
        .B2(inst2_n98), .ZN(inst2_n2563) );
  AOI22_X1 inst2_U860 ( .A1(inst2_n22), .A2(inst2_n2614), .B1(key2[72]), .B2(
        inst2_n2595), .ZN(inst2_n2564) );
  NAND2_X1 inst2_U859 ( .A1(inst2_n2562), .A2(inst2_n2561), .ZN(
        inst2_KeyArray_S12reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U858 ( .A1(inst2_n2586), .A2(inst2_n129), .B1(inst2_n2667),
        .B2(inst2_n97), .ZN(inst2_n2561) );
  AOI22_X1 inst2_U857 ( .A1(inst2_n17), .A2(inst2_n2122), .B1(key2[73]), .B2(
        inst2_n2595), .ZN(inst2_n2562) );
  NAND2_X1 inst2_U856 ( .A1(inst2_n2560), .A2(inst2_n2559), .ZN(
        inst2_KeyArray_S12reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U855 ( .A1(inst2_n2586), .A2(inst2_n128), .B1(inst2_n2667),
        .B2(inst2_n96), .ZN(inst2_n2559) );
  AOI22_X1 inst2_U854 ( .A1(inst2_n14), .A2(inst2_n2568), .B1(key2[74]), .B2(
        inst2_n2595), .ZN(inst2_n2560) );
  NAND2_X1 inst2_U853 ( .A1(inst2_n2558), .A2(inst2_n2557), .ZN(
        inst2_KeyArray_S12reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U852 ( .A1(inst2_n2586), .A2(inst2_n127), .B1(inst2_n2667),
        .B2(inst2_n95), .ZN(inst2_n2557) );
  AOI22_X1 inst2_U851 ( .A1(inst2_n12), .A2(inst2_n2614), .B1(key2[75]), .B2(
        inst2_n2595), .ZN(inst2_n2558) );
  NAND2_X1 inst2_U850 ( .A1(inst2_n2556), .A2(inst2_n2555), .ZN(
        inst2_KeyArray_S12reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U849 ( .A1(inst2_n2586), .A2(inst2_n126), .B1(inst2_n2667),
        .B2(inst2_n94), .ZN(inst2_n2555) );
  AOI22_X1 inst2_U848 ( .A1(inst2_n11), .A2(inst2_n2568), .B1(key2[76]), .B2(
        inst2_n2595), .ZN(inst2_n2556) );
  NAND2_X1 inst2_U847 ( .A1(inst2_n2554), .A2(inst2_n2553), .ZN(
        inst2_KeyArray_S12reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst2_U846 ( .A1(inst2_n2586), .A2(inst2_n125), .B1(inst2_n2667),
        .B2(inst2_n93), .ZN(inst2_n2553) );
  AOI22_X1 inst2_U845 ( .A1(inst2_n10), .A2(inst2_n2122), .B1(key2[77]), .B2(
        inst2_n2595), .ZN(inst2_n2554) );
  INV_X1 inst2_U844 ( .A(inst2_n6), .ZN(inst2_n2595) );
  NAND2_X1 inst2_U843 ( .A1(inst2_n2552), .A2(inst2_n2551), .ZN(
        inst2_KeyArray_S12reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst2_U842 ( .A1(inst2_n2586), .A2(inst2_n124), .B1(inst2_n2667),
        .B2(inst2_n92), .ZN(inst2_n2551) );
  AOI22_X1 inst2_U841 ( .A1(inst2_n24), .A2(inst2_n2122), .B1(key2[78]), .B2(
        inst2_n2550), .ZN(inst2_n2552) );
  NAND2_X1 inst2_U840 ( .A1(inst2_n2549), .A2(inst2_n2548), .ZN(
        inst2_KeyArray_S12reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst2_U839 ( .A1(inst2_n2586), .A2(inst2_n123), .B1(inst2_n2667),
        .B2(inst2_n91), .ZN(inst2_n2548) );
  AOI22_X1 inst2_U838 ( .A1(inst2_n9), .A2(inst2_n2122), .B1(key2[79]), .B2(
        inst2_n2550), .ZN(inst2_n2549) );
  NAND2_X1 inst2_U837 ( .A1(inst2_n2547), .A2(inst2_n2546), .ZN(
        inst2_KeyArray_S13reg_gff_1_SFF_0_n5) );
  AOI22_X1 inst2_U836 ( .A1(inst2_n2586), .A2(inst2_n22), .B1(inst2_n2667),
        .B2(inst2_n90), .ZN(inst2_n2546) );
  AOI22_X1 inst2_U835 ( .A1(inst2_n122), .A2(inst2_n2122), .B1(key2[64]), .B2(
        inst2_n2550), .ZN(inst2_n2547) );
  NAND2_X1 inst2_U834 ( .A1(inst2_n2545), .A2(inst2_n2544), .ZN(
        inst2_KeyArray_S13reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst2_U833 ( .A1(inst2_n2543), .A2(inst2_n17), .B1(inst2_n2667),
        .B2(inst2_n89), .ZN(inst2_n2544) );
  AOI22_X1 inst2_U832 ( .A1(inst2_n121), .A2(inst2_n2122), .B1(key2[65]), .B2(
        inst2_n2550), .ZN(inst2_n2545) );
  NAND2_X1 inst2_U831 ( .A1(inst2_n2542), .A2(inst2_n2541), .ZN(
        inst2_KeyArray_S13reg_gff_1_SFF_2_n5) );
  AOI22_X1 inst2_U830 ( .A1(inst2_n2586), .A2(inst2_n14), .B1(inst2_n2667),
        .B2(inst2_n88), .ZN(inst2_n2541) );
  INV_X1 inst2_U829 ( .A(inst2_n2647), .ZN(inst2_n2586) );
  AOI22_X1 inst2_U828 ( .A1(inst2_n120), .A2(inst2_n2122), .B1(key2[66]), .B2(
        inst2_n2550), .ZN(inst2_n2542) );
  NAND2_X1 inst2_U827 ( .A1(inst2_n2540), .A2(inst2_n2539), .ZN(
        inst2_KeyArray_S13reg_gff_1_SFF_3_n5) );
  AOI22_X1 inst2_U826 ( .A1(inst2_n2586), .A2(inst2_n12), .B1(inst2_n2667),
        .B2(inst2_n87), .ZN(inst2_n2539) );
  AOI22_X1 inst2_U825 ( .A1(inst2_n119), .A2(inst2_n2122), .B1(key2[67]), .B2(
        inst2_n2550), .ZN(inst2_n2540) );
  NAND2_X1 inst2_U824 ( .A1(inst2_n2538), .A2(inst2_n2537), .ZN(
        inst2_KeyArray_S13reg_gff_1_SFF_4_n5) );
  AOI22_X1 inst2_U823 ( .A1(inst2_n2543), .A2(inst2_n11), .B1(inst2_n2667),
        .B2(inst2_n86), .ZN(inst2_n2537) );
  AOI22_X1 inst2_U822 ( .A1(inst2_n118), .A2(inst2_n2122), .B1(key2[68]), .B2(
        inst2_n2550), .ZN(inst2_n2538) );
  NAND2_X1 inst2_U821 ( .A1(inst2_n2536), .A2(inst2_n2535), .ZN(
        inst2_KeyArray_S13reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst2_U820 ( .A1(inst2_n2872), .A2(inst2_n10), .B1(inst2_n2667),
        .B2(inst2_n85), .ZN(inst2_n2535) );
  AOI22_X1 inst2_U819 ( .A1(inst2_n117), .A2(inst2_n2122), .B1(key2[69]), .B2(
        inst2_n2550), .ZN(inst2_n2536) );
  NAND2_X1 inst2_U818 ( .A1(inst2_n2534), .A2(inst2_n2533), .ZN(
        inst2_KeyArray_S13reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst2_U817 ( .A1(inst2_n2586), .A2(inst2_n24), .B1(inst2_n2667),
        .B2(inst2_n84), .ZN(inst2_n2533) );
  AOI22_X1 inst2_U816 ( .A1(inst2_n116), .A2(inst2_n2122), .B1(key2[70]), .B2(
        inst2_n2550), .ZN(inst2_n2534) );
  NAND2_X1 inst2_U815 ( .A1(inst2_n2532), .A2(inst2_n2531), .ZN(
        inst2_KeyArray_S13reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst2_U814 ( .A1(inst2_n2543), .A2(inst2_n9), .B1(inst2_n2667),
        .B2(inst2_n83), .ZN(inst2_n2531) );
  AOI22_X1 inst2_U813 ( .A1(inst2_n115), .A2(inst2_n2614), .B1(key2[71]), .B2(
        inst2_n2550), .ZN(inst2_n2532) );
  NAND2_X1 inst2_U812 ( .A1(inst2_n2530), .A2(inst2_n2529), .ZN(
        inst2_KeyArray_S20reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst2_U811 ( .A1(inst2_n2872), .A2(inst2_n122), .B1(inst2_n2667),
        .B2(inst2_n82), .ZN(inst2_n2529) );
  AOI22_X1 inst2_U810 ( .A1(inst2_n114), .A2(inst2_n2614), .B1(key2[56]), .B2(
        inst2_n2528), .ZN(inst2_n2530) );
  NAND2_X1 inst2_U809 ( .A1(inst2_n2527), .A2(inst2_n2526), .ZN(
        inst2_KeyArray_S20reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U808 ( .A1(inst2_n2586), .A2(inst2_n121), .B1(inst2_n2667),
        .B2(inst2_n81), .ZN(inst2_n2526) );
  AOI22_X1 inst2_U807 ( .A1(inst2_n113), .A2(inst2_n2614), .B1(key2[57]), .B2(
        inst2_n2550), .ZN(inst2_n2527) );
  NAND2_X1 inst2_U806 ( .A1(inst2_n2525), .A2(inst2_n2524), .ZN(
        inst2_KeyArray_S20reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U805 ( .A1(inst2_n2666), .A2(inst2_n120), .B1(inst2_n2667),
        .B2(inst2_n80), .ZN(inst2_n2524) );
  AOI22_X1 inst2_U804 ( .A1(inst2_n112), .A2(inst2_n2614), .B1(key2[58]), .B2(
        inst2_n2528), .ZN(inst2_n2525) );
  NAND2_X1 inst2_U803 ( .A1(inst2_n2523), .A2(inst2_n2522), .ZN(
        inst2_KeyArray_S20reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U802 ( .A1(inst2_n2586), .A2(inst2_n119), .B1(inst2_n2667),
        .B2(inst2_n79), .ZN(inst2_n2522) );
  AOI22_X1 inst2_U801 ( .A1(inst2_n111), .A2(inst2_n2614), .B1(key2[59]), .B2(
        inst2_n2528), .ZN(inst2_n2523) );
  NAND2_X1 inst2_U800 ( .A1(inst2_n2521), .A2(inst2_n2520), .ZN(
        inst2_KeyArray_S20reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U799 ( .A1(inst2_n2586), .A2(inst2_n118), .B1(inst2_n78),
        .B2(inst2_n2667), .ZN(inst2_n2520) );
  AOI22_X1 inst2_U798 ( .A1(inst2_n110), .A2(inst2_n2614), .B1(key2[60]), .B2(
        inst2_n2528), .ZN(inst2_n2521) );
  NAND2_X1 inst2_U797 ( .A1(inst2_n2519), .A2(inst2_n2518), .ZN(
        inst2_KeyArray_S20reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst2_U796 ( .A1(inst2_n2543), .A2(inst2_n117), .B1(inst2_n2667),
        .B2(inst2_n77), .ZN(inst2_n2518) );
  AOI22_X1 inst2_U795 ( .A1(inst2_n109), .A2(inst2_n2614), .B1(key2[61]), .B2(
        inst2_n2528), .ZN(inst2_n2519) );
  NAND2_X1 inst2_U794 ( .A1(inst2_n2517), .A2(inst2_n2516), .ZN(
        inst2_KeyArray_S20reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst2_U793 ( .A1(inst2_n2872), .A2(inst2_n116), .B1(inst2_n2667),
        .B2(inst2_n76), .ZN(inst2_n2516) );
  AOI22_X1 inst2_U792 ( .A1(inst2_n108), .A2(inst2_n2614), .B1(key2[62]), .B2(
        inst2_n2528), .ZN(inst2_n2517) );
  NAND2_X1 inst2_U791 ( .A1(inst2_n2515), .A2(inst2_n2514), .ZN(
        inst2_KeyArray_S20reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst2_U790 ( .A1(inst2_n2543), .A2(inst2_n115), .B1(inst2_n2667),
        .B2(inst2_n75), .ZN(inst2_n2514) );
  AOI22_X1 inst2_U789 ( .A1(inst2_n107), .A2(inst2_n2614), .B1(key2[63]), .B2(
        inst2_n2528), .ZN(inst2_n2515) );
  NAND2_X1 inst2_U788 ( .A1(inst2_n2513), .A2(inst2_n2512), .ZN(
        inst2_KeyArray_S21reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst2_U787 ( .A1(inst2_n2543), .A2(inst2_n114), .B1(inst2_n2667),
        .B2(inst2_n74), .ZN(inst2_n2512) );
  AOI22_X1 inst2_U786 ( .A1(inst2_n98), .A2(inst2_n2614), .B1(key2[48]), .B2(
        inst2_n2528), .ZN(inst2_n2513) );
  NAND2_X1 inst2_U785 ( .A1(inst2_n2511), .A2(inst2_n2510), .ZN(
        inst2_KeyArray_S21reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U784 ( .A1(inst2_n2543), .A2(inst2_n113), .B1(inst2_n2667),
        .B2(inst2_n73), .ZN(inst2_n2510) );
  AOI22_X1 inst2_U783 ( .A1(inst2_n97), .A2(inst2_n2614), .B1(key2[49]), .B2(
        inst2_n2528), .ZN(inst2_n2511) );
  INV_X1 inst2_U782 ( .A(inst2_n2670), .ZN(inst2_n2614) );
  NAND2_X1 inst2_U781 ( .A1(inst2_n2509), .A2(inst2_n2508), .ZN(
        inst2_KeyArray_S21reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U780 ( .A1(inst2_n2543), .A2(inst2_n112), .B1(inst2_n2667),
        .B2(inst2_n72), .ZN(inst2_n2508) );
  AOI22_X1 inst2_U779 ( .A1(inst2_n96), .A2(inst2_n2375), .B1(key2[50]), .B2(
        inst2_n2507), .ZN(inst2_n2509) );
  NAND2_X1 inst2_U778 ( .A1(inst2_n2506), .A2(inst2_n2505), .ZN(
        inst2_KeyArray_S21reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U777 ( .A1(inst2_n2543), .A2(inst2_n111), .B1(inst2_n2667),
        .B2(inst2_n71), .ZN(inst2_n2505) );
  AOI22_X1 inst2_U776 ( .A1(inst2_n95), .A2(inst2_n2568), .B1(key2[51]), .B2(
        inst2_n2528), .ZN(inst2_n2506) );
  NAND2_X1 inst2_U775 ( .A1(inst2_n2504), .A2(inst2_n2503), .ZN(
        inst2_KeyArray_S21reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U774 ( .A1(inst2_n2543), .A2(inst2_n110), .B1(inst2_n70),
        .B2(inst2_n2667), .ZN(inst2_n2503) );
  AOI22_X1 inst2_U773 ( .A1(inst2_n94), .A2(inst2_n2122), .B1(key2[52]), .B2(
        inst2_n2507), .ZN(inst2_n2504) );
  NAND2_X1 inst2_U772 ( .A1(inst2_n2502), .A2(inst2_n2501), .ZN(
        inst2_KeyArray_S21reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst2_U771 ( .A1(inst2_n2543), .A2(inst2_n109), .B1(inst2_n2667),
        .B2(inst2_n69), .ZN(inst2_n2501) );
  AOI22_X1 inst2_U770 ( .A1(inst2_n93), .A2(inst2_n2375), .B1(key2[53]), .B2(
        inst2_n2528), .ZN(inst2_n2502) );
  NAND2_X1 inst2_U769 ( .A1(inst2_n2500), .A2(inst2_n2499), .ZN(
        inst2_KeyArray_S21reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst2_U768 ( .A1(inst2_n2543), .A2(inst2_n108), .B1(inst2_n2667),
        .B2(inst2_n68), .ZN(inst2_n2499) );
  AOI22_X1 inst2_U767 ( .A1(inst2_n92), .A2(inst2_n2568), .B1(key2[54]), .B2(
        inst2_n2507), .ZN(inst2_n2500) );
  NAND2_X1 inst2_U766 ( .A1(inst2_n2498), .A2(inst2_n2497), .ZN(
        inst2_KeyArray_S21reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst2_U765 ( .A1(inst2_n2543), .A2(inst2_n107), .B1(inst2_n2667),
        .B2(inst2_n67), .ZN(inst2_n2497) );
  AOI22_X1 inst2_U764 ( .A1(inst2_n91), .A2(inst2_n2375), .B1(key2[55]), .B2(
        inst2_n2507), .ZN(inst2_n2498) );
  OAI211_X1 inst2_U763 ( .C1(inst2_n1097), .C2(inst2_n2652), .A(inst2_n2496),
        .B(inst2_n2495), .ZN(inst2_KeyArray_S22reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst2_U762 ( .A1(inst2_n2872), .A2(inst2_n98), .ZN(inst2_n2495) );
  AOI22_X1 inst2_U761 ( .A1(inst2_n90), .A2(inst2_n2375), .B1(key2[40]), .B2(
        inst2_n2528), .ZN(inst2_n2496) );
  INV_X1 inst2_U760 ( .A(inst2_n6), .ZN(inst2_n2528) );
  NAND2_X1 inst2_U759 ( .A1(inst2_n2494), .A2(inst2_n2493), .ZN(
        inst2_KeyArray_S22reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U758 ( .A1(inst2_n2543), .A2(inst2_n97), .B1(inst2_n2667),
        .B2(inst2_n65), .ZN(inst2_n2493) );
  AOI22_X1 inst2_U757 ( .A1(inst2_n89), .A2(inst2_n2568), .B1(key2[41]), .B2(
        inst2_n2507), .ZN(inst2_n2494) );
  OAI211_X1 inst2_U756 ( .C1(inst2_n1095), .C2(inst2_n2652), .A(inst2_n2492),
        .B(inst2_n2491), .ZN(inst2_KeyArray_S22reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst2_U755 ( .A1(inst2_n2872), .A2(inst2_n96), .ZN(inst2_n2491) );
  AOI22_X1 inst2_U754 ( .A1(inst2_n88), .A2(inst2_n2568), .B1(key2[42]), .B2(
        inst2_n2507), .ZN(inst2_n2492) );
  OAI211_X1 inst2_U753 ( .C1(inst2_n1094), .C2(inst2_n2652), .A(inst2_n2490),
        .B(inst2_n2489), .ZN(inst2_KeyArray_S22reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst2_U752 ( .A1(inst2_n2098), .A2(inst2_n95), .ZN(inst2_n2489) );
  AOI22_X1 inst2_U751 ( .A1(inst2_n87), .A2(inst2_n2568), .B1(key2[43]), .B2(
        inst2_n2507), .ZN(inst2_n2490) );
  OAI211_X1 inst2_U750 ( .C1(inst2_n1093), .C2(inst2_n2652), .A(inst2_n2488),
        .B(inst2_n2487), .ZN(inst2_KeyArray_S22reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst2_U749 ( .A1(inst2_n2872), .A2(inst2_n94), .ZN(inst2_n2487) );
  AOI22_X1 inst2_U748 ( .A1(inst2_n86), .A2(inst2_n2614), .B1(key2[44]), .B2(
        inst2_n2507), .ZN(inst2_n2488) );
  OAI211_X1 inst2_U747 ( .C1(inst2_n1092), .C2(inst2_n2652), .A(inst2_n2486),
        .B(inst2_n2485), .ZN(inst2_KeyArray_S22reg_gff_1_SFF_5_n5) );
  NAND2_X1 inst2_U746 ( .A1(inst2_n2098), .A2(inst2_n93), .ZN(inst2_n2485) );
  AOI22_X1 inst2_U745 ( .A1(inst2_n85), .A2(inst2_n2614), .B1(key2[45]), .B2(
        inst2_n2484), .ZN(inst2_n2486) );
  OAI211_X1 inst2_U744 ( .C1(inst2_n1091), .C2(inst2_n2652), .A(inst2_n2483),
        .B(inst2_n2482), .ZN(inst2_KeyArray_S22reg_gff_1_SFF_6_n5) );
  NAND2_X1 inst2_U743 ( .A1(inst2_n2098), .A2(inst2_n92), .ZN(inst2_n2482) );
  AOI22_X1 inst2_U742 ( .A1(inst2_n84), .A2(inst2_n2375), .B1(key2[46]), .B2(
        inst2_n2507), .ZN(inst2_n2483) );
  OAI211_X1 inst2_U741 ( .C1(inst2_n1090), .C2(inst2_n2652), .A(inst2_n2481),
        .B(inst2_n2480), .ZN(inst2_KeyArray_S22reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst2_U740 ( .A1(inst2_n2872), .A2(inst2_n91), .ZN(inst2_n2480) );
  AOI22_X1 inst2_U739 ( .A1(inst2_n83), .A2(inst2_n2568), .B1(key2[47]), .B2(
        inst2_n2484), .ZN(inst2_n2481) );
  OAI211_X1 inst2_U738 ( .C1(inst2_n1089), .C2(inst2_n2115), .A(inst2_n2479),
        .B(inst2_n2478), .ZN(inst2_KeyArray_S23reg_gff_1_SFF_0_n5) );
  NAND2_X1 inst2_U737 ( .A1(inst2_n2098), .A2(inst2_n90), .ZN(inst2_n2478) );
  AOI22_X1 inst2_U736 ( .A1(inst2_n82), .A2(inst2_n2375), .B1(key2[32]), .B2(
        inst2_n2507), .ZN(inst2_n2479) );
  NAND2_X1 inst2_U735 ( .A1(inst2_n2477), .A2(inst2_n2476), .ZN(
        inst2_KeyArray_S23reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst2_U734 ( .A1(inst2_n2586), .A2(inst2_n89), .B1(inst2_n2667),
        .B2(inst2_n57), .ZN(inst2_n2476) );
  AOI22_X1 inst2_U733 ( .A1(inst2_n81), .A2(inst2_n2375), .B1(key2[33]), .B2(
        inst2_n2507), .ZN(inst2_n2477) );
  OAI211_X1 inst2_U732 ( .C1(inst2_n1087), .C2(inst2_n2115), .A(inst2_n2475),
        .B(inst2_n2474), .ZN(inst2_KeyArray_S23reg_gff_1_SFF_2_n5) );
  NAND2_X1 inst2_U731 ( .A1(inst2_n2872), .A2(inst2_n88), .ZN(inst2_n2474) );
  AOI22_X1 inst2_U730 ( .A1(inst2_n80), .A2(inst2_n2568), .B1(key2[34]), .B2(
        inst2_n2507), .ZN(inst2_n2475) );
  INV_X1 inst2_U729 ( .A(inst2_n6), .ZN(inst2_n2507) );
  OAI211_X1 inst2_U728 ( .C1(inst2_n1086), .C2(inst2_n2115), .A(inst2_n2473),
        .B(inst2_n2472), .ZN(inst2_KeyArray_S23reg_gff_1_SFF_3_n5) );
  NAND2_X1 inst2_U727 ( .A1(inst2_n2872), .A2(inst2_n87), .ZN(inst2_n2472) );
  AOI22_X1 inst2_U726 ( .A1(inst2_n79), .A2(inst2_n2375), .B1(key2[35]), .B2(
        inst2_n2484), .ZN(inst2_n2473) );
  OAI211_X1 inst2_U725 ( .C1(inst2_n1085), .C2(inst2_n2115), .A(inst2_n2471),
        .B(inst2_n2470), .ZN(inst2_KeyArray_S23reg_gff_1_SFF_4_n5) );
  NAND2_X1 inst2_U724 ( .A1(inst2_n2543), .A2(inst2_n86), .ZN(inst2_n2470) );
  AOI22_X1 inst2_U723 ( .A1(inst2_n2122), .A2(inst2_n78), .B1(key2[36]), .B2(
        inst2_n2484), .ZN(inst2_n2471) );
  OAI211_X1 inst2_U722 ( .C1(inst2_n1084), .C2(inst2_n2115), .A(inst2_n2469),
        .B(inst2_n2468), .ZN(inst2_KeyArray_S23reg_gff_1_SFF_5_n5) );
  NAND2_X1 inst2_U721 ( .A1(inst2_n2543), .A2(inst2_n85), .ZN(inst2_n2468) );
  AOI22_X1 inst2_U720 ( .A1(inst2_n77), .A2(inst2_n2568), .B1(key2[37]), .B2(
        inst2_n2484), .ZN(inst2_n2469) );
  OAI211_X1 inst2_U719 ( .C1(inst2_n1083), .C2(inst2_n2115), .A(inst2_n2467),
        .B(inst2_n2466), .ZN(inst2_KeyArray_S23reg_gff_1_SFF_6_n5) );
  NAND2_X1 inst2_U718 ( .A1(inst2_n2543), .A2(inst2_n84), .ZN(inst2_n2466) );
  AOI22_X1 inst2_U717 ( .A1(inst2_n76), .A2(inst2_n2375), .B1(key2[38]), .B2(
        inst2_n2484), .ZN(inst2_n2467) );
  OAI211_X1 inst2_U716 ( .C1(inst2_n1082), .C2(inst2_n2115), .A(inst2_n2465),
        .B(inst2_n2464), .ZN(inst2_KeyArray_S23reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst2_U715 ( .A1(inst2_n2543), .A2(inst2_n83), .ZN(inst2_n2464) );
  AOI22_X1 inst2_U714 ( .A1(inst2_n75), .A2(inst2_n2568), .B1(key2[39]), .B2(
        inst2_n2484), .ZN(inst2_n2465) );
  OAI211_X1 inst2_U713 ( .C1(inst2_n1097), .C2(inst2_n2463), .A(inst2_n2462),
        .B(inst2_n2461), .ZN(inst2_KeyArray_S31reg_gff_1_SFF_0_n6) );
  OR2_X1 inst2_U712 ( .A1(inst2_n2652), .A2(inst2_n1193), .ZN(inst2_n2461) );
  AOI22_X1 inst2_U711 ( .A1(inst2_n74), .A2(inst2_n2586), .B1(key2[16]), .B2(
        inst2_n2657), .ZN(inst2_n2462) );
  OAI211_X1 inst2_U710 ( .C1(inst2_n1192), .C2(inst2_n2652), .A(inst2_n2460),
        .B(inst2_n2459), .ZN(inst2_KeyArray_S31reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst2_U709 ( .A1(inst2_n2543), .A2(inst2_n73), .ZN(inst2_n2459) );
  AOI22_X1 inst2_U708 ( .A1(inst2_n65), .A2(inst2_n2375), .B1(key2[17]), .B2(
        inst2_n2484), .ZN(inst2_n2460) );
  OAI211_X1 inst2_U707 ( .C1(inst2_n1095), .C2(inst2_n2670), .A(inst2_n2458),
        .B(inst2_n2457), .ZN(inst2_KeyArray_S31reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst2_U706 ( .A1(inst2_n2667), .A2(inst2_n2825), .ZN(inst2_n2457)
         );
  AOI22_X1 inst2_U705 ( .A1(inst2_n72), .A2(inst2_n2543), .B1(key2[18]), .B2(
        inst2_n2713), .ZN(inst2_n2458) );
  OAI211_X1 inst2_U704 ( .C1(inst2_n1094), .C2(inst2_n2670), .A(inst2_n2456),
        .B(inst2_n2455), .ZN(inst2_KeyArray_S31reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst2_U703 ( .A1(inst2_n2667), .A2(inst2_n2824), .ZN(inst2_n2455)
         );
  AOI22_X1 inst2_U702 ( .A1(inst2_n71), .A2(inst2_n2098), .B1(key2[19]), .B2(
        inst2_n2484), .ZN(inst2_n2456) );
  OAI21_X1 inst2_U701 ( .B1(inst2_n1189), .B2(inst2_n2652), .A(inst2_n2454),
        .ZN(inst2_KeyArray_S31reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst2_U700 ( .B1(key2[20]), .B2(inst2_n2722), .A(inst2_n2453), .ZN(
        inst2_n2454) );
  OAI22_X1 inst2_U699 ( .A1(inst2_n1093), .A2(inst2_n2463), .B1(inst2_n2796),
        .B2(inst2_n2828), .ZN(inst2_n2453) );
  OAI211_X1 inst2_U698 ( .C1(inst2_n1092), .C2(inst2_n2670), .A(inst2_n2452),
        .B(inst2_n2451), .ZN(inst2_KeyArray_S31reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst2_U697 ( .A1(inst2_n2667), .A2(inst2_n2823), .ZN(inst2_n2451)
         );
  AOI22_X1 inst2_U696 ( .A1(inst2_n69), .A2(inst2_n2666), .B1(key2[21]), .B2(
        inst2_n2484), .ZN(inst2_n2452) );
  OAI211_X1 inst2_U695 ( .C1(inst2_n1091), .C2(inst2_n2670), .A(inst2_n2450),
        .B(inst2_n2449), .ZN(inst2_KeyArray_S31reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst2_U694 ( .A1(inst2_n2667), .A2(inst2_n2822), .ZN(inst2_n2449)
         );
  AOI22_X1 inst2_U693 ( .A1(inst2_n68), .A2(inst2_n2872), .B1(key2[22]), .B2(
        inst2_n2484), .ZN(inst2_n2450) );
  OAI211_X1 inst2_U692 ( .C1(inst2_n1090), .C2(inst2_n2670), .A(inst2_n2448),
        .B(inst2_n2447), .ZN(inst2_KeyArray_S31reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst2_U691 ( .A1(inst2_n2667), .A2(inst2_n2821), .ZN(inst2_n2447)
         );
  AOI22_X1 inst2_U690 ( .A1(inst2_n67), .A2(inst2_n2586), .B1(key2[23]), .B2(
        inst2_n2528), .ZN(inst2_n2448) );
  OAI211_X1 inst2_U689 ( .C1(inst2_n1184), .C2(inst2_n2652), .A(inst2_n2446),
        .B(inst2_n2445), .ZN(inst2_KeyArray_S32reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst2_U688 ( .A1(inst2_n2543), .A2(inst2_n65), .ZN(inst2_n2445) );
  AOI22_X1 inst2_U687 ( .A1(inst2_n57), .A2(inst2_n2568), .B1(key2[9]), .B2(
        inst2_n2484), .ZN(inst2_n2446) );
  INV_X1 inst2_U686 ( .A(inst2_n6), .ZN(inst2_n2484) );
  OAI21_X1 inst2_U685 ( .B1(inst2_n1265), .B2(inst2_n2444), .A(inst2_n2443),
        .ZN(inst2_stateArray_S10reg_gff_1_SFF_0_n5) );
  AOI22_X1 inst2_U684 ( .A1(inst2_n2788), .A2(ciphertext2[88]), .B1(
        plaintext2[88]), .B2(inst2_n2550), .ZN(inst2_n2443) );
  INV_X1 inst2_U683 ( .A(inst2_n6), .ZN(inst2_n2550) );
  OAI21_X1 inst2_U682 ( .B1(inst2_n1264), .B2(inst2_n2444), .A(inst2_n2442),
        .ZN(inst2_stateArray_S10reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst2_U681 ( .A1(done2), .A2(ciphertext2[89]), .B1(plaintext2[89]),
        .B2(inst2_n2582), .ZN(inst2_n2442) );
  OAI21_X1 inst2_U680 ( .B1(inst2_n1263), .B2(inst2_n2444), .A(inst2_n2441),
        .ZN(inst2_stateArray_S10reg_gff_1_SFF_2_n5) );
  AOI22_X1 inst2_U679 ( .A1(inst2_n2788), .A2(ciphertext2[90]), .B1(
        plaintext2[90]), .B2(inst2_n2722), .ZN(inst2_n2441) );
  OAI21_X1 inst2_U678 ( .B1(inst2_n1262), .B2(inst2_n2444), .A(inst2_n2440),
        .ZN(inst2_stateArray_S10reg_gff_1_SFF_3_n5) );
  AOI22_X1 inst2_U677 ( .A1(done2), .A2(ciphertext2[91]), .B1(plaintext2[91]),
        .B2(inst2_n2484), .ZN(inst2_n2440) );
  OAI21_X1 inst2_U676 ( .B1(inst2_n1261), .B2(inst2_n2444), .A(inst2_n2439),
        .ZN(inst2_stateArray_S10reg_gff_1_SFF_4_n5) );
  AOI22_X1 inst2_U675 ( .A1(inst2_n2788), .A2(ciphertext2[92]), .B1(
        plaintext2[92]), .B2(inst2_n2582), .ZN(inst2_n2439) );
  OAI21_X1 inst2_U674 ( .B1(inst2_n1260), .B2(inst2_n2444), .A(inst2_n2438),
        .ZN(inst2_stateArray_S10reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst2_U673 ( .A1(inst2_n2788), .A2(ciphertext2[93]), .B1(
        plaintext2[93]), .B2(inst2_n2657), .ZN(inst2_n2438) );
  OAI21_X1 inst2_U672 ( .B1(inst2_n1259), .B2(inst2_n2444), .A(inst2_n2437),
        .ZN(inst2_stateArray_S10reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst2_U671 ( .A1(inst2_n2788), .A2(ciphertext2[94]), .B1(
        plaintext2[94]), .B2(inst2_n2722), .ZN(inst2_n2437) );
  OAI21_X1 inst2_U670 ( .B1(inst2_n1258), .B2(inst2_n2444), .A(inst2_n2436),
        .ZN(inst2_stateArray_S10reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst2_U669 ( .A1(inst2_n2788), .A2(ciphertext2[95]), .B1(
        plaintext2[95]), .B2(inst2_n2595), .ZN(inst2_n2436) );
  INV_X1 inst2_U668 ( .A(inst2_n2435), .ZN(inst2_n2444) );
  OAI21_X1 inst2_U667 ( .B1(inst2_n1265), .B2(inst2_n2711), .A(inst2_n2434),
        .ZN(inst2_stateArray_S11reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst2_U666 ( .A1(inst2_n2435), .A2(ciphertext2[72]), .B1(
        plaintext2[80]), .B2(inst2_n2550), .ZN(inst2_n2434) );
  OAI21_X1 inst2_U665 ( .B1(inst2_n1264), .B2(inst2_n2711), .A(inst2_n2433),
        .ZN(inst2_stateArray_S11reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U664 ( .A1(inst2_n2435), .A2(ciphertext2[73]), .B1(
        plaintext2[81]), .B2(inst2_n2550), .ZN(inst2_n2433) );
  OAI21_X1 inst2_U663 ( .B1(inst2_n1263), .B2(inst2_n2711), .A(inst2_n2432),
        .ZN(inst2_stateArray_S11reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U662 ( .A1(inst2_n2435), .A2(ciphertext2[74]), .B1(
        plaintext2[82]), .B2(inst2_n2713), .ZN(inst2_n2432) );
  OAI21_X1 inst2_U661 ( .B1(inst2_n1262), .B2(inst2_n2711), .A(inst2_n2431),
        .ZN(inst2_stateArray_S11reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U660 ( .A1(inst2_n2435), .A2(ciphertext2[75]), .B1(
        plaintext2[83]), .B2(inst2_n2713), .ZN(inst2_n2431) );
  OAI21_X1 inst2_U659 ( .B1(inst2_n1250), .B2(inst2_n2711), .A(inst2_n2430),
        .ZN(inst2_stateArray_S12reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst2_U658 ( .A1(inst2_n2435), .A2(ciphertext2[71]), .B1(
        plaintext2[79]), .B2(inst2_n2582), .ZN(inst2_n2430) );
  OAI21_X1 inst2_U657 ( .B1(inst2_n1261), .B2(inst2_n2711), .A(inst2_n2429),
        .ZN(inst2_stateArray_S11reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U656 ( .A1(inst2_n2435), .A2(ciphertext2[76]), .B1(
        plaintext2[84]), .B2(inst2_n2722), .ZN(inst2_n2429) );
  OAI21_X1 inst2_U655 ( .B1(inst2_n1260), .B2(inst2_n2711), .A(inst2_n2428),
        .ZN(inst2_stateArray_S11reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst2_U654 ( .A1(inst2_n2435), .A2(ciphertext2[77]), .B1(
        plaintext2[85]), .B2(inst2_n2722), .ZN(inst2_n2428) );
  OAI21_X1 inst2_U653 ( .B1(inst2_n1259), .B2(inst2_n2711), .A(inst2_n2427),
        .ZN(inst2_stateArray_S11reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst2_U652 ( .A1(inst2_n2435), .A2(ciphertext2[78]), .B1(
        plaintext2[86]), .B2(inst2_n2722), .ZN(inst2_n2427) );
  OAI21_X1 inst2_U651 ( .B1(inst2_n1258), .B2(inst2_n2711), .A(inst2_n2426),
        .ZN(inst2_stateArray_S11reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst2_U650 ( .A1(inst2_n2435), .A2(ciphertext2[79]), .B1(
        plaintext2[87]), .B2(inst2_n2595), .ZN(inst2_n2426) );
  OAI21_X1 inst2_U649 ( .B1(inst2_n1257), .B2(inst2_n2711), .A(inst2_n2425),
        .ZN(inst2_stateArray_S12reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst2_U648 ( .A1(inst2_n2435), .A2(ciphertext2[64]), .B1(
        plaintext2[72]), .B2(inst2_n2550), .ZN(inst2_n2425) );
  OAI21_X1 inst2_U647 ( .B1(inst2_n1256), .B2(inst2_n2711), .A(inst2_n2424),
        .ZN(inst2_stateArray_S12reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U646 ( .A1(inst2_n2435), .A2(ciphertext2[65]), .B1(
        plaintext2[73]), .B2(inst2_n2713), .ZN(inst2_n2424) );
  OAI21_X1 inst2_U645 ( .B1(inst2_n1255), .B2(inst2_n2711), .A(inst2_n2423),
        .ZN(inst2_stateArray_S12reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U644 ( .A1(inst2_n2435), .A2(ciphertext2[66]), .B1(
        plaintext2[74]), .B2(inst2_n2722), .ZN(inst2_n2423) );
  INV_X1 inst2_U643 ( .A(inst2_n6), .ZN(inst2_n2722) );
  OAI21_X1 inst2_U642 ( .B1(inst2_n1254), .B2(inst2_n2711), .A(inst2_n2422),
        .ZN(inst2_stateArray_S12reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U641 ( .A1(inst2_n2435), .A2(ciphertext2[67]), .B1(
        plaintext2[75]), .B2(inst2_n2550), .ZN(inst2_n2422) );
  OAI21_X1 inst2_U640 ( .B1(inst2_n1253), .B2(inst2_n2711), .A(inst2_n2421),
        .ZN(inst2_stateArray_S12reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U639 ( .A1(inst2_n2435), .A2(ciphertext2[68]), .B1(
        plaintext2[76]), .B2(inst2_n2582), .ZN(inst2_n2421) );
  OAI21_X1 inst2_U638 ( .B1(inst2_n1252), .B2(inst2_n2711), .A(inst2_n2420),
        .ZN(inst2_stateArray_S12reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst2_U637 ( .A1(inst2_n2435), .A2(ciphertext2[69]), .B1(
        plaintext2[77]), .B2(inst2_n2713), .ZN(inst2_n2420) );
  OAI21_X1 inst2_U636 ( .B1(inst2_n1251), .B2(inst2_n2711), .A(inst2_n2419),
        .ZN(inst2_stateArray_S12reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst2_U635 ( .A1(inst2_n2435), .A2(ciphertext2[70]), .B1(
        plaintext2[78]), .B2(inst2_n2595), .ZN(inst2_n2419) );
  NOR2_X2 inst2_U634 ( .A1(done2), .A2(inst2_n2528), .ZN(inst2_n2435) );
  OAI211_X1 inst2_U633 ( .C1(inst2_n1176), .C2(inst2_n2115), .A(inst2_n2418),
        .B(inst2_n2417), .ZN(inst2_KeyArray_S33reg_gff_1_SFF_1_n5) );
  NAND2_X1 inst2_U632 ( .A1(inst2_n2543), .A2(inst2_n57), .ZN(inst2_n2417) );
  AOI22_X1 inst2_U631 ( .A1(inst2_n2375), .A2(inst2_n2813), .B1(key2[1]), .B2(
        inst2_n2713), .ZN(inst2_n2418) );
  OAI21_X1 inst2_U630 ( .B1(inst2_n1175), .B2(inst2_n2115), .A(inst2_n2416),
        .ZN(inst2_KeyArray_S33reg_gff_1_SFF_2_n5) );
  AOI21_X1 inst2_U629 ( .B1(key2[2]), .B2(inst2_n2582), .A(inst2_n2415), .ZN(
        inst2_n2416) );
  OAI22_X1 inst2_U628 ( .A1(inst2_n225), .A2(inst2_n2463), .B1(inst2_n1087),
        .B2(inst2_n2647), .ZN(inst2_n2415) );
  OAI21_X1 inst2_U627 ( .B1(inst2_n1174), .B2(inst2_n2652), .A(inst2_n2414),
        .ZN(inst2_KeyArray_S33reg_gff_1_SFF_3_n5) );
  AOI21_X1 inst2_U626 ( .B1(key2[3]), .B2(inst2_n2722), .A(inst2_n2413), .ZN(
        inst2_n2414) );
  OAI22_X1 inst2_U625 ( .A1(inst2_n224), .A2(inst2_n2463), .B1(inst2_n1086),
        .B2(inst2_n2647), .ZN(inst2_n2413) );
  OAI211_X1 inst2_U624 ( .C1(inst2_n1203), .C2(inst2_n2771), .A(inst2_n2412),
        .B(inst2_n2411), .ZN(inst2_stateArray_S31reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst2_U623 ( .A1(plaintext2[22]), .A2(inst2_n2713), .ZN(inst2_n2411) );
  AOI22_X1 inst2_U622 ( .A1(ciphertext2[22]), .A2(done2), .B1(inst2_n2791),
        .B2(ciphertext2[30]), .ZN(inst2_n2412) );
  OAI211_X1 inst2_U621 ( .C1(inst2_n1202), .C2(inst2_n2771), .A(inst2_n2410),
        .B(inst2_n2409), .ZN(inst2_stateArray_S31reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst2_U620 ( .A1(plaintext2[23]), .A2(inst2_n2582), .ZN(inst2_n2409) );
  AOI22_X1 inst2_U619 ( .A1(inst2_n2788), .A2(ciphertext2[23]), .B1(
        inst2_n2791), .B2(ciphertext2[31]), .ZN(inst2_n2410) );
  OAI21_X1 inst2_U618 ( .B1(inst2_n1220), .B2(inst2_n2771), .A(inst2_n2408),
        .ZN(inst2_stateArray_S22reg_gff_1_SFF_5_n6) );
  AOI21_X1 inst2_U617 ( .B1(plaintext2[45]), .B2(inst2_n2595), .A(inst2_n2407),
        .ZN(inst2_n2408) );
  OAI22_X1 inst2_U616 ( .A1(inst2_n1228), .A2(inst2_n2711), .B1(inst2_n2757),
        .B2(inst2_n2820), .ZN(inst2_n2407) );
  OAI21_X1 inst2_U615 ( .B1(inst2_n1177), .B2(inst2_n2652), .A(inst2_n2406),
        .ZN(inst2_KeyArray_S33reg_gff_1_SFF_0_n5) );
  AOI21_X1 inst2_U614 ( .B1(key2[0]), .B2(inst2_n2582), .A(inst2_n2405), .ZN(
        inst2_n2406) );
  OAI22_X1 inst2_U613 ( .A1(inst2_n227), .A2(inst2_n2463), .B1(inst2_n1089),
        .B2(inst2_n2647), .ZN(inst2_n2405) );
  OAI21_X1 inst2_U612 ( .B1(inst2_n1173), .B2(inst2_n2652), .A(inst2_n2404),
        .ZN(inst2_KeyArray_S33reg_gff_1_SFF_4_n5) );
  AOI21_X1 inst2_U611 ( .B1(key2[4]), .B2(inst2_n2582), .A(inst2_n2403), .ZN(
        inst2_n2404) );
  OAI22_X1 inst2_U610 ( .A1(inst2_n223), .A2(inst2_n2463), .B1(inst2_n1085),
        .B2(inst2_n2647), .ZN(inst2_n2403) );
  OAI21_X1 inst2_U609 ( .B1(inst2_n1172), .B2(inst2_n2652), .A(inst2_n2402),
        .ZN(inst2_KeyArray_S33reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst2_U608 ( .B1(key2[5]), .B2(inst2_n2582), .A(inst2_n2401), .ZN(
        inst2_n2402) );
  OAI22_X1 inst2_U607 ( .A1(inst2_n228), .A2(inst2_n2463), .B1(inst2_n1084),
        .B2(inst2_n2647), .ZN(inst2_n2401) );
  OAI21_X1 inst2_U606 ( .B1(inst2_n1171), .B2(inst2_n2652), .A(inst2_n2400),
        .ZN(inst2_KeyArray_S33reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst2_U605 ( .B1(key2[6]), .B2(inst2_n2582), .A(inst2_n2399), .ZN(
        inst2_n2400) );
  OAI22_X1 inst2_U604 ( .A1(inst2_n222), .A2(inst2_n2463), .B1(inst2_n1083),
        .B2(inst2_n2647), .ZN(inst2_n2399) );
  OAI21_X1 inst2_U603 ( .B1(inst2_n1170), .B2(inst2_n2115), .A(inst2_n2398),
        .ZN(inst2_KeyArray_S33reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst2_U602 ( .B1(key2[7]), .B2(inst2_n2582), .A(inst2_n2397), .ZN(
        inst2_n2398) );
  OAI22_X1 inst2_U601 ( .A1(inst2_n221), .A2(inst2_n2463), .B1(inst2_n1082),
        .B2(inst2_n2565), .ZN(inst2_n2397) );
  OAI211_X1 inst2_U600 ( .C1(inst2_n210), .C2(inst2_n2396), .A(inst2_n2395),
        .B(inst2_n2394), .ZN(inst2_stateArray_S03reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst2_U599 ( .A1(inst2_n2568), .A2(ciphertext2[88]), .B1(
        inst2_n2393), .B2(inst2_n2392), .ZN(inst2_n2394) );
  XNOR2_X1 inst2_U598 ( .A(inst2_n2782), .B(inst2_n2391), .ZN(inst2_n2392) );
  AOI22_X1 inst2_U597 ( .A1(inst2_n2390), .A2(ciphertext2[88]), .B1(inst2_n209), .B2(inst2_n2389), .ZN(inst2_n2391) );
  AOI22_X1 inst2_U596 ( .A1(inst2_n2586), .A2(ciphertext2[96]), .B1(
        plaintext2[96]), .B2(inst2_n2713), .ZN(inst2_n2395) );
  OAI211_X1 inst2_U595 ( .C1(inst2_n1169), .C2(inst2_n2115), .A(inst2_n2388),
        .B(inst2_n2387), .ZN(inst2_KeyArray_S00reg_gff_1_SFF_0_n6) );
  OAI21_X1 inst2_U594 ( .B1(inst2_n1193), .B2(inst2_n2386), .A(inst2_n2385),
        .ZN(inst2_n2387) );
  AOI21_X1 inst2_U593 ( .B1(inst2_n1193), .B2(inst2_n2386), .A(inst2_n2776),
        .ZN(inst2_n2385) );
  NAND2_X1 inst2_U592 ( .A1(inst2_n2384), .A2(inst2_n2819), .ZN(inst2_n2386)
         );
  AOI22_X1 inst2_U591 ( .A1(inst2_n2666), .A2(inst2_n2819), .B1(key2[120]),
        .B2(inst2_n2713), .ZN(inst2_n2388) );
  OAI211_X1 inst2_U590 ( .C1(inst2_n1168), .C2(inst2_n2652), .A(inst2_n2383),
        .B(inst2_n2382), .ZN(inst2_KeyArray_S00reg_gff_1_SFF_1_n6) );
  OAI21_X1 inst2_U589 ( .B1(inst2_n1192), .B2(inst2_n2381), .A(inst2_n2380),
        .ZN(inst2_n2382) );
  AOI21_X1 inst2_U588 ( .B1(inst2_n1192), .B2(inst2_n2381), .A(inst2_n2670),
        .ZN(inst2_n2380) );
  NAND2_X1 inst2_U587 ( .A1(inst2_n2384), .A2(inst2_n2813), .ZN(inst2_n2381)
         );
  AOI22_X1 inst2_U586 ( .A1(inst2_n2872), .A2(inst2_n2813), .B1(key2[121]),
        .B2(inst2_n2528), .ZN(inst2_n2383) );
  OAI211_X1 inst2_U585 ( .C1(inst2_n1167), .C2(inst2_n2115), .A(inst2_n2379),
        .B(inst2_n2378), .ZN(inst2_KeyArray_S00reg_gff_1_SFF_2_n6) );
  OAI21_X1 inst2_U584 ( .B1(inst2_n1191), .B2(inst2_n2377), .A(inst2_n2376),
        .ZN(inst2_n2378) );
  AOI21_X1 inst2_U583 ( .B1(inst2_n1191), .B2(inst2_n2377), .A(inst2_n2776),
        .ZN(inst2_n2376) );
  INV_X1 inst2_U582 ( .A(inst2_n2375), .ZN(inst2_n2776) );
  INV_X1 inst2_U581 ( .A(inst2_n2670), .ZN(inst2_n2375) );
  NAND2_X1 inst2_U580 ( .A1(inst2_n2384), .A2(inst2_n2814), .ZN(inst2_n2377)
         );
  AOI22_X1 inst2_U579 ( .A1(inst2_n2872), .A2(inst2_n2814), .B1(key2[122]),
        .B2(inst2_n2803), .ZN(inst2_n2379) );
  OAI211_X1 inst2_U578 ( .C1(inst2_n1166), .C2(inst2_n2652), .A(inst2_n2374),
        .B(inst2_n2373), .ZN(inst2_KeyArray_S00reg_gff_1_SFF_3_n6) );
  OAI21_X1 inst2_U577 ( .B1(inst2_n1190), .B2(inst2_n2372), .A(inst2_n2371),
        .ZN(inst2_n2373) );
  AOI21_X1 inst2_U576 ( .B1(inst2_n1190), .B2(inst2_n2372), .A(inst2_n2463),
        .ZN(inst2_n2371) );
  NAND2_X1 inst2_U575 ( .A1(inst2_n2384), .A2(inst2_n2818), .ZN(inst2_n2372)
         );
  AOI22_X1 inst2_U574 ( .A1(inst2_n2872), .A2(inst2_n2818), .B1(key2[123]),
        .B2(inst2_n2803), .ZN(inst2_n2374) );
  OAI211_X1 inst2_U573 ( .C1(inst2_n1165), .C2(inst2_n2652), .A(inst2_n2370),
        .B(inst2_n2369), .ZN(inst2_KeyArray_S00reg_gff_1_SFF_4_n6) );
  OAI21_X1 inst2_U572 ( .B1(inst2_n1189), .B2(inst2_n2368), .A(inst2_n2367),
        .ZN(inst2_n2369) );
  AOI21_X1 inst2_U571 ( .B1(inst2_n1189), .B2(inst2_n2368), .A(inst2_n2670),
        .ZN(inst2_n2367) );
  NAND2_X1 inst2_U570 ( .A1(inst2_n2384), .A2(inst2_n2817), .ZN(inst2_n2368)
         );
  AOI22_X1 inst2_U569 ( .A1(inst2_n2666), .A2(inst2_n2817), .B1(key2[124]),
        .B2(inst2_n2803), .ZN(inst2_n2370) );
  OAI211_X1 inst2_U568 ( .C1(inst2_n1164), .C2(inst2_n2115), .A(inst2_n2366),
        .B(inst2_n2365), .ZN(inst2_KeyArray_S00reg_gff_1_SFF_5_n6) );
  OAI21_X1 inst2_U567 ( .B1(inst2_n1188), .B2(inst2_n2364), .A(inst2_n2363),
        .ZN(inst2_n2365) );
  AOI21_X1 inst2_U566 ( .B1(inst2_n1188), .B2(inst2_n2364), .A(inst2_n2776),
        .ZN(inst2_n2363) );
  NAND2_X1 inst2_U565 ( .A1(inst2_n2384), .A2(inst2_n2816), .ZN(inst2_n2364)
         );
  AOI22_X1 inst2_U564 ( .A1(inst2_n2543), .A2(inst2_n2816), .B1(key2[125]),
        .B2(inst2_n2803), .ZN(inst2_n2366) );
  INV_X1 inst2_U563 ( .A(inst2_n2796), .ZN(inst2_n2543) );
  OAI211_X1 inst2_U562 ( .C1(inst2_n1163), .C2(inst2_n2652), .A(inst2_n2362),
        .B(inst2_n2361), .ZN(inst2_KeyArray_S00reg_gff_1_SFF_6_n6) );
  OAI21_X1 inst2_U561 ( .B1(inst2_n1187), .B2(inst2_n2360), .A(inst2_n2359),
        .ZN(inst2_n2361) );
  AOI21_X1 inst2_U560 ( .B1(inst2_n1187), .B2(inst2_n2360), .A(inst2_n2776),
        .ZN(inst2_n2359) );
  NAND2_X1 inst2_U559 ( .A1(inst2_n2384), .A2(inst2_n2815), .ZN(inst2_n2360)
         );
  AOI22_X1 inst2_U558 ( .A1(inst2_n2666), .A2(inst2_n2815), .B1(key2[126]),
        .B2(inst2_n2803), .ZN(inst2_n2362) );
  OAI211_X1 inst2_U557 ( .C1(inst2_n1162), .C2(inst2_n2652), .A(inst2_n2358),
        .B(inst2_n2357), .ZN(inst2_KeyArray_S00reg_gff_1_SFF_7_n6) );
  OAI21_X1 inst2_U556 ( .B1(inst2_n1186), .B2(inst2_n2356), .A(inst2_n2355),
        .ZN(inst2_n2357) );
  AOI21_X1 inst2_U555 ( .B1(inst2_n1186), .B2(inst2_n2356), .A(inst2_n2463),
        .ZN(inst2_n2355) );
  NAND2_X1 inst2_U554 ( .A1(inst2_n2384), .A2(inst2_n2802), .ZN(inst2_n2356)
         );
  AOI22_X1 inst2_U553 ( .A1(inst2_n2354), .A2(inst2_n2353), .B1(inst2_n236),
        .B2(inst2_n2811), .ZN(inst2_n2384) );
  AND4_X1 inst2_U552 ( .A1(inst2_n2801), .A2(inst2_n2812), .A3(inst2_n2837),
        .A4(inst2_n718), .ZN(inst2_n2353) );
  AND4_X1 inst2_U551 ( .A1(inst2_n2836), .A2(inst2_n499), .A3(inst2_n1081),
        .A4(inst2_n1080), .ZN(inst2_n2354) );
  AOI22_X1 inst2_U550 ( .A1(inst2_n2666), .A2(inst2_n2802), .B1(key2[127]),
        .B2(inst2_n2803), .ZN(inst2_n2358) );
  OAI211_X1 inst2_U549 ( .C1(inst2_n1206), .C2(inst2_n2771), .A(inst2_n2352),
        .B(inst2_n2351), .ZN(inst2_stateArray_S31reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst2_U548 ( .A1(plaintext2[19]), .A2(inst2_n2550), .ZN(inst2_n2351) );
  AOI22_X1 inst2_U547 ( .A1(inst2_n2788), .A2(ciphertext2[19]), .B1(
        inst2_n2791), .B2(ciphertext2[27]), .ZN(inst2_n2352) );
  OAI211_X1 inst2_U546 ( .C1(inst2_n198), .C2(inst2_n2396), .A(inst2_n2350),
        .B(inst2_n2349), .ZN(inst2_stateArray_S03reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U545 ( .A1(inst2_n2375), .A2(ciphertext2[89]), .B1(
        inst2_n2393), .B2(inst2_n2348), .ZN(inst2_n2349) );
  XNOR2_X1 inst2_U544 ( .A(inst2_n2347), .B(inst2_n2346), .ZN(inst2_n2348) );
  AOI22_X1 inst2_U543 ( .A1(inst2_n2390), .A2(ciphertext2[89]), .B1(inst2_n197), .B2(inst2_n2389), .ZN(inst2_n2346) );
  AOI22_X1 inst2_U542 ( .A1(inst2_n2345), .A2(inst2_n2772), .B1(inst2_n2773),
        .B2(inst2_n2344), .ZN(inst2_n2347) );
  INV_X1 inst2_U541 ( .A(inst2_n2345), .ZN(inst2_n2344) );
  INV_X1 inst2_U540 ( .A(inst2_n2772), .ZN(inst2_n2773) );
  AOI22_X1 inst2_U539 ( .A1(inst2_n2872), .A2(ciphertext2[97]), .B1(
        plaintext2[97]), .B2(inst2_n2803), .ZN(inst2_n2350) );
  OAI211_X1 inst2_U538 ( .C1(inst2_n202), .C2(inst2_n2396), .A(inst2_n2343),
        .B(inst2_n2342), .ZN(inst2_stateArray_S03reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U537 ( .A1(inst2_n2614), .A2(ciphertext2[91]), .B1(
        inst2_n2393), .B2(inst2_n2341), .ZN(inst2_n2342) );
  XNOR2_X1 inst2_U536 ( .A(inst2_n2340), .B(inst2_n2339), .ZN(inst2_n2341) );
  AOI22_X1 inst2_U535 ( .A1(inst2_n201), .A2(inst2_n2390), .B1(inst2_n2389),
        .B2(ciphertext2[91]), .ZN(inst2_n2339) );
  AOI22_X1 inst2_U534 ( .A1(inst2_n2775), .A2(inst2_n2762), .B1(inst2_n2761),
        .B2(inst2_n2338), .ZN(inst2_n2340) );
  INV_X1 inst2_U533 ( .A(inst2_n2775), .ZN(inst2_n2338) );
  INV_X1 inst2_U532 ( .A(inst2_n2762), .ZN(inst2_n2761) );
  AOI22_X1 inst2_U531 ( .A1(inst2_n2666), .A2(ciphertext2[99]), .B1(
        plaintext2[99]), .B2(inst2_n2803), .ZN(inst2_n2343) );
  OAI211_X1 inst2_U530 ( .C1(inst2_n216), .C2(inst2_n2396), .A(inst2_n2337),
        .B(inst2_n2336), .ZN(inst2_stateArray_S03reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst2_U529 ( .A1(inst2_n2122), .A2(ciphertext2[94]), .B1(
        inst2_n2393), .B2(inst2_n2335), .ZN(inst2_n2336) );
  XNOR2_X1 inst2_U528 ( .A(inst2_n2334), .B(inst2_n2333), .ZN(inst2_n2335) );
  AOI22_X1 inst2_U527 ( .A1(inst2_n214), .A2(ciphertext2[30]), .B1(inst2_n215),
        .B2(ciphertext2[125]), .ZN(inst2_n2333) );
  AOI22_X1 inst2_U526 ( .A1(inst2_n2332), .A2(inst2_n190), .B1(ciphertext2[93]), .B2(inst2_n2331), .ZN(inst2_n2334) );
  INV_X1 inst2_U525 ( .A(inst2_n2332), .ZN(inst2_n2331) );
  AOI22_X1 inst2_U524 ( .A1(inst2_n2872), .A2(ciphertext2[102]), .B1(
        plaintext2[102]), .B2(inst2_n2803), .ZN(inst2_n2337) );
  OAI211_X1 inst2_U523 ( .C1(inst2_n2800), .C2(inst2_n2396), .A(inst2_n2330),
        .B(inst2_n2329), .ZN(inst2_stateArray_S03reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U522 ( .A1(inst2_n2122), .A2(ciphertext2[90]), .B1(
        inst2_n2393), .B2(inst2_n2328), .ZN(inst2_n2329) );
  XNOR2_X1 inst2_U521 ( .A(inst2_n2327), .B(inst2_n2326), .ZN(inst2_n2328) );
  AOI22_X1 inst2_U520 ( .A1(inst2_n203), .A2(inst2_n2783), .B1(inst2_n2325),
        .B2(ciphertext2[26]), .ZN(inst2_n2326) );
  INV_X1 inst2_U519 ( .A(inst2_n2783), .ZN(inst2_n2325) );
  AOI22_X1 inst2_U518 ( .A1(inst2_n2666), .A2(ciphertext2[98]), .B1(
        plaintext2[98]), .B2(inst2_n2803), .ZN(inst2_n2330) );
  OAI211_X1 inst2_U517 ( .C1(inst2_n214), .C2(inst2_n2396), .A(inst2_n2324),
        .B(inst2_n2323), .ZN(inst2_stateArray_S03reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst2_U516 ( .A1(inst2_n2568), .A2(ciphertext2[93]), .B1(
        inst2_n2393), .B2(inst2_n2322), .ZN(inst2_n2323) );
  XNOR2_X1 inst2_U515 ( .A(inst2_n2321), .B(inst2_n2320), .ZN(inst2_n2322) );
  AOI22_X1 inst2_U514 ( .A1(ciphertext2[124]), .A2(inst2_n2804), .B1(
        ciphertext2[29]), .B2(inst2_n2799), .ZN(inst2_n2320) );
  AOI22_X1 inst2_U513 ( .A1(inst2_n212), .A2(inst2_n2319), .B1(inst2_n2318),
        .B2(ciphertext2[92]), .ZN(inst2_n2321) );
  INV_X1 inst2_U512 ( .A(inst2_n2319), .ZN(inst2_n2318) );
  AOI22_X1 inst2_U511 ( .A1(inst2_n2666), .A2(ciphertext2[101]), .B1(
        plaintext2[101]), .B2(inst2_n2803), .ZN(inst2_n2324) );
  OAI211_X1 inst2_U510 ( .C1(inst2_n2799), .C2(inst2_n2396), .A(inst2_n2317),
        .B(inst2_n2316), .ZN(inst2_stateArray_S03reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U509 ( .A1(inst2_n2614), .A2(ciphertext2[92]), .B1(
        inst2_n2393), .B2(inst2_n2315), .ZN(inst2_n2316) );
  XNOR2_X1 inst2_U508 ( .A(inst2_n2314), .B(inst2_n2313), .ZN(inst2_n2315) );
  AOI22_X1 inst2_U507 ( .A1(inst2_n207), .A2(inst2_n2312), .B1(inst2_n2311),
        .B2(ciphertext2[28]), .ZN(inst2_n2313) );
  INV_X1 inst2_U506 ( .A(inst2_n2311), .ZN(inst2_n2312) );
  AOI22_X1 inst2_U505 ( .A1(inst2_n2310), .A2(inst2_n2390), .B1(inst2_n2389),
        .B2(inst2_n2309), .ZN(inst2_n2314) );
  AOI22_X1 inst2_U504 ( .A1(inst2_n2586), .A2(ciphertext2[100]), .B1(
        plaintext2[100]), .B2(inst2_n2528), .ZN(inst2_n2317) );
  OAI211_X1 inst2_U503 ( .C1(inst2_n1208), .C2(inst2_n2771), .A(inst2_n2308),
        .B(inst2_n2307), .ZN(inst2_stateArray_S31reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst2_U502 ( .A1(plaintext2[17]), .A2(inst2_n2595), .ZN(inst2_n2307) );
  AOI22_X1 inst2_U501 ( .A1(done2), .A2(ciphertext2[17]), .B1(inst2_n2791),
        .B2(ciphertext2[25]), .ZN(inst2_n2308) );
  OAI211_X1 inst2_U500 ( .C1(inst2_n1209), .C2(inst2_n2771), .A(inst2_n2306),
        .B(inst2_n2305), .ZN(inst2_stateArray_S31reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst2_U499 ( .A1(plaintext2[16]), .A2(inst2_n2722), .ZN(inst2_n2305) );
  AOI22_X1 inst2_U498 ( .A1(inst2_n2788), .A2(ciphertext2[16]), .B1(
        inst2_n2791), .B2(ciphertext2[24]), .ZN(inst2_n2306) );
  OAI211_X1 inst2_U497 ( .C1(inst2_n218), .C2(inst2_n2396), .A(inst2_n2304),
        .B(inst2_n2303), .ZN(inst2_stateArray_S03reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst2_U496 ( .A1(inst2_n2375), .A2(ciphertext2[95]), .B1(
        inst2_n2393), .B2(inst2_n2302), .ZN(inst2_n2303) );
  XNOR2_X1 inst2_U495 ( .A(inst2_n2301), .B(inst2_n2300), .ZN(inst2_n2302) );
  AOI22_X1 inst2_U494 ( .A1(inst2_n216), .A2(ciphertext2[94]), .B1(inst2_n206),
        .B2(ciphertext2[126]), .ZN(inst2_n2300) );
  AOI22_X1 inst2_U493 ( .A1(inst2_n220), .A2(inst2_n2785), .B1(inst2_n2784),
        .B2(ciphertext2[95]), .ZN(inst2_n2301) );
  AOI22_X1 inst2_U492 ( .A1(inst2_n2586), .A2(ciphertext2[103]), .B1(
        plaintext2[103]), .B2(inst2_n2507), .ZN(inst2_n2304) );
  OAI211_X1 inst2_U491 ( .C1(inst2_n1207), .C2(inst2_n2771), .A(inst2_n2299),
        .B(inst2_n2298), .ZN(inst2_stateArray_S31reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst2_U490 ( .A1(plaintext2[18]), .A2(inst2_n2550), .ZN(inst2_n2298) );
  AOI22_X1 inst2_U489 ( .A1(inst2_n2788), .A2(ciphertext2[18]), .B1(
        inst2_n2791), .B2(ciphertext2[26]), .ZN(inst2_n2299) );
  OAI211_X1 inst2_U488 ( .C1(inst2_n1205), .C2(inst2_n2771), .A(inst2_n2297),
        .B(inst2_n2296), .ZN(inst2_stateArray_S31reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst2_U487 ( .A1(plaintext2[20]), .A2(inst2_n2582), .ZN(inst2_n2296) );
  AOI22_X1 inst2_U486 ( .A1(inst2_n2788), .A2(ciphertext2[20]), .B1(
        inst2_n2791), .B2(ciphertext2[28]), .ZN(inst2_n2297) );
  OAI211_X1 inst2_U485 ( .C1(inst2_n2794), .C2(inst2_n2295), .A(inst2_n2294),
        .B(inst2_n2293), .ZN(inst2_stateArray_S13reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst2_U484 ( .A1(inst2_n2375), .A2(ciphertext2[56]), .B1(
        ciphertext2[88]), .B2(inst2_n2292), .ZN(inst2_n2293) );
  AOI22_X1 inst2_U483 ( .A1(done2), .A2(ciphertext2[64]), .B1(plaintext2[64]),
        .B2(inst2_n2657), .ZN(inst2_n2294) );
  XNOR2_X1 inst2_U482 ( .A(inst2_n2782), .B(inst2_n2291), .ZN(inst2_n2295) );
  AOI22_X1 inst2_U481 ( .A1(inst2_n210), .A2(inst2_n2290), .B1(inst2_n2289),
        .B2(ciphertext2[120]), .ZN(inst2_n2291) );
  AOI22_X1 inst2_U480 ( .A1(inst2_n199), .A2(ciphertext2[56]), .B1(inst2_n2808), .B2(ciphertext2[24]), .ZN(inst2_n2782) );
  OAI211_X1 inst2_U479 ( .C1(inst2_n2288), .C2(inst2_n2780), .A(inst2_n2287),
        .B(inst2_n2286), .ZN(inst2_stateArray_S13reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U478 ( .A1(inst2_n2568), .A2(ciphertext2[57]), .B1(
        ciphertext2[89]), .B2(inst2_n2292), .ZN(inst2_n2286) );
  AOI22_X1 inst2_U477 ( .A1(done2), .A2(ciphertext2[65]), .B1(plaintext2[65]),
        .B2(inst2_n2713), .ZN(inst2_n2287) );
  XNOR2_X1 inst2_U476 ( .A(inst2_n2285), .B(inst2_n2284), .ZN(inst2_n2288) );
  AOI22_X1 inst2_U475 ( .A1(inst2_n209), .A2(inst2_n2290), .B1(inst2_n2289),
        .B2(ciphertext2[88]), .ZN(inst2_n2284) );
  XNOR2_X1 inst2_U474 ( .A(inst2_n2772), .B(inst2_n2283), .ZN(inst2_n2285) );
  AOI22_X1 inst2_U473 ( .A1(inst2_n198), .A2(ciphertext2[56]), .B1(inst2_n2808), .B2(ciphertext2[121]), .ZN(inst2_n2283) );
  AOI22_X1 inst2_U472 ( .A1(inst2_n191), .A2(ciphertext2[57]), .B1(inst2_n2810), .B2(ciphertext2[25]), .ZN(inst2_n2772) );
  OAI211_X1 inst2_U471 ( .C1(inst2_n2282), .C2(inst2_n2780), .A(inst2_n2281),
        .B(inst2_n2280), .ZN(inst2_stateArray_S13reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U470 ( .A1(inst2_n2614), .A2(ciphertext2[58]), .B1(
        ciphertext2[90]), .B2(inst2_n2292), .ZN(inst2_n2280) );
  AOI22_X1 inst2_U469 ( .A1(done2), .A2(ciphertext2[66]), .B1(plaintext2[66]),
        .B2(inst2_n2713), .ZN(inst2_n2281) );
  XNOR2_X1 inst2_U468 ( .A(inst2_n2279), .B(inst2_n2278), .ZN(inst2_n2282) );
  AOI22_X1 inst2_U467 ( .A1(inst2_n197), .A2(ciphertext2[57]), .B1(inst2_n2810), .B2(ciphertext2[89]), .ZN(inst2_n2278) );
  XNOR2_X1 inst2_U466 ( .A(inst2_n2277), .B(inst2_n193), .ZN(inst2_n2279) );
  OAI211_X1 inst2_U465 ( .C1(inst2_n2794), .C2(inst2_n2276), .A(inst2_n2275),
        .B(inst2_n2274), .ZN(inst2_stateArray_S13reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U464 ( .A1(inst2_n2614), .A2(ciphertext2[59]), .B1(
        ciphertext2[91]), .B2(inst2_n2292), .ZN(inst2_n2274) );
  AOI22_X1 inst2_U463 ( .A1(done2), .A2(ciphertext2[67]), .B1(plaintext2[67]),
        .B2(inst2_n2713), .ZN(inst2_n2275) );
  XNOR2_X1 inst2_U462 ( .A(inst2_n2273), .B(inst2_n2272), .ZN(inst2_n2276) );
  AOI22_X1 inst2_U461 ( .A1(inst2_n202), .A2(inst2_n2289), .B1(inst2_n2290),
        .B2(ciphertext2[123]), .ZN(inst2_n2272) );
  INV_X1 inst2_U460 ( .A(inst2_n2290), .ZN(inst2_n2289) );
  XNOR2_X1 inst2_U459 ( .A(inst2_n2762), .B(inst2_n2327), .ZN(inst2_n2273) );
  AOI22_X1 inst2_U458 ( .A1(inst2_n194), .A2(inst2_n193), .B1(ciphertext2[58]),
        .B2(ciphertext2[90]), .ZN(inst2_n2327) );
  AOI22_X1 inst2_U457 ( .A1(ciphertext2[27]), .A2(inst2_n196), .B1(
        ciphertext2[59]), .B2(inst2_n2806), .ZN(inst2_n2762) );
  OAI211_X1 inst2_U456 ( .C1(inst2_n2271), .C2(inst2_n2794), .A(inst2_n2270),
        .B(inst2_n2269), .ZN(inst2_stateArray_S13reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U455 ( .A1(inst2_n2122), .A2(ciphertext2[60]), .B1(
        ciphertext2[92]), .B2(inst2_n2292), .ZN(inst2_n2269) );
  AOI22_X1 inst2_U454 ( .A1(done2), .A2(ciphertext2[68]), .B1(plaintext2[68]),
        .B2(inst2_n2484), .ZN(inst2_n2270) );
  XNOR2_X1 inst2_U453 ( .A(inst2_n2268), .B(inst2_n2267), .ZN(inst2_n2271) );
  AOI22_X1 inst2_U452 ( .A1(inst2_n201), .A2(inst2_n2764), .B1(inst2_n2763),
        .B2(ciphertext2[91]), .ZN(inst2_n2267) );
  INV_X1 inst2_U451 ( .A(inst2_n2764), .ZN(inst2_n2763) );
  XNOR2_X1 inst2_U450 ( .A(inst2_n2290), .B(inst2_n2266), .ZN(inst2_n2268) );
  AOI22_X1 inst2_U449 ( .A1(ciphertext2[60]), .A2(inst2_n196), .B1(
        ciphertext2[59]), .B2(inst2_n2809), .ZN(inst2_n2266) );
  AOI22_X1 inst2_U448 ( .A1(inst2_n219), .A2(inst2_n220), .B1(ciphertext2[95]),
        .B2(ciphertext2[63]), .ZN(inst2_n2290) );
  OAI211_X1 inst2_U447 ( .C1(inst2_n2794), .C2(inst2_n2265), .A(inst2_n2264),
        .B(inst2_n2263), .ZN(inst2_stateArray_S13reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst2_U446 ( .A1(inst2_n2122), .A2(ciphertext2[61]), .B1(
        ciphertext2[93]), .B2(inst2_n2292), .ZN(inst2_n2263) );
  AOI22_X1 inst2_U445 ( .A1(inst2_n2788), .A2(ciphertext2[69]), .B1(
        plaintext2[69]), .B2(inst2_n2713), .ZN(inst2_n2264) );
  XNOR2_X1 inst2_U444 ( .A(inst2_n2311), .B(inst2_n2262), .ZN(inst2_n2265) );
  AOI22_X1 inst2_U443 ( .A1(inst2_n2261), .A2(ciphertext2[61]), .B1(
        inst2_n2820), .B2(inst2_n2260), .ZN(inst2_n2262) );
  OAI211_X1 inst2_U442 ( .C1(inst2_n2259), .C2(inst2_n2794), .A(inst2_n2258),
        .B(inst2_n2257), .ZN(inst2_stateArray_S13reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst2_U441 ( .A1(inst2_n2614), .A2(ciphertext2[62]), .B1(
        ciphertext2[94]), .B2(inst2_n2292), .ZN(inst2_n2257) );
  AOI22_X1 inst2_U440 ( .A1(inst2_n2788), .A2(ciphertext2[70]), .B1(
        plaintext2[70]), .B2(inst2_n2484), .ZN(inst2_n2258) );
  XNOR2_X1 inst2_U439 ( .A(inst2_n2319), .B(inst2_n2256), .ZN(inst2_n2259) );
  AOI22_X1 inst2_U438 ( .A1(ciphertext2[62]), .A2(inst2_n2255), .B1(
        inst2_n2254), .B2(inst2_n2807), .ZN(inst2_n2256) );
  OAI211_X1 inst2_U437 ( .C1(inst2_n2253), .C2(inst2_n2794), .A(inst2_n2252),
        .B(inst2_n2251), .ZN(inst2_stateArray_S13reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst2_U436 ( .A1(inst2_n2375), .A2(ciphertext2[63]), .B1(
        ciphertext2[95]), .B2(inst2_n2292), .ZN(inst2_n2251) );
  NAND2_X1 inst2_U435 ( .A1(inst2_n2789), .A2(inst2_n2760), .ZN(inst2_n2292)
         );
  AOI22_X1 inst2_U434 ( .A1(done2), .A2(ciphertext2[71]), .B1(plaintext2[71]),
        .B2(inst2_n2657), .ZN(inst2_n2252) );
  XNOR2_X1 inst2_U433 ( .A(inst2_n2332), .B(inst2_n2250), .ZN(inst2_n2253) );
  AOI22_X1 inst2_U432 ( .A1(inst2_n218), .A2(inst2_n2784), .B1(inst2_n2785),
        .B2(ciphertext2[127]), .ZN(inst2_n2250) );
  OAI211_X1 inst2_U431 ( .C1(inst2_n2791), .C2(inst2_n444), .A(inst2_n6), .B(
        inst2_n2249), .ZN(inst2_calcRCon_n51) );
  NAND2_X1 inst2_U430 ( .A1(inst2_n2791), .A2(inst2_n2801), .ZN(inst2_n2249)
         );
  OAI221_X1 inst2_U429 ( .B1(inst2_n2791), .B2(inst2_n581), .C1(inst2_n2760),
        .C2(inst2_n499), .A(inst2_n6), .ZN(inst2_calcRCon_n49) );
  OAI221_X1 inst2_U428 ( .B1(inst2_n2791), .B2(inst2_n1071), .C1(inst2_n2757),
        .C2(inst2_n718), .A(inst2_n6), .ZN(inst2_calcRCon_n44) );
  OAI21_X1 inst2_U427 ( .B1(inst2_n210), .B2(inst2_n2647), .A(inst2_n2248),
        .ZN(inst2_stateArray_S00reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst2_U426 ( .A1(ciphertext2[112]), .A2(inst2_n1917), .B1(
        plaintext2[120]), .B2(inst2_n2722), .ZN(inst2_n2248) );
  OAI21_X1 inst2_U425 ( .B1(inst2_n198), .B2(inst2_n2647), .A(inst2_n2247),
        .ZN(inst2_stateArray_S00reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U424 ( .A1(ciphertext2[113]), .A2(inst2_n1917), .B1(
        plaintext2[121]), .B2(inst2_n2484), .ZN(inst2_n2247) );
  OAI21_X1 inst2_U423 ( .B1(inst2_n2647), .B2(inst2_n2800), .A(inst2_n2246),
        .ZN(inst2_stateArray_S00reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U422 ( .A1(ciphertext2[114]), .A2(inst2_n1917), .B1(
        plaintext2[122]), .B2(inst2_n2595), .ZN(inst2_n2246) );
  OAI21_X1 inst2_U421 ( .B1(inst2_n202), .B2(inst2_n2565), .A(inst2_n2245),
        .ZN(inst2_stateArray_S00reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U420 ( .A1(ciphertext2[115]), .A2(inst2_n1917), .B1(
        plaintext2[123]), .B2(inst2_n2657), .ZN(inst2_n2245) );
  OAI21_X1 inst2_U419 ( .B1(inst2_n2565), .B2(inst2_n2799), .A(inst2_n2244),
        .ZN(inst2_stateArray_S00reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U418 ( .A1(ciphertext2[116]), .A2(inst2_n1917), .B1(
        plaintext2[124]), .B2(inst2_n2722), .ZN(inst2_n2244) );
  OAI21_X1 inst2_U417 ( .B1(inst2_n214), .B2(inst2_n2565), .A(inst2_n2243),
        .ZN(inst2_stateArray_S00reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst2_U416 ( .A1(ciphertext2[117]), .A2(inst2_n1917), .B1(
        plaintext2[125]), .B2(inst2_n2713), .ZN(inst2_n2243) );
  OAI21_X1 inst2_U415 ( .B1(inst2_n216), .B2(inst2_n2565), .A(inst2_n2242),
        .ZN(inst2_stateArray_S00reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst2_U414 ( .A1(ciphertext2[118]), .A2(inst2_n1917), .B1(
        plaintext2[126]), .B2(inst2_n2582), .ZN(inst2_n2242) );
  OAI21_X1 inst2_U413 ( .B1(inst2_n218), .B2(inst2_n2565), .A(inst2_n2241),
        .ZN(inst2_stateArray_S00reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst2_U412 ( .A1(ciphertext2[119]), .A2(inst2_n1917), .B1(
        plaintext2[127]), .B2(inst2_n2528), .ZN(inst2_n2241) );
  OAI21_X1 inst2_U411 ( .B1(inst2_n2796), .B2(inst2_n2862), .A(inst2_n2240),
        .ZN(inst2_stateArray_S01reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst2_U410 ( .A1(ciphertext2[104]), .A2(inst2_n1917), .B1(
        plaintext2[112]), .B2(inst2_n2507), .ZN(inst2_n2240) );
  OAI21_X1 inst2_U409 ( .B1(inst2_n2796), .B2(inst2_n2861), .A(inst2_n2239),
        .ZN(inst2_stateArray_S01reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U408 ( .A1(ciphertext2[105]), .A2(inst2_n1917), .B1(
        plaintext2[113]), .B2(inst2_n2550), .ZN(inst2_n2239) );
  OAI21_X1 inst2_U407 ( .B1(inst2_n2565), .B2(inst2_n2860), .A(inst2_n2238),
        .ZN(inst2_stateArray_S01reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U406 ( .A1(ciphertext2[106]), .A2(inst2_n1917), .B1(
        plaintext2[114]), .B2(inst2_n2582), .ZN(inst2_n2238) );
  OAI21_X1 inst2_U405 ( .B1(inst2_n2796), .B2(inst2_n2859), .A(inst2_n2237),
        .ZN(inst2_stateArray_S01reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U404 ( .A1(ciphertext2[107]), .A2(inst2_n1917), .B1(
        plaintext2[115]), .B2(inst2_n2595), .ZN(inst2_n2237) );
  OAI21_X1 inst2_U403 ( .B1(inst2_n2565), .B2(inst2_n2858), .A(inst2_n2236),
        .ZN(inst2_stateArray_S01reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U402 ( .A1(ciphertext2[108]), .A2(inst2_n1917), .B1(
        plaintext2[116]), .B2(inst2_n2550), .ZN(inst2_n2236) );
  OAI21_X1 inst2_U401 ( .B1(inst2_n2565), .B2(inst2_n2857), .A(inst2_n2235),
        .ZN(inst2_stateArray_S01reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst2_U400 ( .A1(ciphertext2[109]), .A2(inst2_n1917), .B1(
        plaintext2[117]), .B2(inst2_n2550), .ZN(inst2_n2235) );
  OAI21_X1 inst2_U399 ( .B1(inst2_n2565), .B2(inst2_n2856), .A(inst2_n2234),
        .ZN(inst2_stateArray_S01reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst2_U398 ( .A1(ciphertext2[110]), .A2(inst2_n1917), .B1(
        plaintext2[118]), .B2(inst2_n2595), .ZN(inst2_n2234) );
  OAI21_X1 inst2_U397 ( .B1(inst2_n2565), .B2(inst2_n2855), .A(inst2_n2233),
        .ZN(inst2_stateArray_S01reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst2_U396 ( .A1(ciphertext2[111]), .A2(inst2_n1917), .B1(
        plaintext2[119]), .B2(inst2_n2722), .ZN(inst2_n2233) );
  OAI21_X1 inst2_U395 ( .B1(inst2_n1273), .B2(inst2_n2771), .A(inst2_n2232),
        .ZN(inst2_stateArray_S02reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst2_U394 ( .A1(ciphertext2[104]), .A2(inst2_n2872), .B1(
        plaintext2[104]), .B2(inst2_n2657), .ZN(inst2_n2232) );
  OAI21_X1 inst2_U393 ( .B1(inst2_n1272), .B2(inst2_n2771), .A(inst2_n2231),
        .ZN(inst2_stateArray_S02reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst2_U392 ( .A1(ciphertext2[105]), .A2(inst2_n2872), .B1(
        plaintext2[105]), .B2(inst2_n2507), .ZN(inst2_n2231) );
  OAI21_X1 inst2_U391 ( .B1(inst2_n1271), .B2(inst2_n2771), .A(inst2_n2230),
        .ZN(inst2_stateArray_S02reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst2_U390 ( .A1(ciphertext2[106]), .A2(inst2_n2666), .B1(
        plaintext2[106]), .B2(inst2_n2507), .ZN(inst2_n2230) );
  OAI21_X1 inst2_U389 ( .B1(inst2_n1270), .B2(inst2_n2771), .A(inst2_n2229),
        .ZN(inst2_stateArray_S02reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst2_U388 ( .A1(ciphertext2[107]), .A2(inst2_n2872), .B1(
        plaintext2[107]), .B2(inst2_n2484), .ZN(inst2_n2229) );
  OAI21_X1 inst2_U387 ( .B1(inst2_n1269), .B2(inst2_n2771), .A(inst2_n2228),
        .ZN(inst2_stateArray_S02reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst2_U386 ( .A1(ciphertext2[108]), .A2(inst2_n2872), .B1(
        plaintext2[108]), .B2(inst2_n2528), .ZN(inst2_n2228) );
  OAI21_X1 inst2_U385 ( .B1(inst2_n1268), .B2(inst2_n2771), .A(inst2_n2227),
        .ZN(inst2_stateArray_S02reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst2_U384 ( .A1(ciphertext2[109]), .A2(inst2_n2098), .B1(
        plaintext2[109]), .B2(inst2_n2657), .ZN(inst2_n2227) );
  OAI21_X1 inst2_U383 ( .B1(inst2_n1267), .B2(inst2_n2771), .A(inst2_n2226),
        .ZN(inst2_stateArray_S02reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst2_U382 ( .A1(ciphertext2[110]), .A2(inst2_n2098), .B1(
        plaintext2[110]), .B2(inst2_n2713), .ZN(inst2_n2226) );
  OAI21_X1 inst2_U381 ( .B1(inst2_n1266), .B2(inst2_n2771), .A(inst2_n2225),
        .ZN(inst2_stateArray_S02reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst2_U380 ( .A1(ciphertext2[111]), .A2(inst2_n2098), .B1(
        plaintext2[111]), .B2(inst2_n2484), .ZN(inst2_n2225) );
  OAI211_X1 inst2_U379 ( .C1(inst2_n2794), .C2(inst2_n2224), .A(inst2_n2223),
        .B(inst2_n2222), .ZN(inst2_stateArray_S23reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst2_U378 ( .B1(inst2_n2791), .B2(ciphertext2[48]), .A(inst2_n2221), .ZN(inst2_n2222) );
  OAI22_X1 inst2_U377 ( .A1(inst2_n199), .A2(inst2_n2463), .B1(inst2_n2396),
        .B2(inst2_n2808), .ZN(inst2_n2221) );
  AOI22_X1 inst2_U376 ( .A1(done2), .A2(ciphertext2[32]), .B1(plaintext2[32]),
        .B2(inst2_n2582), .ZN(inst2_n2223) );
  XNOR2_X1 inst2_U375 ( .A(inst2_n2345), .B(inst2_n2220), .ZN(inst2_n2224) );
  AOI22_X1 inst2_U374 ( .A1(inst2_n199), .A2(inst2_n2785), .B1(inst2_n2784),
        .B2(ciphertext2[24]), .ZN(inst2_n2220) );
  INV_X1 inst2_U373 ( .A(inst2_n2785), .ZN(inst2_n2784) );
  OAI211_X1 inst2_U372 ( .C1(inst2_n2219), .C2(inst2_n2794), .A(inst2_n2218),
        .B(inst2_n2217), .ZN(inst2_stateArray_S23reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst2_U371 ( .B1(inst2_n2791), .B2(ciphertext2[53]), .A(inst2_n2216), .ZN(inst2_n2217) );
  OAI22_X1 inst2_U370 ( .A1(inst2_n2463), .A2(inst2_n2804), .B1(inst2_n2396),
        .B2(inst2_n2820), .ZN(inst2_n2216) );
  AOI22_X1 inst2_U369 ( .A1(done2), .A2(ciphertext2[37]), .B1(plaintext2[37]),
        .B2(inst2_n2803), .ZN(inst2_n2218) );
  XNOR2_X1 inst2_U368 ( .A(inst2_n2215), .B(inst2_n2214), .ZN(inst2_n2219) );
  AOI22_X1 inst2_U367 ( .A1(inst2_n2261), .A2(ciphertext2[28]), .B1(inst2_n207), .B2(inst2_n2260), .ZN(inst2_n2214) );
  INV_X1 inst2_U366 ( .A(inst2_n2261), .ZN(inst2_n2260) );
  AOI22_X1 inst2_U365 ( .A1(ciphertext2[60]), .A2(inst2_n190), .B1(
        ciphertext2[93]), .B2(inst2_n2809), .ZN(inst2_n2215) );
  OAI211_X1 inst2_U364 ( .C1(inst2_n2213), .C2(inst2_n2780), .A(inst2_n2212),
        .B(inst2_n2211), .ZN(inst2_stateArray_S23reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst2_U363 ( .B1(inst2_n2791), .B2(ciphertext2[54]), .A(inst2_n2210), .ZN(inst2_n2211) );
  OAI22_X1 inst2_U362 ( .A1(inst2_n215), .A2(inst2_n2463), .B1(inst2_n2396),
        .B2(inst2_n2807), .ZN(inst2_n2210) );
  AOI22_X1 inst2_U361 ( .A1(inst2_n2788), .A2(ciphertext2[38]), .B1(
        plaintext2[38]), .B2(inst2_n2803), .ZN(inst2_n2212) );
  INV_X1 inst2_U360 ( .A(inst2_n2711), .ZN(inst2_n2788) );
  XNOR2_X1 inst2_U359 ( .A(inst2_n2209), .B(inst2_n2208), .ZN(inst2_n2213) );
  AOI22_X1 inst2_U358 ( .A1(inst2_n206), .A2(inst2_n2804), .B1(ciphertext2[29]), .B2(ciphertext2[94]), .ZN(inst2_n2208) );
  AOI22_X1 inst2_U357 ( .A1(inst2_n2254), .A2(ciphertext2[61]), .B1(
        inst2_n2820), .B2(inst2_n2255), .ZN(inst2_n2209) );
  INV_X1 inst2_U356 ( .A(inst2_n2254), .ZN(inst2_n2255) );
  OAI211_X1 inst2_U355 ( .C1(inst2_n2207), .C2(inst2_n2794), .A(inst2_n2206),
        .B(inst2_n2205), .ZN(inst2_stateArray_S23reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst2_U354 ( .B1(inst2_n2791), .B2(ciphertext2[55]), .A(inst2_n2204), .ZN(inst2_n2205) );
  OAI22_X1 inst2_U353 ( .A1(inst2_n219), .A2(inst2_n2789), .B1(inst2_n2463),
        .B2(inst2_n2805), .ZN(inst2_n2204) );
  AOI22_X1 inst2_U352 ( .A1(done2), .A2(ciphertext2[39]), .B1(plaintext2[39]),
        .B2(inst2_n2803), .ZN(inst2_n2206) );
  XNOR2_X1 inst2_U351 ( .A(inst2_n2203), .B(inst2_n2202), .ZN(inst2_n2207) );
  AOI22_X1 inst2_U350 ( .A1(inst2_n215), .A2(inst2_n2807), .B1(ciphertext2[62]), .B2(ciphertext2[30]), .ZN(inst2_n2202) );
  AOI22_X1 inst2_U349 ( .A1(ciphertext2[31]), .A2(inst2_n2390), .B1(
        inst2_n2389), .B2(inst2_n2805), .ZN(inst2_n2203) );
  INV_X1 inst2_U348 ( .A(inst2_n2390), .ZN(inst2_n2389) );
  OAI211_X1 inst2_U347 ( .C1(inst2_n2201), .C2(inst2_n2780), .A(inst2_n2200),
        .B(inst2_n2199), .ZN(inst2_stateArray_S23reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst2_U346 ( .B1(inst2_n2791), .B2(ciphertext2[51]), .A(inst2_n2198), .ZN(inst2_n2199) );
  OAI22_X1 inst2_U345 ( .A1(inst2_n196), .A2(inst2_n2789), .B1(inst2_n2463),
        .B2(inst2_n2806), .ZN(inst2_n2198) );
  AOI22_X1 inst2_U344 ( .A1(done2), .A2(ciphertext2[35]), .B1(plaintext2[35]),
        .B2(inst2_n2803), .ZN(inst2_n2200) );
  XNOR2_X1 inst2_U343 ( .A(inst2_n2197), .B(inst2_n2196), .ZN(inst2_n2201) );
  AOI22_X1 inst2_U342 ( .A1(ciphertext2[27]), .A2(inst2_n2310), .B1(
        inst2_n2309), .B2(inst2_n2806), .ZN(inst2_n2196) );
  INV_X1 inst2_U341 ( .A(inst2_n2310), .ZN(inst2_n2309) );
  XNOR2_X1 inst2_U340 ( .A(inst2_n2785), .B(inst2_n2195), .ZN(inst2_n2197) );
  AOI22_X1 inst2_U339 ( .A1(inst2_n203), .A2(inst2_n193), .B1(ciphertext2[58]),
        .B2(ciphertext2[26]), .ZN(inst2_n2195) );
  AOI22_X1 inst2_U338 ( .A1(ciphertext2[31]), .A2(inst2_n219), .B1(
        ciphertext2[63]), .B2(inst2_n2805), .ZN(inst2_n2785) );
  NAND2_X1 inst2_U337 ( .A1(inst2_n2194), .A2(inst2_n2193), .ZN(
        inst2_stateArray_S33reg_gff_1_SFF_0_n5) );
  AOI22_X1 inst2_U336 ( .A1(inst2_n2192), .A2(inst2_n2191), .B1(inst2_n2190),
        .B2(inst2_n2189), .ZN(inst2_n2193) );
  AOI211_X1 inst2_U335 ( .C1(plaintext2[0]), .C2(inst2_n2803), .A(inst2_n2188),
        .B(inst2_n2187), .ZN(inst2_n2194) );
  OAI22_X1 inst2_U334 ( .A1(inst2_n2186), .A2(inst2_n2780), .B1(inst2_n1201),
        .B2(inst2_n2711), .ZN(inst2_n2187) );
  XNOR2_X1 inst2_U333 ( .A(inst2_n2345), .B(inst2_n2185), .ZN(inst2_n2186) );
  AOI22_X1 inst2_U332 ( .A1(inst2_n2184), .A2(inst2_n2808), .B1(
        ciphertext2[56]), .B2(inst2_n2183), .ZN(inst2_n2185) );
  AOI22_X1 inst2_U331 ( .A1(inst2_n210), .A2(inst2_n209), .B1(ciphertext2[88]),
        .B2(ciphertext2[120]), .ZN(inst2_n2345) );
  OAI22_X1 inst2_U330 ( .A1(inst2_n199), .A2(inst2_n2789), .B1(inst2_n1209),
        .B2(inst2_n2757), .ZN(inst2_n2188) );
  NAND2_X1 inst2_U329 ( .A1(inst2_n2182), .A2(inst2_n2181), .ZN(
        inst2_stateArray_S33reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst2_U328 ( .A1(inst2_n2180), .A2(inst2_n2191), .B1(inst2_n2190),
        .B2(inst2_n2179), .ZN(inst2_n2181) );
  AOI211_X1 inst2_U327 ( .C1(plaintext2[1]), .C2(inst2_n2803), .A(inst2_n2178),
        .B(inst2_n2177), .ZN(inst2_n2182) );
  OAI22_X1 inst2_U326 ( .A1(inst2_n2176), .A2(inst2_n2780), .B1(inst2_n1200),
        .B2(inst2_n2711), .ZN(inst2_n2177) );
  XNOR2_X1 inst2_U325 ( .A(inst2_n2175), .B(inst2_n2174), .ZN(inst2_n2176) );
  AOI22_X1 inst2_U324 ( .A1(inst2_n210), .A2(inst2_n2184), .B1(inst2_n2183),
        .B2(ciphertext2[120]), .ZN(inst2_n2174) );
  XNOR2_X1 inst2_U323 ( .A(inst2_n2783), .B(inst2_n2173), .ZN(inst2_n2175) );
  AOI22_X1 inst2_U322 ( .A1(inst2_n199), .A2(ciphertext2[57]), .B1(inst2_n2810), .B2(ciphertext2[24]), .ZN(inst2_n2173) );
  AOI22_X1 inst2_U321 ( .A1(inst2_n198), .A2(inst2_n197), .B1(ciphertext2[89]),
        .B2(ciphertext2[121]), .ZN(inst2_n2783) );
  OAI22_X1 inst2_U320 ( .A1(inst2_n191), .A2(inst2_n2789), .B1(inst2_n1208),
        .B2(inst2_n2757), .ZN(inst2_n2178) );
  NAND2_X1 inst2_U319 ( .A1(inst2_n2172), .A2(inst2_n2171), .ZN(
        inst2_stateArray_S33reg_gff_1_SFF_2_n5) );
  AOI22_X1 inst2_U318 ( .A1(inst2_n2170), .A2(inst2_n2190), .B1(inst2_n2191),
        .B2(inst2_n2169), .ZN(inst2_n2171) );
  AOI211_X1 inst2_U317 ( .C1(plaintext2[2]), .C2(inst2_n2803), .A(inst2_n2168),
        .B(inst2_n2167), .ZN(inst2_n2172) );
  OAI22_X1 inst2_U316 ( .A1(inst2_n1199), .A2(inst2_n2711), .B1(inst2_n2780),
        .B2(inst2_n2166), .ZN(inst2_n2167) );
  XNOR2_X1 inst2_U315 ( .A(inst2_n2165), .B(inst2_n2164), .ZN(inst2_n2166) );
  AOI22_X1 inst2_U314 ( .A1(inst2_n198), .A2(ciphertext2[58]), .B1(inst2_n193),
        .B2(ciphertext2[121]), .ZN(inst2_n2164) );
  XNOR2_X1 inst2_U313 ( .A(inst2_n191), .B(inst2_n2775), .ZN(inst2_n2165) );
  AOI22_X1 inst2_U312 ( .A1(ciphertext2[122]), .A2(inst2_n194), .B1(
        ciphertext2[90]), .B2(inst2_n2800), .ZN(inst2_n2775) );
  OAI22_X1 inst2_U311 ( .A1(inst2_n203), .A2(inst2_n2789), .B1(inst2_n1207),
        .B2(inst2_n2757), .ZN(inst2_n2168) );
  NAND2_X1 inst2_U310 ( .A1(inst2_n2163), .A2(inst2_n2162), .ZN(
        inst2_stateArray_S33reg_gff_1_SFF_3_n5) );
  AOI22_X1 inst2_U309 ( .A1(inst2_n2161), .A2(inst2_n2191), .B1(inst2_n2160),
        .B2(inst2_n2190), .ZN(inst2_n2162) );
  AOI211_X1 inst2_U308 ( .C1(plaintext2[3]), .C2(inst2_n2803), .A(inst2_n2159),
        .B(inst2_n2158), .ZN(inst2_n2163) );
  OAI22_X1 inst2_U307 ( .A1(inst2_n2157), .A2(inst2_n2780), .B1(inst2_n1198),
        .B2(inst2_n2711), .ZN(inst2_n2158) );
  XNOR2_X1 inst2_U306 ( .A(inst2_n2156), .B(inst2_n2155), .ZN(inst2_n2157) );
  AOI22_X1 inst2_U305 ( .A1(inst2_n2184), .A2(inst2_n196), .B1(ciphertext2[59]), .B2(inst2_n2183), .ZN(inst2_n2155) );
  INV_X1 inst2_U304 ( .A(inst2_n2184), .ZN(inst2_n2183) );
  XNOR2_X1 inst2_U303 ( .A(inst2_n2310), .B(inst2_n2277), .ZN(inst2_n2156) );
  AOI22_X1 inst2_U302 ( .A1(ciphertext2[122]), .A2(inst2_n203), .B1(
        ciphertext2[26]), .B2(inst2_n2800), .ZN(inst2_n2277) );
  AOI22_X1 inst2_U301 ( .A1(inst2_n202), .A2(inst2_n201), .B1(ciphertext2[91]),
        .B2(ciphertext2[123]), .ZN(inst2_n2310) );
  OAI22_X1 inst2_U300 ( .A1(inst2_n1206), .A2(inst2_n2760), .B1(inst2_n2789),
        .B2(inst2_n2806), .ZN(inst2_n2159) );
  NAND2_X1 inst2_U299 ( .A1(inst2_n2154), .A2(inst2_n2153), .ZN(
        inst2_stateArray_S33reg_gff_1_SFF_4_n5) );
  AOI22_X1 inst2_U298 ( .A1(inst2_n2190), .A2(inst2_n2152), .B1(inst2_n2191),
        .B2(inst2_n2151), .ZN(inst2_n2153) );
  AOI211_X1 inst2_U297 ( .C1(plaintext2[4]), .C2(inst2_n2803), .A(inst2_n2150),
        .B(inst2_n2149), .ZN(inst2_n2154) );
  OAI22_X1 inst2_U296 ( .A1(inst2_n2148), .A2(inst2_n2780), .B1(inst2_n1197),
        .B2(inst2_n2711), .ZN(inst2_n2149) );
  XNOR2_X1 inst2_U295 ( .A(inst2_n2147), .B(inst2_n2146), .ZN(inst2_n2148) );
  XNOR2_X1 inst2_U294 ( .A(inst2_n202), .B(inst2_n2311), .ZN(inst2_n2146) );
  AOI22_X1 inst2_U293 ( .A1(inst2_n212), .A2(ciphertext2[60]), .B1(inst2_n2809), .B2(ciphertext2[92]), .ZN(inst2_n2311) );
  XOR2_X1 inst2_U292 ( .A(inst2_n2145), .B(inst2_n2184), .Z(inst2_n2147) );
  AOI22_X1 inst2_U291 ( .A1(inst2_n218), .A2(ciphertext2[31]), .B1(inst2_n2805), .B2(ciphertext2[127]), .ZN(inst2_n2184) );
  AOI22_X1 inst2_U290 ( .A1(ciphertext2[124]), .A2(ciphertext2[27]), .B1(
        inst2_n2806), .B2(inst2_n2799), .ZN(inst2_n2145) );
  OAI22_X1 inst2_U289 ( .A1(inst2_n207), .A2(inst2_n2789), .B1(inst2_n1205),
        .B2(inst2_n2757), .ZN(inst2_n2150) );
  NAND2_X1 inst2_U288 ( .A1(inst2_n2144), .A2(inst2_n2143), .ZN(
        inst2_stateArray_S33reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst2_U287 ( .A1(inst2_n2142), .A2(inst2_n2191), .B1(inst2_n2190),
        .B2(inst2_n2141), .ZN(inst2_n2143) );
  AOI211_X1 inst2_U286 ( .C1(plaintext2[5]), .C2(inst2_n2803), .A(inst2_n2140),
        .B(inst2_n2139), .ZN(inst2_n2144) );
  OAI22_X1 inst2_U285 ( .A1(inst2_n2138), .A2(inst2_n2780), .B1(inst2_n1196),
        .B2(inst2_n2711), .ZN(inst2_n2139) );
  XNOR2_X1 inst2_U284 ( .A(inst2_n2137), .B(inst2_n2319), .ZN(inst2_n2138) );
  AOI22_X1 inst2_U283 ( .A1(ciphertext2[61]), .A2(inst2_n190), .B1(
        ciphertext2[93]), .B2(inst2_n2820), .ZN(inst2_n2319) );
  XNOR2_X1 inst2_U282 ( .A(inst2_n214), .B(inst2_n2764), .ZN(inst2_n2137) );
  AOI22_X1 inst2_U281 ( .A1(ciphertext2[124]), .A2(inst2_n207), .B1(
        ciphertext2[28]), .B2(inst2_n2799), .ZN(inst2_n2764) );
  OAI22_X1 inst2_U280 ( .A1(inst2_n1204), .A2(inst2_n2760), .B1(inst2_n2396),
        .B2(inst2_n2804), .ZN(inst2_n2140) );
  NAND2_X1 inst2_U279 ( .A1(inst2_n2136), .A2(inst2_n2135), .ZN(
        inst2_stateArray_S33reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst2_U278 ( .A1(inst2_n2134), .A2(inst2_n2191), .B1(inst2_n2190),
        .B2(inst2_n2133), .ZN(inst2_n2135) );
  AOI211_X1 inst2_U277 ( .C1(plaintext2[6]), .C2(inst2_n2803), .A(inst2_n2132),
        .B(inst2_n2131), .ZN(inst2_n2136) );
  OAI22_X1 inst2_U276 ( .A1(inst2_n2130), .A2(inst2_n2780), .B1(inst2_n1195),
        .B2(inst2_n2711), .ZN(inst2_n2131) );
  XNOR2_X1 inst2_U275 ( .A(inst2_n2129), .B(inst2_n2261), .ZN(inst2_n2130) );
  AOI22_X1 inst2_U274 ( .A1(inst2_n214), .A2(ciphertext2[29]), .B1(inst2_n2804), .B2(ciphertext2[125]), .ZN(inst2_n2261) );
  XNOR2_X1 inst2_U273 ( .A(inst2_n216), .B(inst2_n2332), .ZN(inst2_n2129) );
  AOI22_X1 inst2_U272 ( .A1(ciphertext2[62]), .A2(inst2_n206), .B1(
        ciphertext2[94]), .B2(inst2_n2807), .ZN(inst2_n2332) );
  OAI22_X1 inst2_U271 ( .A1(inst2_n215), .A2(inst2_n2789), .B1(inst2_n1203),
        .B2(inst2_n2757), .ZN(inst2_n2132) );
  INV_X1 inst2_U270 ( .A(inst2_n2791), .ZN(inst2_n2757) );
  OAI211_X1 inst2_U269 ( .C1(inst2_n2128), .C2(inst2_n2127), .A(inst2_n2126),
        .B(inst2_n2125), .ZN(inst2_stateArray_S33reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst2_U268 ( .A1(inst2_n2124), .A2(inst2_n2191), .ZN(inst2_n2125)
         );
  NOR2_X1 inst2_U267 ( .A1(inst2_n2463), .A2(inst2_n2123), .ZN(inst2_n2191) );
  INV_X1 inst2_U266 ( .A(inst2_n2122), .ZN(inst2_n2463) );
  INV_X1 inst2_U265 ( .A(inst2_n2670), .ZN(inst2_n2122) );
  AOI211_X1 inst2_U264 ( .C1(plaintext2[7]), .C2(inst2_n2803), .A(inst2_n2121),
        .B(inst2_n2120), .ZN(inst2_n2126) );
  OAI22_X1 inst2_U263 ( .A1(inst2_n2119), .A2(inst2_n2780), .B1(inst2_n1194),
        .B2(inst2_n2711), .ZN(inst2_n2120) );
  INV_X1 inst2_U262 ( .A(inst2_n2393), .ZN(inst2_n2780) );
  INV_X1 inst2_U261 ( .A(inst2_n2794), .ZN(inst2_n2393) );
  NAND2_X1 inst2_U260 ( .A1(inst2_n2667), .A2(inst2_n2123), .ZN(inst2_n2794)
         );
  INV_X1 inst2_U259 ( .A(inst2_n2118), .ZN(inst2_n2123) );
  XNOR2_X1 inst2_U258 ( .A(inst2_n2117), .B(inst2_n2254), .ZN(inst2_n2119) );
  AOI22_X1 inst2_U257 ( .A1(inst2_n216), .A2(inst2_n215), .B1(ciphertext2[30]),
        .B2(ciphertext2[126]), .ZN(inst2_n2254) );
  XNOR2_X1 inst2_U256 ( .A(inst2_n219), .B(inst2_n2390), .ZN(inst2_n2117) );
  AOI22_X1 inst2_U255 ( .A1(inst2_n218), .A2(inst2_n220), .B1(ciphertext2[95]),
        .B2(ciphertext2[127]), .ZN(inst2_n2390) );
  OAI22_X1 inst2_U254 ( .A1(inst2_n1202), .A2(inst2_n2760), .B1(inst2_n2789),
        .B2(inst2_n2805), .ZN(inst2_n2121) );
  INV_X1 inst2_U253 ( .A(inst2_n2116), .ZN(inst2_n2789) );
  INV_X1 inst2_U252 ( .A(inst2_n2396), .ZN(inst2_n2116) );
  NAND2_X1 inst2_U251 ( .A1(inst2_n2667), .A2(inst2_n2118), .ZN(inst2_n2396)
         );
  INV_X1 inst2_U250 ( .A(inst2_n2791), .ZN(inst2_n2760) );
  AND2_X2 inst2_U249 ( .A1(inst2_n2872), .A2(inst2_n2711), .ZN(inst2_n2791) );
  INV_X1 inst2_U248 ( .A(inst2_n2190), .ZN(inst2_n2127) );
  NOR2_X1 inst2_U247 ( .A1(inst2_n2118), .A2(inst2_n2463), .ZN(inst2_n2190) );
  OAI211_X1 inst2_U246 ( .C1(inst2_n2854), .C2(inst2_n2565), .A(inst2_n2114),
        .B(inst2_n2113), .ZN(inst2_KeyArray_S30reg_gff_1_SFF_3_n6) );
  OAI21_X1 inst2_U245 ( .B1(inst2_n224), .B2(inst2_n2112), .A(inst2_n2111),
        .ZN(inst2_n2113) );
  AOI21_X1 inst2_U244 ( .B1(inst2_n224), .B2(inst2_n2112), .A(inst2_n2652),
        .ZN(inst2_n2111) );
  XNOR2_X1 inst2_U243 ( .A(inst2_n2160), .B(inst2_n2110), .ZN(inst2_n2112) );
  NOR2_X1 inst2_U242 ( .A1(inst2_n321), .A2(inst2_n706), .ZN(inst2_n2110) );
  XNOR2_X1 inst2_U241 ( .A(inst2_n2109), .B(inst2_n2108), .ZN(inst2_n2160) );
  XNOR2_X1 inst2_U240 ( .A(inst2_n2107), .B(inst2_n2106), .ZN(inst2_n2109) );
  AOI22_X1 inst2_U239 ( .A1(inst2_n71), .A2(inst2_n2375), .B1(key2[27]), .B2(
        inst2_n2803), .ZN(inst2_n2114) );
  OAI211_X1 inst2_U238 ( .C1(inst2_n2853), .C2(inst2_n2796), .A(inst2_n2105),
        .B(inst2_n2104), .ZN(inst2_KeyArray_S30reg_gff_1_SFF_6_n6) );
  OAI21_X1 inst2_U237 ( .B1(inst2_n222), .B2(inst2_n2103), .A(inst2_n2102),
        .ZN(inst2_n2104) );
  AOI21_X1 inst2_U236 ( .B1(inst2_n222), .B2(inst2_n2103), .A(inst2_n2652),
        .ZN(inst2_n2102) );
  XNOR2_X1 inst2_U235 ( .A(inst2_n2101), .B(inst2_n2133), .ZN(inst2_n2103) );
  XNOR2_X1 inst2_U234 ( .A(inst2_n2100), .B(inst2_n2099), .ZN(inst2_n2133) );
  NOR2_X1 inst2_U233 ( .A1(inst2_n718), .A2(inst2_n321), .ZN(inst2_n2101) );
  AOI22_X1 inst2_U232 ( .A1(inst2_n68), .A2(inst2_n2122), .B1(key2[30]), .B2(
        inst2_n2803), .ZN(inst2_n2105) );
  OAI211_X1 inst2_U231 ( .C1(inst2_n2852), .C2(inst2_n2565), .A(inst2_n2097),
        .B(inst2_n2096), .ZN(inst2_KeyArray_S30reg_gff_1_SFF_1_n6) );
  OAI21_X1 inst2_U230 ( .B1(inst2_n226), .B2(inst2_n2095), .A(inst2_n2094),
        .ZN(inst2_n2096) );
  AOI21_X1 inst2_U229 ( .B1(inst2_n226), .B2(inst2_n2095), .A(inst2_n2652),
        .ZN(inst2_n2094) );
  XNOR2_X1 inst2_U228 ( .A(inst2_n2093), .B(inst2_n2179), .ZN(inst2_n2095) );
  XNOR2_X1 inst2_U227 ( .A(inst2_n2092), .B(inst2_n2091), .ZN(inst2_n2179) );
  XNOR2_X1 inst2_U226 ( .A(inst2_n2108), .B(inst2_n2090), .ZN(inst2_n2092) );
  XNOR2_X1 inst2_U225 ( .A(inst2_n2089), .B(inst2_n2088), .ZN(inst2_n2090) );
  XOR2_X1 inst2_U224 ( .A(inst2_n2087), .B(inst2_n2086), .Z(inst2_n2088) );
  XNOR2_X1 inst2_U223 ( .A(inst2_n2085), .B(inst2_n2084), .ZN(inst2_n2108) );
  NOR2_X1 inst2_U222 ( .A1(inst2_n499), .A2(inst2_n321), .ZN(inst2_n2093) );
  AOI22_X1 inst2_U221 ( .A1(inst2_n73), .A2(inst2_n2568), .B1(key2[25]), .B2(
        inst2_n2803), .ZN(inst2_n2097) );
  OAI211_X1 inst2_U220 ( .C1(inst2_n2851), .C2(inst2_n2565), .A(inst2_n2083),
        .B(inst2_n2082), .ZN(inst2_KeyArray_S30reg_gff_1_SFF_2_n6) );
  OAI21_X1 inst2_U219 ( .B1(inst2_n225), .B2(inst2_n2081), .A(inst2_n2080),
        .ZN(inst2_n2082) );
  AOI21_X1 inst2_U218 ( .B1(inst2_n225), .B2(inst2_n2081), .A(inst2_n2652),
        .ZN(inst2_n2080) );
  XNOR2_X1 inst2_U217 ( .A(inst2_n2079), .B(inst2_n2170), .ZN(inst2_n2081) );
  XNOR2_X1 inst2_U216 ( .A(inst2_n2078), .B(inst2_n2077), .ZN(inst2_n2170) );
  XNOR2_X1 inst2_U215 ( .A(inst2_n2091), .B(inst2_n2076), .ZN(inst2_n2077) );
  XNOR2_X1 inst2_U214 ( .A(inst2_n2075), .B(inst2_n2074), .ZN(inst2_n2078) );
  XOR2_X1 inst2_U213 ( .A(inst2_n2073), .B(inst2_n2072), .Z(inst2_n2074) );
  NOR2_X1 inst2_U212 ( .A1(inst2_n2071), .A2(inst2_n2070), .ZN(inst2_n2075) );
  AOI21_X1 inst2_U211 ( .B1(inst2_n2069), .B2(inst2_n2068), .A(inst2_n2067),
        .ZN(inst2_n2071) );
  NOR2_X1 inst2_U210 ( .A1(inst2_n581), .A2(inst2_n321), .ZN(inst2_n2079) );
  AOI22_X1 inst2_U209 ( .A1(inst2_n72), .A2(inst2_n2375), .B1(key2[26]), .B2(
        inst2_n2803), .ZN(inst2_n2083) );
  OAI211_X1 inst2_U208 ( .C1(inst2_n2828), .C2(inst2_n2670), .A(inst2_n2066),
        .B(inst2_n2065), .ZN(inst2_KeyArray_S30reg_gff_1_SFF_4_n6) );
  OAI21_X1 inst2_U207 ( .B1(inst2_n223), .B2(inst2_n2064), .A(inst2_n2063),
        .ZN(inst2_n2065) );
  AOI21_X1 inst2_U206 ( .B1(inst2_n223), .B2(inst2_n2064), .A(inst2_n2652),
        .ZN(inst2_n2063) );
  XNOR2_X1 inst2_U205 ( .A(inst2_n2062), .B(inst2_n2152), .ZN(inst2_n2064) );
  XNOR2_X1 inst2_U204 ( .A(inst2_n2073), .B(inst2_n2100), .ZN(inst2_n2152) );
  XNOR2_X1 inst2_U203 ( .A(inst2_n2061), .B(inst2_n2107), .ZN(inst2_n2100) );
  XNOR2_X1 inst2_U202 ( .A(inst2_n2060), .B(inst2_n2059), .ZN(inst2_n2107) );
  NAND2_X1 inst2_U201 ( .A1(inst2_n2058), .A2(inst2_n2057), .ZN(inst2_n2060)
         );
  NOR2_X1 inst2_U200 ( .A1(inst2_n321), .A2(inst2_n1081), .ZN(inst2_n2062) );
  AOI22_X1 inst2_U199 ( .A1(inst2_n78), .A2(inst2_n2872), .B1(key2[28]), .B2(
        inst2_n2803), .ZN(inst2_n2066) );
  OAI211_X1 inst2_U198 ( .C1(inst2_n2850), .C2(inst2_n2796), .A(inst2_n2056),
        .B(inst2_n2055), .ZN(inst2_KeyArray_S30reg_gff_1_SFF_7_n6) );
  OAI21_X1 inst2_U197 ( .B1(inst2_n2054), .B2(inst2_n2802), .A(inst2_n2053),
        .ZN(inst2_n2055) );
  AOI21_X1 inst2_U196 ( .B1(inst2_n2054), .B2(inst2_n2802), .A(inst2_n2652),
        .ZN(inst2_n2053) );
  XNOR2_X1 inst2_U195 ( .A(inst2_n2052), .B(inst2_n2128), .ZN(inst2_n2054) );
  XNOR2_X1 inst2_U194 ( .A(inst2_n2051), .B(inst2_n2099), .ZN(inst2_n2128) );
  XNOR2_X1 inst2_U193 ( .A(inst2_n2091), .B(inst2_n2050), .ZN(inst2_n2099) );
  OAI221_X1 inst2_U192 ( .B1(inst2_n2049), .B2(inst2_n2048), .C1(inst2_n2047),
        .C2(inst2_n2046), .A(inst2_n2045), .ZN(inst2_n2091) );
  INV_X1 inst2_U191 ( .A(inst2_n2046), .ZN(inst2_n2048) );
  XNOR2_X1 inst2_U190 ( .A(inst2_n2073), .B(inst2_n2059), .ZN(inst2_n2051) );
  XNOR2_X1 inst2_U189 ( .A(inst2_n2044), .B(inst2_n2072), .ZN(inst2_n2059) );
  XNOR2_X1 inst2_U188 ( .A(inst2_n2043), .B(inst2_n2042), .ZN(inst2_n2072) );
  NAND2_X1 inst2_U187 ( .A1(inst2_n2058), .A2(inst2_n2041), .ZN(inst2_n2043)
         );
  XNOR2_X1 inst2_U186 ( .A(inst2_n2040), .B(inst2_n2039), .ZN(inst2_n2058) );
  XNOR2_X1 inst2_U185 ( .A(inst2_n2038), .B(inst2_n2037), .ZN(inst2_n2040) );
  NAND2_X1 inst2_U184 ( .A1(inst2_n2036), .A2(inst2_n2035), .ZN(inst2_n2044)
         );
  XNOR2_X1 inst2_U183 ( .A(inst2_n2034), .B(inst2_n2084), .ZN(inst2_n2073) );
  NAND2_X1 inst2_U182 ( .A1(inst2_n2033), .A2(inst2_n2032), .ZN(inst2_n2084)
         );
  NOR2_X1 inst2_U181 ( .A1(inst2_n1071), .A2(inst2_n321), .ZN(inst2_n2052) );
  AOI22_X1 inst2_U180 ( .A1(inst2_n67), .A2(inst2_n2568), .B1(key2[31]), .B2(
        inst2_n2803), .ZN(inst2_n2056) );
  OAI211_X1 inst2_U179 ( .C1(inst2_n2849), .C2(inst2_n2647), .A(inst2_n2031),
        .B(inst2_n2030), .ZN(inst2_KeyArray_S30reg_gff_1_SFF_0_n6) );
  OAI21_X1 inst2_U178 ( .B1(inst2_n227), .B2(inst2_n2029), .A(inst2_n2028),
        .ZN(inst2_n2030) );
  AOI21_X1 inst2_U177 ( .B1(inst2_n227), .B2(inst2_n2029), .A(inst2_n2652),
        .ZN(inst2_n2028) );
  XNOR2_X1 inst2_U176 ( .A(inst2_n2027), .B(inst2_n2189), .ZN(inst2_n2029) );
  XNOR2_X1 inst2_U175 ( .A(inst2_n2034), .B(inst2_n2026), .ZN(inst2_n2189) );
  XNOR2_X1 inst2_U174 ( .A(inst2_n2025), .B(inst2_n2089), .ZN(inst2_n2026) );
  XOR2_X1 inst2_U173 ( .A(inst2_n2042), .B(inst2_n2024), .Z(inst2_n2089) );
  OAI211_X1 inst2_U172 ( .C1(inst2_n2023), .C2(inst2_n2022), .A(inst2_n2021),
        .B(inst2_n2032), .ZN(inst2_n2024) );
  MUX2_X1 inst2_U171 ( .A(inst2_n2020), .B(inst2_n2038), .S(inst2_n2019), .Z(
        inst2_n2032) );
  XOR2_X1 inst2_U170 ( .A(inst2_n2018), .B(inst2_n2017), .Z(inst2_n2042) );
  NAND2_X1 inst2_U169 ( .A1(inst2_n2045), .A2(inst2_n2016), .ZN(inst2_n2017)
         );
  XNOR2_X1 inst2_U168 ( .A(inst2_n2015), .B(inst2_n2014), .ZN(inst2_n2045) );
  XNOR2_X1 inst2_U167 ( .A(inst2_n2013), .B(inst2_n2012), .ZN(inst2_n2014) );
  XOR2_X1 inst2_U166 ( .A(inst2_n2011), .B(inst2_n2010), .Z(inst2_n2015) );
  XNOR2_X1 inst2_U165 ( .A(inst2_n2085), .B(inst2_n2009), .ZN(inst2_n2025) );
  NOR2_X1 inst2_U164 ( .A1(inst2_n2008), .A2(inst2_n2007), .ZN(inst2_n2085) );
  AND2_X1 inst2_U163 ( .A1(inst2_n2006), .A2(inst2_n2005), .ZN(inst2_n2034) );
  NOR2_X1 inst2_U162 ( .A1(inst2_n444), .A2(inst2_n321), .ZN(inst2_n2027) );
  AOI22_X1 inst2_U161 ( .A1(inst2_n74), .A2(inst2_n2375), .B1(key2[24]), .B2(
        inst2_n2484), .ZN(inst2_n2031) );
  OAI211_X1 inst2_U160 ( .C1(inst2_n2848), .C2(inst2_n2796), .A(inst2_n2004),
        .B(inst2_n2003), .ZN(inst2_KeyArray_S30reg_gff_1_SFF_5_n6) );
  OAI21_X1 inst2_U159 ( .B1(inst2_n228), .B2(inst2_n2002), .A(inst2_n2001),
        .ZN(inst2_n2003) );
  AOI21_X1 inst2_U158 ( .B1(inst2_n228), .B2(inst2_n2002), .A(inst2_n2652),
        .ZN(inst2_n2001) );
  INV_X4 inst2_U157 ( .A(inst2_n2115), .ZN(inst2_n2667) );
  INV_X1 inst2_U156 ( .A(inst2_n2098), .ZN(inst2_n2565) );
  XNOR2_X1 inst2_U155 ( .A(inst2_n1999), .B(inst2_n2141), .ZN(inst2_n2002) );
  XOR2_X1 inst2_U154 ( .A(inst2_n1998), .B(inst2_n2018), .Z(inst2_n2141) );
  NAND2_X1 inst2_U153 ( .A1(inst2_n1997), .A2(inst2_n1996), .ZN(inst2_n2018)
         );
  XNOR2_X1 inst2_U152 ( .A(inst2_n1995), .B(inst2_n1994), .ZN(inst2_n1998) );
  NAND2_X1 inst2_U151 ( .A1(inst2_n1993), .A2(inst2_n1992), .ZN(inst2_n1994)
         );
  XNOR2_X1 inst2_U150 ( .A(inst2_n2050), .B(inst2_n2076), .ZN(inst2_n1995) );
  XNOR2_X1 inst2_U149 ( .A(inst2_n1991), .B(inst2_n2009), .ZN(inst2_n2076) );
  XNOR2_X1 inst2_U148 ( .A(inst2_n1990), .B(inst2_n2087), .ZN(inst2_n2009) );
  NAND2_X1 inst2_U147 ( .A1(inst2_n1989), .A2(inst2_n2005), .ZN(inst2_n2087)
         );
  XOR2_X1 inst2_U146 ( .A(inst2_n1988), .B(inst2_n1987), .Z(inst2_n2005) );
  XOR2_X1 inst2_U145 ( .A(inst2_n1986), .B(inst2_n2020), .Z(inst2_n1988) );
  XOR2_X1 inst2_U144 ( .A(inst2_n2038), .B(inst2_n1985), .Z(inst2_n2020) );
  XNOR2_X1 inst2_U143 ( .A(inst2_n2061), .B(inst2_n2106), .ZN(inst2_n1990) );
  NOR2_X1 inst2_U142 ( .A1(inst2_n2069), .A2(inst2_n2070), .ZN(inst2_n2106) );
  XOR2_X1 inst2_U141 ( .A(inst2_n2010), .B(inst2_n1984), .Z(inst2_n2070) );
  AND2_X1 inst2_U140 ( .A1(inst2_n1983), .A2(inst2_n2036), .ZN(inst2_n2061) );
  AOI22_X1 inst2_U139 ( .A1(inst2_n1982), .A2(inst2_n1981), .B1(inst2_n2038),
        .B2(inst2_n1980), .ZN(inst2_n2036) );
  INV_X1 inst2_U138 ( .A(inst2_n1979), .ZN(inst2_n1980) );
  XNOR2_X1 inst2_U137 ( .A(inst2_n1978), .B(inst2_n2086), .ZN(inst2_n1991) );
  NAND2_X1 inst2_U136 ( .A1(inst2_n1977), .A2(inst2_n1992), .ZN(inst2_n2086)
         );
  XNOR2_X1 inst2_U135 ( .A(inst2_n1976), .B(inst2_n2011), .ZN(inst2_n1992) );
  XNOR2_X1 inst2_U134 ( .A(inst2_n1975), .B(inst2_n1985), .ZN(inst2_n2011) );
  NAND3_X1 inst2_U133 ( .A1(inst2_n1974), .A2(inst2_n1973), .A3(inst2_n1972),
        .ZN(inst2_n1985) );
  INV_X1 inst2_U132 ( .A(inst2_n1971), .ZN(inst2_n1974) );
  XNOR2_X1 inst2_U131 ( .A(inst2_n2039), .B(inst2_n1970), .ZN(inst2_n1975) );
  XNOR2_X1 inst2_U130 ( .A(inst2_n1969), .B(inst2_n2021), .ZN(inst2_n2039) );
  NOR2_X1 inst2_U129 ( .A1(inst2_n1981), .A2(inst2_n1982), .ZN(inst2_n1969) );
  NAND2_X1 inst2_U128 ( .A1(inst2_n1979), .A2(inst2_n1968), .ZN(inst2_n1982)
         );
  XNOR2_X1 inst2_U127 ( .A(inst2_n2067), .B(inst2_n1967), .ZN(inst2_n1976) );
  NOR2_X1 inst2_U126 ( .A1(inst2_n2007), .A2(inst2_n1966), .ZN(inst2_n1978) );
  XNOR2_X1 inst2_U125 ( .A(inst2_n2012), .B(inst2_n1965), .ZN(inst2_n2007) );
  NAND2_X1 inst2_U124 ( .A1(inst2_n1964), .A2(inst2_n1996), .ZN(inst2_n2050)
         );
  XNOR2_X1 inst2_U123 ( .A(inst2_n1963), .B(inst2_n1962), .ZN(inst2_n1996) );
  XOR2_X1 inst2_U122 ( .A(inst2_n1987), .B(inst2_n2010), .Z(inst2_n1962) );
  XOR2_X1 inst2_U121 ( .A(inst2_n1961), .B(inst2_n1960), .Z(inst2_n2010) );
  OAI211_X1 inst2_U120 ( .C1(inst2_n2038), .C2(inst2_n1968), .A(inst2_n1979),
        .B(inst2_n1959), .ZN(inst2_n1960) );
  NAND2_X1 inst2_U119 ( .A1(inst2_n2038), .A2(inst2_n1968), .ZN(inst2_n1959)
         );
  XNOR2_X1 inst2_U118 ( .A(inst2_n2037), .B(inst2_n2021), .ZN(inst2_n1979) );
  NAND2_X1 inst2_U117 ( .A1(inst2_n2023), .A2(inst2_n2022), .ZN(inst2_n2021)
         );
  XOR2_X1 inst2_U116 ( .A(inst2_n1958), .B(inst2_n1957), .Z(inst2_n2037) );
  XNOR2_X1 inst2_U115 ( .A(inst2_n1956), .B(inst2_n1955), .ZN(inst2_n1958) );
  XNOR2_X1 inst2_U114 ( .A(inst2_n1954), .B(inst2_n1965), .ZN(inst2_n1968) );
  XNOR2_X1 inst2_U113 ( .A(inst2_n1953), .B(inst2_n1952), .ZN(inst2_n1965) );
  XNOR2_X1 inst2_U112 ( .A(inst2_n2013), .B(inst2_n2067), .ZN(inst2_n1953) );
  XNOR2_X1 inst2_U111 ( .A(inst2_n1951), .B(inst2_n2012), .ZN(inst2_n1987) );
  XNOR2_X1 inst2_U110 ( .A(inst2_n1954), .B(inst2_n1950), .ZN(inst2_n2012) );
  AOI211_X1 inst2_U109 ( .C1(inst2_n1973), .C2(inst2_n2038), .A(inst2_n2019),
        .B(inst2_n1949), .ZN(inst2_n1950) );
  NOR2_X1 inst2_U108 ( .A1(inst2_n1973), .A2(inst2_n2038), .ZN(inst2_n1949) );
  INV_X1 inst2_U107 ( .A(inst2_n1972), .ZN(inst2_n2019) );
  XNOR2_X1 inst2_U106 ( .A(inst2_n2067), .B(inst2_n1948), .ZN(inst2_n1972) );
  XNOR2_X1 inst2_U105 ( .A(inst2_n1947), .B(inst2_n1946), .ZN(inst2_n1948) );
  NAND2_X1 inst2_U104 ( .A1(inst2_n1956), .A2(inst2_n1945), .ZN(inst2_n1946)
         );
  XOR2_X1 inst2_U103 ( .A(inst2_n1970), .B(inst2_n1955), .Z(inst2_n1947) );
  NOR2_X1 inst2_U102 ( .A1(inst2_n1981), .A2(inst2_n1971), .ZN(inst2_n2038) );
  XNOR2_X1 inst2_U101 ( .A(inst2_n1944), .B(inst2_n1954), .ZN(inst2_n1971) );
  XNOR2_X1 inst2_U100 ( .A(inst2_n1951), .B(inst2_n1986), .ZN(inst2_n1944) );
  XNOR2_X1 inst2_U99 ( .A(inst2_n1943), .B(inst2_n1942), .ZN(inst2_n1986) );
  INV_X1 inst2_U98 ( .A(inst2_n1941), .ZN(inst2_n1942) );
  XOR2_X1 inst2_U97 ( .A(inst2_n1970), .B(inst2_n1956), .Z(inst2_n1943) );
  NAND2_X1 inst2_U96 ( .A1(inst2_n2016), .A2(inst2_n1945), .ZN(inst2_n1956) );
  XOR2_X1 inst2_U95 ( .A(inst2_n1940), .B(inst2_n2046), .Z(inst2_n2016) );
  NAND2_X1 inst2_U94 ( .A1(inst2_n2041), .A2(inst2_n2057), .ZN(inst2_n1970) );
  XNOR2_X1 inst2_U93 ( .A(inst2_n2069), .B(inst2_n1983), .ZN(inst2_n2057) );
  XNOR2_X1 inst2_U92 ( .A(inst2_n1939), .B(inst2_n1938), .ZN(inst2_n2041) );
  XNOR2_X1 inst2_U91 ( .A(inst2_n2023), .B(inst2_n2049), .ZN(inst2_n1939) );
  INV_X1 inst2_U90 ( .A(inst2_n2047), .ZN(inst2_n2049) );
  XNOR2_X1 inst2_U89 ( .A(inst2_n1940), .B(inst2_n1945), .ZN(inst2_n2047) );
  XNOR2_X1 inst2_U88 ( .A(inst2_n1937), .B(inst2_n1936), .ZN(inst2_n1981) );
  XNOR2_X1 inst2_U87 ( .A(inst2_n1935), .B(inst2_n1934), .ZN(inst2_n1937) );
  NAND2_X1 inst2_U86 ( .A1(inst2_n2033), .A2(inst2_n2023), .ZN(inst2_n1934) );
  INV_X1 inst2_U85 ( .A(inst2_n2022), .ZN(inst2_n2033) );
  XOR2_X1 inst2_U84 ( .A(inst2_n2013), .B(inst2_n1933), .Z(inst2_n2022) );
  XNOR2_X1 inst2_U83 ( .A(inst2_n1961), .B(inst2_n1932), .ZN(inst2_n1935) );
  XOR2_X1 inst2_U82 ( .A(inst2_n1931), .B(inst2_n1930), .Z(inst2_n1932) );
  AOI21_X1 inst2_U81 ( .B1(inst2_n2046), .B2(inst2_n1945), .A(inst2_n1929),
        .ZN(inst2_n1930) );
  NOR2_X1 inst2_U80 ( .A1(inst2_n1940), .A2(inst2_n1945), .ZN(inst2_n1929) );
  XOR2_X1 inst2_U79 ( .A(inst2_n1961), .B(inst2_n1984), .Z(inst2_n1973) );
  XNOR2_X1 inst2_U78 ( .A(inst2_n1967), .B(inst2_n1952), .ZN(inst2_n1984) );
  XNOR2_X1 inst2_U77 ( .A(inst2_n1941), .B(inst2_n1955), .ZN(inst2_n1952) );
  NAND2_X1 inst2_U76 ( .A1(inst2_n1977), .A2(inst2_n1993), .ZN(inst2_n1955) );
  XOR2_X1 inst2_U75 ( .A(inst2_n1940), .B(inst2_n1951), .Z(inst2_n1993) );
  XNOR2_X1 inst2_U74 ( .A(inst2_n1928), .B(inst2_n1927), .ZN(inst2_n1977) );
  XOR2_X1 inst2_U73 ( .A(inst2_n1926), .B(inst2_n1945), .Z(inst2_n1928) );
  XNOR2_X1 inst2_U72 ( .A(inst2_n1925), .B(inst2_n1936), .ZN(inst2_n1941) );
  NAND2_X1 inst2_U71 ( .A1(inst2_n1997), .A2(inst2_n1964), .ZN(inst2_n1936) );
  AOI21_X1 inst2_U70 ( .B1(inst2_n1925), .B2(inst2_n1924), .A(inst2_n1923),
        .ZN(inst2_n1967) );
  NOR2_X1 inst2_U69 ( .A1(inst2_n1945), .A2(inst2_n1938), .ZN(inst2_n1923) );
  NAND2_X1 inst2_U68 ( .A1(inst2_n1945), .A2(inst2_n1938), .ZN(inst2_n1924) );
  NAND2_X1 inst2_U67 ( .A1(inst2_n2006), .A2(inst2_n1989), .ZN(inst2_n1961) );
  XOR2_X1 inst2_U66 ( .A(inst2_n2023), .B(inst2_n1951), .Z(inst2_n1989) );
  XOR2_X1 inst2_U65 ( .A(inst2_n2013), .B(inst2_n1925), .Z(inst2_n2006) );
  XNOR2_X1 inst2_U64 ( .A(inst2_n1922), .B(inst2_n1921), .ZN(inst2_n1954) );
  INV_X1 inst2_U63 ( .A(inst2_n1927), .ZN(inst2_n1921) );
  NAND2_X1 inst2_U62 ( .A1(inst2_n2035), .A2(inst2_n1983), .ZN(inst2_n1922) );
  XNOR2_X1 inst2_U61 ( .A(inst2_n1926), .B(inst2_n1920), .ZN(inst2_n1983) );
  INV_X1 inst2_U60 ( .A(inst2_n1997), .ZN(inst2_n1920) );
  XNOR2_X1 inst2_U59 ( .A(inst2_n1940), .B(inst2_n1919), .ZN(inst2_n2035) );
  XNOR2_X1 inst2_U58 ( .A(inst2_n2023), .B(inst2_n1997), .ZN(inst2_n1919) );
  XOR2_X1 inst2_U57 ( .A(inst2_n1951), .B(inst2_n2046), .Z(inst2_n1997) );
  NOR2_X1 inst2_U56 ( .A1(inst2_n2067), .A2(inst2_n1957), .ZN(inst2_n1963) );
  NOR2_X1 inst2_U55 ( .A1(inst2_n2008), .A2(inst2_n1966), .ZN(inst2_n1957) );
  XNOR2_X1 inst2_U54 ( .A(inst2_n1945), .B(inst2_n1938), .ZN(inst2_n1966) );
  XNOR2_X1 inst2_U53 ( .A(inst2_n2013), .B(inst2_n1951), .ZN(inst2_n1945) );
  AOI22_X1 inst2_U52 ( .A1(inst2_n2000), .A2(inst2_n9), .B1(inst2_n2124), .B2(
        inst2_n2797), .ZN(inst2_n1951) );
  AOI22_X1 inst2_U51 ( .A1(inst2_n221), .A2(inst2_n218), .B1(ciphertext2[127]),
        .B2(inst2_n2802), .ZN(inst2_n2124) );
  XNOR2_X1 inst2_U50 ( .A(inst2_n1925), .B(inst2_n1938), .ZN(inst2_n2008) );
  INV_X1 inst2_U49 ( .A(inst2_n1933), .ZN(inst2_n1938) );
  XOR2_X1 inst2_U48 ( .A(inst2_n2069), .B(inst2_n1918), .Z(inst2_n1933) );
  NOR2_X1 inst2_U47 ( .A1(inst2_n2069), .A2(inst2_n2068), .ZN(inst2_n2067) );
  XNOR2_X1 inst2_U46 ( .A(inst2_n2013), .B(inst2_n1927), .ZN(inst2_n2068) );
  XOR2_X1 inst2_U45 ( .A(inst2_n1918), .B(inst2_n2046), .Z(inst2_n1927) );
  AOI22_X1 inst2_U44 ( .A1(inst2_n2000), .A2(inst2_n11), .B1(inst2_n2151),
        .B2(inst2_n2797), .ZN(inst2_n2046) );
  AOI22_X1 inst2_U43 ( .A1(inst2_n223), .A2(inst2_n2799), .B1(ciphertext2[124]), .B2(inst2_n2817), .ZN(inst2_n2151) );
  AOI22_X1 inst2_U42 ( .A1(inst2_n2000), .A2(inst2_n10), .B1(inst2_n2142),
        .B2(inst2_n2797), .ZN(inst2_n2013) );
  AOI22_X1 inst2_U41 ( .A1(inst2_n228), .A2(inst2_n214), .B1(ciphertext2[125]),
        .B2(inst2_n2816), .ZN(inst2_n2142) );
  AOI22_X1 inst2_U40 ( .A1(inst2_n2000), .A2(inst2_n22), .B1(inst2_n2192),
        .B2(inst2_n2797), .ZN(inst2_n2069) );
  AOI22_X1 inst2_U39 ( .A1(inst2_n227), .A2(inst2_n210), .B1(ciphertext2[120]),
        .B2(inst2_n2819), .ZN(inst2_n2192) );
  XOR2_X1 inst2_U38 ( .A(inst2_n1925), .B(inst2_n1918), .Z(inst2_n1964) );
  AOI22_X1 inst2_U37 ( .A1(inst2_n2000), .A2(inst2_n24), .B1(inst2_n2134),
        .B2(inst2_n2797), .ZN(inst2_n1918) );
  AOI22_X1 inst2_U36 ( .A1(inst2_n222), .A2(inst2_n216), .B1(ciphertext2[126]),
        .B2(inst2_n2815), .ZN(inst2_n2134) );
  XOR2_X1 inst2_U35 ( .A(inst2_n1940), .B(inst2_n1926), .Z(inst2_n1925) );
  XOR2_X1 inst2_U34 ( .A(inst2_n2023), .B(inst2_n1931), .Z(inst2_n1926) );
  AOI22_X1 inst2_U33 ( .A1(inst2_n2000), .A2(inst2_n12), .B1(inst2_n2161),
        .B2(inst2_n2797), .ZN(inst2_n1931) );
  AOI22_X1 inst2_U32 ( .A1(inst2_n224), .A2(inst2_n202), .B1(ciphertext2[123]),
        .B2(inst2_n2818), .ZN(inst2_n2161) );
  AOI22_X1 inst2_U31 ( .A1(inst2_n2000), .A2(inst2_n17), .B1(inst2_n2180),
        .B2(inst2_n2797), .ZN(inst2_n2023) );
  AOI22_X1 inst2_U30 ( .A1(inst2_n198), .A2(inst2_n226), .B1(inst2_n2813),
        .B2(ciphertext2[121]), .ZN(inst2_n2180) );
  AOI22_X1 inst2_U29 ( .A1(inst2_n2000), .A2(inst2_n14), .B1(inst2_n2169),
        .B2(inst2_n2797), .ZN(inst2_n1940) );
  AOI22_X1 inst2_U28 ( .A1(ciphertext2[122]), .A2(inst2_n2814), .B1(inst2_n225), .B2(inst2_n2800), .ZN(inst2_n2169) );
  NOR2_X1 inst2_U27 ( .A1(inst2_n1080), .A2(inst2_n321), .ZN(inst2_n1999) );
  AOI22_X1 inst2_U26 ( .A1(inst2_n69), .A2(inst2_n2375), .B1(key2[29]), .B2(
        inst2_n2507), .ZN(inst2_n2004) );
  NAND2_X1 inst2_U25 ( .A1(inst2_n6), .A2(inst2_ctrl_n6), .ZN(inst2_n2797) );
  NAND2_X1 inst2_U24 ( .A1(inst2_n1917), .A2(inst2_n2826), .ZN(
        inst2_ctrl_seq4_SFF_0_n5) );
  INV_X1 inst2_U23 ( .A(inst2_n1915), .ZN(inst2_n1916) );
  OAI221_X1 inst2_U22 ( .B1(inst2_n232), .B2(inst2_n1290), .C1(inst2_n1914),
        .C2(done2), .A(inst2_n6), .ZN(inst2_ctrl_seq6_SFF_0_n5) );
  NAND2_X1 inst2_U21 ( .A1(inst2_n232), .A2(inst2_n1290), .ZN(inst2_n1914) );
  NAND2_X1 inst2_U20 ( .A1(inst2_n6), .A2(inst2_n231), .ZN(
        inst2_ctrl_seq6_SFF_4_n5) );
  NOR4_X2 inst2_U19 ( .A1(inst2_n1081), .A2(inst2_n499), .A3(inst2_n581), .A4(
        inst2_n1080), .ZN(inst2_n2118) );
  NAND4_X1 inst2_U18 ( .A1(inst2_n233), .A2(inst2_n232), .A3(inst2_n1290),
        .A4(inst2_n231), .ZN(inst2_n1915) );
  NAND2_X1 inst2_U17 ( .A1(inst2_n6), .A2(inst2_n230), .ZN(
        inst2_ctrl_seq6_SFF_2_n5) );
  INV_X1 inst2_U16 ( .A(reset2), .ZN(inst2_n1096) );
  INV_X1 inst2_U15 ( .A(inst2_n2666), .ZN(inst2_n2796) );
  NAND2_X1 inst2_U14 ( .A1(inst2_n1917), .A2(inst2_n2797), .ZN(inst2_n2670) );
  NOR2_X1 inst2_U13 ( .A1(inst2_ctrl_seq6_SFF_2_n5), .A2(inst2_n1915), .ZN(
        inst2_n2098) );
  INV_X1 inst2_U12 ( .A(inst2_n6), .ZN(inst2_n2582) );
  INV_X1 inst2_U11 ( .A(inst2_n2797), .ZN(inst2_n2000) );
  NAND2_X1 inst2_U10 ( .A1(inst2_n2000), .A2(inst2_n2565), .ZN(inst2_n2115) );
  AOI21_X4 inst2_U9 ( .B1(inst2_n230), .B2(inst2_n1916), .A(inst2_n2507), .ZN(
        inst2_n1917) );
  INV_X4 inst2_U8 ( .A(inst2_n1917), .ZN(inst2_n2771) );
  NAND4_X4 inst2_U7 ( .A1(inst2_n2872), .A2(inst2_n2118), .A3(inst2_n143),
        .A4(inst2_n236), .ZN(inst2_n2711) );
  INV_X2 inst2_U6 ( .A(inst2_n2711), .ZN(done2) );
  INV_X4 inst2_U5 ( .A(inst2_n2667), .ZN(inst2_n2652) );
  INV_X2 inst2_U4 ( .A(inst2_n2098), .ZN(inst2_n2647) );
  INV_X2 inst2_U3 ( .A(inst2_n2565), .ZN(inst2_n2872) );
  DFF_X2 inst2_nReset_reg_FF_FF ( .D(inst2_n1096), .CK(clk), .Q(inst2_n6),
        .QN(inst2_n2803) );
  DFF_X1 inst2_calcRCon_s_current_state_reg_7__FF_FF ( .D(inst2_calcRCon_n44),
        .CK(clk), .Q(inst2_n2801), .QN(inst2_n1071) );
  DFF_X1 inst2_calcRCon_s_current_state_reg_6__FF_FF ( .D(inst2_calcRCon_n45),
        .CK(clk), .QN(inst2_n718) );
  DFF_X1 inst2_calcRCon_s_current_state_reg_5__FF_FF ( .D(inst2_calcRCon_n46),
        .CK(clk), .QN(inst2_n1080) );
  DFF_X1 inst2_calcRCon_s_current_state_reg_4__FF_FF ( .D(inst2_calcRCon_n47),
        .CK(clk), .QN(inst2_n1081) );
  DFF_X1 inst2_calcRCon_s_current_state_reg_3__FF_FF ( .D(inst2_calcRCon_n48),
        .CK(clk), .Q(inst2_n2812), .QN(inst2_n706) );
  DFF_X1 inst2_calcRCon_s_current_state_reg_2__FF_FF ( .D(inst2_calcRCon_n49),
        .CK(clk), .Q(inst2_n2836), .QN(inst2_n581) );
  DFF_X1 inst2_calcRCon_s_current_state_reg_1__FF_FF ( .D(inst2_calcRCon_n50),
        .CK(clk), .QN(inst2_n499) );
  DFF_X1 inst2_calcRCon_s_current_state_reg_0__FF_FF ( .D(inst2_calcRCon_n51),
        .CK(clk), .Q(inst2_n2837), .QN(inst2_n444) );
  DFF_X1 inst2_KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S33reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst2_n1082) );
  DFF_X1 inst2_KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S33reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst2_n1083) );
  DFF_X1 inst2_KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S33reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst2_n1084) );
  DFF_X1 inst2_KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S33reg_gff_1_SFF_4_n5), .CK(clk), .QN(inst2_n1085) );
  DFF_X1 inst2_KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S33reg_gff_1_SFF_3_n5), .CK(clk), .QN(inst2_n1086) );
  DFF_X1 inst2_KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S33reg_gff_1_SFF_2_n5), .CK(clk), .QN(inst2_n1087) );
  DFF_X1 inst2_KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S33reg_gff_1_SFF_1_n5), .CK(clk), .Q(inst2_n57) );
  DFF_X1 inst2_KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S33reg_gff_1_SFF_0_n5), .CK(clk), .QN(inst2_n1089) );
  DFF_X1 inst2_KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S32reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst2_n1090) );
  DFF_X1 inst2_KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S32reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst2_n1091) );
  DFF_X1 inst2_KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S32reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst2_n1092) );
  DFF_X1 inst2_KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S32reg_gff_1_SFF_4_n6), .CK(clk), .QN(inst2_n1093) );
  DFF_X1 inst2_KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S32reg_gff_1_SFF_3_n6), .CK(clk), .QN(inst2_n1094) );
  DFF_X1 inst2_KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S32reg_gff_1_SFF_2_n6), .CK(clk), .QN(inst2_n1095) );
  DFF_X1 inst2_KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S32reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst2_n65) );
  DFF_X1 inst2_KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S32reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst2_n1097) );
  DFF_X1 inst2_KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S31reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst2_n67) );
  DFF_X1 inst2_KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S31reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst2_n68) );
  DFF_X1 inst2_KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S31reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst2_n69) );
  DFF_X1 inst2_KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S31reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst2_n70), .QN(
        inst2_n2828) );
  DFF_X1 inst2_KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S31reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst2_n71) );
  DFF_X1 inst2_KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S31reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst2_n72) );
  DFF_X1 inst2_KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S31reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst2_n73) );
  DFF_X1 inst2_KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S31reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst2_n74) );
  DFF_X1 inst2_KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S30reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst2_n75), .QN(
        inst2_n2850) );
  DFF_X1 inst2_KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S30reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst2_n76), .QN(
        inst2_n2853) );
  DFF_X1 inst2_KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S30reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst2_n77), .QN(
        inst2_n2848) );
  DFF_X1 inst2_KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S30reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst2_n78) );
  DFF_X1 inst2_KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S30reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst2_n79), .QN(
        inst2_n2854) );
  DFF_X1 inst2_KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S30reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst2_n80), .QN(
        inst2_n2851) );
  DFF_X1 inst2_KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S30reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst2_n81), .QN(
        inst2_n2852) );
  DFF_X1 inst2_KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S30reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst2_n82), .QN(
        inst2_n2849) );
  DFF_X1 inst2_KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S23reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst2_n83) );
  DFF_X1 inst2_KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S23reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst2_n84) );
  DFF_X1 inst2_KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S23reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst2_n85) );
  DFF_X1 inst2_KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S23reg_gff_1_SFF_4_n5), .CK(clk), .Q(inst2_n86) );
  DFF_X1 inst2_KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S23reg_gff_1_SFF_3_n5), .CK(clk), .Q(inst2_n87) );
  DFF_X1 inst2_KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S23reg_gff_1_SFF_2_n5), .CK(clk), .Q(inst2_n88) );
  DFF_X1 inst2_KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S23reg_gff_1_SFF_1_n5), .CK(clk), .Q(inst2_n89) );
  DFF_X1 inst2_KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S23reg_gff_1_SFF_0_n5), .CK(clk), .Q(inst2_n90) );
  DFF_X1 inst2_KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S22reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst2_n91) );
  DFF_X1 inst2_KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S22reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst2_n92) );
  DFF_X1 inst2_KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S22reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst2_n93) );
  DFF_X1 inst2_KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S22reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst2_n94) );
  DFF_X1 inst2_KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S22reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst2_n95) );
  DFF_X1 inst2_KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S22reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst2_n96) );
  DFF_X1 inst2_KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S22reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst2_n97) );
  DFF_X1 inst2_KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S22reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst2_n98) );
  DFF_X1 inst2_KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S21reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst2_n107) );
  DFF_X1 inst2_KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S21reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst2_n108) );
  DFF_X1 inst2_KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S21reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst2_n109) );
  DFF_X1 inst2_KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S21reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst2_n110) );
  DFF_X1 inst2_KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S21reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst2_n111) );
  DFF_X1 inst2_KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S21reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst2_n112) );
  DFF_X1 inst2_KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S21reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst2_n113) );
  DFF_X1 inst2_KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S21reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst2_n114) );
  DFF_X1 inst2_KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S20reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst2_n115) );
  DFF_X1 inst2_KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S20reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst2_n116) );
  DFF_X1 inst2_KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S20reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst2_n117) );
  DFF_X1 inst2_KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S20reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst2_n118) );
  DFF_X1 inst2_KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S20reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst2_n119) );
  DFF_X1 inst2_KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S20reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst2_n120) );
  DFF_X1 inst2_KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S20reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst2_n121) );
  DFF_X1 inst2_KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S20reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst2_n122), .QN(
        inst2_n2863) );
  DFF_X1 inst2_KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S13reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst2_n9), .QN(
        inst2_n2840) );
  DFF_X1 inst2_KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S13reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst2_n24), .QN(
        inst2_n2841) );
  DFF_X1 inst2_KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S13reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst2_n10), .QN(
        inst2_n2842) );
  DFF_X1 inst2_KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S13reg_gff_1_SFF_4_n5), .CK(clk), .Q(inst2_n11), .QN(
        inst2_n2843) );
  DFF_X1 inst2_KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S13reg_gff_1_SFF_3_n5), .CK(clk), .Q(inst2_n12), .QN(
        inst2_n2844) );
  DFF_X1 inst2_KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S13reg_gff_1_SFF_2_n5), .CK(clk), .Q(inst2_n14), .QN(
        inst2_n2845) );
  DFF_X1 inst2_KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S13reg_gff_1_SFF_1_n5), .CK(clk), .Q(inst2_n17), .QN(
        inst2_n2846) );
  DFF_X1 inst2_KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S13reg_gff_1_SFF_0_n5), .CK(clk), .Q(inst2_n22), .QN(
        inst2_n2847) );
  DFF_X1 inst2_KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S12reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst2_n123), .QN(
        inst2_n2864) );
  DFF_X1 inst2_KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S12reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst2_n124), .QN(
        inst2_n2865) );
  DFF_X1 inst2_KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S12reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst2_n125), .QN(
        inst2_n2866) );
  DFF_X1 inst2_KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S12reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst2_n126), .QN(
        inst2_n2867) );
  DFF_X1 inst2_KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S12reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst2_n127), .QN(
        inst2_n2868) );
  DFF_X1 inst2_KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S12reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst2_n128), .QN(
        inst2_n2869) );
  DFF_X1 inst2_KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S12reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst2_n129), .QN(
        inst2_n2870) );
  DFF_X1 inst2_KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S12reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst2_n130), .QN(
        inst2_n2871) );
  DFF_X1 inst2_KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S11reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst2_n131) );
  DFF_X1 inst2_KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S11reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst2_n132) );
  DFF_X1 inst2_KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S11reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst2_n133) );
  DFF_X1 inst2_KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S11reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst2_n134) );
  DFF_X1 inst2_KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S11reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst2_n135) );
  DFF_X1 inst2_KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S11reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst2_n136) );
  DFF_X1 inst2_KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S11reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst2_n137) );
  DFF_X1 inst2_KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S11reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst2_n1161) );
  DFF_X1 inst2_KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S10reg_gff_1_SFF_7_n6), .CK(clk), .QN(inst2_n1162) );
  DFF_X1 inst2_KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S10reg_gff_1_SFF_6_n6), .CK(clk), .QN(inst2_n1163) );
  DFF_X1 inst2_KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S10reg_gff_1_SFF_5_n6), .CK(clk), .QN(inst2_n1164) );
  DFF_X1 inst2_KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S10reg_gff_1_SFF_4_n6), .CK(clk), .QN(inst2_n1165) );
  DFF_X1 inst2_KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S10reg_gff_1_SFF_3_n6), .CK(clk), .QN(inst2_n1166) );
  DFF_X1 inst2_KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S10reg_gff_1_SFF_2_n6), .CK(clk), .QN(inst2_n1167) );
  DFF_X1 inst2_KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S10reg_gff_1_SFF_1_n6), .CK(clk), .QN(inst2_n1168) );
  DFF_X1 inst2_KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S10reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst2_n1169) );
  DFF_X1 inst2_KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S03reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst2_n1170) );
  DFF_X1 inst2_KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S03reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst2_n1171) );
  DFF_X1 inst2_KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S03reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst2_n1172) );
  DFF_X1 inst2_KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S03reg_gff_1_SFF_4_n5), .CK(clk), .QN(inst2_n1173) );
  DFF_X1 inst2_KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S03reg_gff_1_SFF_3_n5), .CK(clk), .QN(inst2_n1174) );
  DFF_X1 inst2_KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S03reg_gff_1_SFF_2_n5), .CK(clk), .QN(inst2_n1175) );
  DFF_X1 inst2_KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S03reg_gff_1_SFF_1_n5), .CK(clk), .QN(inst2_n1176) );
  DFF_X1 inst2_KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S03reg_gff_1_SFF_0_n5), .CK(clk), .QN(inst2_n1177) );
  DFF_X1 inst2_KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S02reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst2_n1178) );
  DFF_X1 inst2_KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S02reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst2_n1179) );
  DFF_X1 inst2_KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S02reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst2_n1180) );
  DFF_X1 inst2_KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S02reg_gff_1_SFF_4_n6), .CK(clk), .QN(inst2_n1181) );
  DFF_X1 inst2_KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S02reg_gff_1_SFF_3_n6), .CK(clk), .QN(inst2_n1182) );
  DFF_X1 inst2_KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S02reg_gff_1_SFF_2_n6), .CK(clk), .QN(inst2_n1183) );
  DFF_X1 inst2_KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S02reg_gff_1_SFF_1_n6), .CK(clk), .QN(inst2_n1184) );
  DFF_X1 inst2_KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S02reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst2_n1185) );
  DFF_X1 inst2_KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S01reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst2_n2821), .QN(
        inst2_n1186) );
  DFF_X1 inst2_KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S01reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst2_n2822), .QN(
        inst2_n1187) );
  DFF_X1 inst2_KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S01reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst2_n2823), .QN(
        inst2_n1188) );
  DFF_X1 inst2_KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S01reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst2_n2838), .QN(
        inst2_n1189) );
  DFF_X1 inst2_KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S01reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst2_n2824), .QN(
        inst2_n1190) );
  DFF_X1 inst2_KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S01reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst2_n2825), .QN(
        inst2_n1191) );
  DFF_X1 inst2_KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S01reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst2_n2839), .QN(
        inst2_n1192) );
  DFF_X1 inst2_KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S01reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst2_n1193) );
  DFF_X1 inst2_KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S00reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst2_n2802), .QN(
        inst2_n221) );
  DFF_X1 inst2_KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S00reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst2_n2815), .QN(
        inst2_n222) );
  DFF_X1 inst2_KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S00reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst2_n2816), .QN(
        inst2_n228) );
  DFF_X1 inst2_KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S00reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst2_n2817), .QN(
        inst2_n223) );
  DFF_X1 inst2_KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S00reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst2_n2818), .QN(
        inst2_n224) );
  DFF_X1 inst2_KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S00reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst2_n2814), .QN(
        inst2_n225) );
  DFF_X1 inst2_KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S00reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst2_n2813), .QN(
        inst2_n226) );
  DFF_X1 inst2_KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_KeyArray_S00reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst2_n2819), .QN(
        inst2_n227) );
  DFF_X1 inst2_stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S33reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext2[7]),
        .QN(inst2_n1194) );
  DFF_X1 inst2_stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S33reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext2[6]),
        .QN(inst2_n1195) );
  DFF_X1 inst2_stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S33reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext2[5]),
        .QN(inst2_n1196) );
  DFF_X1 inst2_stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S33reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext2[4]),
        .QN(inst2_n1197) );
  DFF_X1 inst2_stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S33reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext2[3]),
        .QN(inst2_n1198) );
  DFF_X1 inst2_stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S33reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext2[2]),
        .QN(inst2_n1199) );
  DFF_X1 inst2_stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S33reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext2[1]),
        .QN(inst2_n1200) );
  DFF_X1 inst2_stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S33reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext2[0]),
        .QN(inst2_n1201) );
  DFF_X1 inst2_stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S32reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext2[15]),
        .QN(inst2_n1202) );
  DFF_X1 inst2_stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S32reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext2[14]),
        .QN(inst2_n1203) );
  DFF_X1 inst2_stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S32reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext2[13]),
        .QN(inst2_n1204) );
  DFF_X1 inst2_stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S32reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[12]),
        .QN(inst2_n1205) );
  DFF_X1 inst2_stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S32reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[11]),
        .QN(inst2_n1206) );
  DFF_X1 inst2_stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S32reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[10]),
        .QN(inst2_n1207) );
  DFF_X1 inst2_stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S32reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[9]),
        .QN(inst2_n1208) );
  DFF_X1 inst2_stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S32reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[8]),
        .QN(inst2_n1209) );
  DFF_X1 inst2_stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S31reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext2[23]),
        .QN(inst2_n2829) );
  DFF_X1 inst2_stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S31reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext2[22]),
        .QN(inst2_n2827) );
  DFF_X1 inst2_stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S31reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext2[21]),
        .QN(inst2_n2830) );
  DFF_X1 inst2_stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S31reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[20]),
        .QN(inst2_n2831) );
  DFF_X1 inst2_stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S31reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[19]),
        .QN(inst2_n2832) );
  DFF_X1 inst2_stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S31reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[18]),
        .QN(inst2_n2833) );
  DFF_X1 inst2_stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S31reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[17]),
        .QN(inst2_n2834) );
  DFF_X1 inst2_stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S31reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[16]),
        .QN(inst2_n2835) );
  DFF_X1 inst2_stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S30reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext2[31]),
        .QN(inst2_n2805) );
  DFF_X1 inst2_stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S30reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext2[30]),
        .QN(inst2_n215) );
  DFF_X1 inst2_stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S30reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext2[29]),
        .QN(inst2_n2804) );
  DFF_X1 inst2_stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S30reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext2[28]),
        .QN(inst2_n207) );
  DFF_X1 inst2_stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S30reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext2[27]),
        .QN(inst2_n2806) );
  DFF_X1 inst2_stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S30reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext2[26]),
        .QN(inst2_n203) );
  DFF_X1 inst2_stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S30reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext2[25]),
        .QN(inst2_n191) );
  DFF_X1 inst2_stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S30reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext2[24]),
        .QN(inst2_n199) );
  DFF_X1 inst2_stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S23reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext2[39]),
        .QN(inst2_n1218) );
  DFF_X1 inst2_stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S23reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext2[38]),
        .QN(inst2_n1219) );
  DFF_X1 inst2_stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S23reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext2[37]),
        .QN(inst2_n1220) );
  DFF_X1 inst2_stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S23reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[36]),
        .QN(inst2_n1221) );
  DFF_X1 inst2_stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S23reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[35]),
        .QN(inst2_n1222) );
  DFF_X1 inst2_stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S23reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[34]),
        .QN(inst2_n1223) );
  DFF_X1 inst2_stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S23reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[33]),
        .QN(inst2_n1224) );
  DFF_X1 inst2_stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S23reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[32]),
        .QN(inst2_n1225) );
  DFF_X1 inst2_stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S22reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext2[47]),
        .QN(inst2_n1226) );
  DFF_X1 inst2_stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S22reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext2[46]),
        .QN(inst2_n1227) );
  DFF_X1 inst2_stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S22reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext2[45]),
        .QN(inst2_n1228) );
  DFF_X1 inst2_stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S22reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[44]),
        .QN(inst2_n1229) );
  DFF_X1 inst2_stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S22reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[43]),
        .QN(inst2_n1230) );
  DFF_X1 inst2_stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S22reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[42]),
        .QN(inst2_n1231) );
  DFF_X1 inst2_stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S22reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[41]),
        .QN(inst2_n1232) );
  DFF_X1 inst2_stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S22reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[40]),
        .QN(inst2_n1233) );
  DFF_X1 inst2_stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S21reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext2[55])
         );
  DFF_X1 inst2_stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S21reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext2[54])
         );
  DFF_X1 inst2_stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S21reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext2[53])
         );
  DFF_X1 inst2_stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S21reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[52])
         );
  DFF_X1 inst2_stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S21reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[51])
         );
  DFF_X1 inst2_stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S21reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[50])
         );
  DFF_X1 inst2_stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S21reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[49])
         );
  DFF_X1 inst2_stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S21reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[48])
         );
  DFF_X1 inst2_stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S20reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext2[63]),
        .QN(inst2_n219) );
  DFF_X1 inst2_stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S20reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext2[62]),
        .QN(inst2_n2807) );
  DFF_X1 inst2_stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S20reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext2[61]),
        .QN(inst2_n2820) );
  DFF_X1 inst2_stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S20reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext2[60]),
        .QN(inst2_n2809) );
  DFF_X1 inst2_stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S20reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext2[59]),
        .QN(inst2_n196) );
  DFF_X1 inst2_stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S20reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext2[58]),
        .QN(inst2_n193) );
  DFF_X1 inst2_stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S20reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext2[57]),
        .QN(inst2_n2810) );
  DFF_X1 inst2_stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S20reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext2[56]),
        .QN(inst2_n2808) );
  DFF_X1 inst2_stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S13reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext2[71])
         );
  DFF_X1 inst2_stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S13reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext2[70])
         );
  DFF_X1 inst2_stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S13reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext2[69])
         );
  DFF_X1 inst2_stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S13reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[68])
         );
  DFF_X1 inst2_stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S13reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[67])
         );
  DFF_X1 inst2_stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S13reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[66])
         );
  DFF_X1 inst2_stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S13reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[65])
         );
  DFF_X1 inst2_stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S13reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[64])
         );
  DFF_X1 inst2_stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S12reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext2[79]),
        .QN(inst2_n1250) );
  DFF_X1 inst2_stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S12reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext2[78]),
        .QN(inst2_n1251) );
  DFF_X1 inst2_stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S12reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext2[77]),
        .QN(inst2_n1252) );
  DFF_X1 inst2_stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S12reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[76]),
        .QN(inst2_n1253) );
  DFF_X1 inst2_stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S12reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[75]),
        .QN(inst2_n1254) );
  DFF_X1 inst2_stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S12reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[74]),
        .QN(inst2_n1255) );
  DFF_X1 inst2_stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S12reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[73]),
        .QN(inst2_n1256) );
  DFF_X1 inst2_stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S12reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[72]),
        .QN(inst2_n1257) );
  DFF_X1 inst2_stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S11reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext2[87]),
        .QN(inst2_n1258) );
  DFF_X1 inst2_stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S11reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext2[86]),
        .QN(inst2_n1259) );
  DFF_X1 inst2_stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S11reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext2[85]),
        .QN(inst2_n1260) );
  DFF_X1 inst2_stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S11reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[84]),
        .QN(inst2_n1261) );
  DFF_X1 inst2_stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S11reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[83]),
        .QN(inst2_n1262) );
  DFF_X1 inst2_stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S11reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[82]),
        .QN(inst2_n1263) );
  DFF_X1 inst2_stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S11reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[81]),
        .QN(inst2_n1264) );
  DFF_X1 inst2_stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S11reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[80]),
        .QN(inst2_n1265) );
  DFF_X1 inst2_stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S10reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext2[95]),
        .QN(inst2_n220) );
  DFF_X1 inst2_stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S10reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext2[94]),
        .QN(inst2_n206) );
  DFF_X1 inst2_stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S10reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext2[93]),
        .QN(inst2_n190) );
  DFF_X1 inst2_stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S10reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext2[92]),
        .QN(inst2_n212) );
  DFF_X1 inst2_stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S10reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext2[91]),
        .QN(inst2_n201) );
  DFF_X1 inst2_stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S10reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext2[90]),
        .QN(inst2_n194) );
  DFF_X1 inst2_stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S10reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext2[89]),
        .QN(inst2_n197) );
  DFF_X1 inst2_stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S10reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext2[88]),
        .QN(inst2_n209) );
  DFF_X1 inst2_stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S03reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext2[103]), .QN(inst2_n1266) );
  DFF_X1 inst2_stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S03reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext2[102]), .QN(inst2_n1267) );
  DFF_X1 inst2_stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S03reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext2[101]), .QN(inst2_n1268) );
  DFF_X1 inst2_stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S03reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[100]), .QN(inst2_n1269) );
  DFF_X1 inst2_stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S03reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[99]),
        .QN(inst2_n1270) );
  DFF_X1 inst2_stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S03reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[98]),
        .QN(inst2_n1271) );
  DFF_X1 inst2_stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S03reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[97]),
        .QN(inst2_n1272) );
  DFF_X1 inst2_stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S03reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[96]),
        .QN(inst2_n1273) );
  DFF_X1 inst2_stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S02reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext2[111]) );
  DFF_X1 inst2_stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S02reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext2[110]) );
  DFF_X1 inst2_stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S02reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext2[109]) );
  DFF_X1 inst2_stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S02reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[108]) );
  DFF_X1 inst2_stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S02reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[107]) );
  DFF_X1 inst2_stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S02reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[106]) );
  DFF_X1 inst2_stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S02reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[105]) );
  DFF_X1 inst2_stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S02reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[104]) );
  DFF_X1 inst2_stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S01reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext2[119]), .QN(inst2_n2855) );
  DFF_X1 inst2_stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S01reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext2[118]), .QN(inst2_n2856) );
  DFF_X1 inst2_stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S01reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext2[117]), .QN(inst2_n2857) );
  DFF_X1 inst2_stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S01reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[116]), .QN(inst2_n2858) );
  DFF_X1 inst2_stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S01reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[115]), .QN(inst2_n2859) );
  DFF_X1 inst2_stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S01reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[114]), .QN(inst2_n2860) );
  DFF_X1 inst2_stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S01reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[113]), .QN(inst2_n2861) );
  DFF_X1 inst2_stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S01reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[112]), .QN(inst2_n2862) );
  DFF_X1 inst2_stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst2_stateArray_S00reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext2[127]), .QN(inst2_n218) );
  DFF_X1 inst2_stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst2_stateArray_S00reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext2[126]), .QN(inst2_n216) );
  DFF_X1 inst2_stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst2_stateArray_S00reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext2[125]), .QN(inst2_n214) );
  DFF_X1 inst2_stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst2_stateArray_S00reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext2[124]), .QN(inst2_n2799) );
  DFF_X1 inst2_stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst2_stateArray_S00reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext2[123]), .QN(inst2_n202) );
  DFF_X1 inst2_stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst2_stateArray_S00reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext2[122]), .QN(inst2_n2800) );
  DFF_X1 inst2_stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst2_stateArray_S00reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext2[121]), .QN(inst2_n198) );
  DFF_X1 inst2_stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst2_stateArray_S00reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext2[120]), .QN(inst2_n210) );
  DFF_X1 inst2_ctrl_CSenRC_reg_FF_FF ( .D(inst2_n2872), .CK(clk), .QN(
        inst2_n321) );
  DFF_X1 inst2_ctrl_CSselMC_reg_FF_FF ( .D(inst2_n1088), .CK(clk), .Q(
        inst2_ctrl_n6) );
  DFF_X1 inst2_ctrl_seq4_SFF_1_Q_reg_FF_FF ( .D(inst2_ctrl_seq4_SFF_1_n5),
        .CK(clk), .Q(inst2_n2826), .QN(inst2_n236) );
  DFF_X1 inst2_ctrl_seq4_SFF_0_Q_reg_FF_FF ( .D(inst2_ctrl_seq4_SFF_0_n5),
        .CK(clk), .Q(inst2_n143), .QN(inst2_n2811) );
  DFF_X1 inst2_ctrl_seq6_SFF_4_Q_reg_FF_FF ( .D(inst2_ctrl_seq6_SFF_4_n5),
        .CK(clk), .QN(inst2_n1290) );
  DFF_X1 inst2_ctrl_seq6_SFF_3_Q_reg_FF_FF ( .D(inst2_ctrl_seq6_SFF_3_n5),
        .CK(clk), .QN(inst2_n231) );
  DFF_X1 inst2_ctrl_seq6_SFF_2_Q_reg_FF_FF ( .D(inst2_ctrl_seq6_SFF_2_n5),
        .CK(clk), .QN(inst2_n233) );
  DFF_X1 inst2_ctrl_seq6_SFF_1_Q_reg_FF_FF ( .D(inst2_ctrl_seq6_SFF_1_n5),
        .CK(clk), .QN(inst2_n230) );
  DFF_X1 inst2_ctrl_seq6_SFF_0_Q_reg_FF_FF ( .D(inst2_ctrl_seq6_SFF_0_n5),
        .CK(clk), .QN(inst2_n232) );
  OAI21_X1 inst3_U1163 ( .B1(inst3_n2801), .B2(inst3_n2800), .A(inst3_n2799),
        .ZN(inst3_n1088) );
  OAI211_X1 inst3_U1162 ( .C1(inst3_n2798), .C2(inst3_n2797), .A(inst3_n2796),
        .B(inst3_n2795), .ZN(inst3_stateArray_S23reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst3_U1161 ( .B1(inst3_n2794), .B2(ciphertext3[49]), .A(
        inst3_n2793), .ZN(inst3_n2795) );
  OAI22_X1 inst3_U1160 ( .A1(inst3_n191), .A2(inst3_n2780), .B1(inst3_n2792),
        .B2(inst3_n2811), .ZN(inst3_n2793) );
  AOI22_X1 inst3_U1159 ( .A1(done3), .A2(ciphertext3[33]), .B1(plaintext3[33]),
        .B2(inst3_n2806), .ZN(inst3_n2796) );
  XNOR2_X1 inst3_U1158 ( .A(inst3_n2791), .B(inst3_n2790), .ZN(inst3_n2798) );
  AOI22_X1 inst3_U1157 ( .A1(inst3_n191), .A2(inst3_n2789), .B1(inst3_n2788),
        .B2(ciphertext3[25]), .ZN(inst3_n2790) );
  XNOR2_X1 inst3_U1156 ( .A(inst3_n2787), .B(inst3_n2786), .ZN(inst3_n2791) );
  OAI211_X1 inst3_U1155 ( .C1(inst3_n2785), .C2(inst3_n2784), .A(inst3_n2783),
        .B(inst3_n2782), .ZN(inst3_stateArray_S23reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst3_U1154 ( .B1(inst3_n2794), .B2(ciphertext3[50]), .A(
        inst3_n2781), .ZN(inst3_n2782) );
  OAI22_X1 inst3_U1153 ( .A1(inst3_n203), .A2(inst3_n2780), .B1(inst3_n193),
        .B2(inst3_n2792), .ZN(inst3_n2781) );
  AOI22_X1 inst3_U1152 ( .A1(done3), .A2(ciphertext3[34]), .B1(plaintext3[34]),
        .B2(inst3_n2806), .ZN(inst3_n2783) );
  XNOR2_X1 inst3_U1151 ( .A(inst3_n2779), .B(inst3_n2778), .ZN(inst3_n2785) );
  AOI22_X1 inst3_U1150 ( .A1(inst3_n203), .A2(inst3_n2777), .B1(inst3_n2776),
        .B2(ciphertext3[26]), .ZN(inst3_n2778) );
  NOR2_X1 inst3_U1149 ( .A1(inst3_n2775), .A2(inst3_n2812), .ZN(
        inst3_ctrl_seq4_SFF_1_n5) );
  NOR2_X1 inst3_U1148 ( .A1(inst3_n232), .A2(inst3_n2774), .ZN(
        inst3_ctrl_seq6_SFF_1_n5) );
  NOR2_X1 inst3_U1147 ( .A1(inst3_n233), .A2(inst3_n2774), .ZN(
        inst3_ctrl_seq6_SFF_3_n5) );
  OAI211_X1 inst3_U1146 ( .C1(inst3_n2797), .C2(inst3_n2773), .A(inst3_n2772),
        .B(inst3_n2771), .ZN(inst3_stateArray_S23reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst3_U1145 ( .B1(inst3_n2794), .B2(ciphertext3[52]), .A(
        inst3_n2770), .ZN(inst3_n2771) );
  OAI22_X1 inst3_U1144 ( .A1(inst3_n207), .A2(inst3_n2780), .B1(inst3_n2792),
        .B2(inst3_n2822), .ZN(inst3_n2770) );
  AOI22_X1 inst3_U1143 ( .A1(done3), .A2(ciphertext3[36]), .B1(plaintext3[36]),
        .B2(inst3_n2806), .ZN(inst3_n2772) );
  XNOR2_X1 inst3_U1142 ( .A(inst3_n2769), .B(inst3_n2768), .ZN(inst3_n2773) );
  AOI22_X1 inst3_U1141 ( .A1(inst3_n212), .A2(inst3_n2767), .B1(inst3_n2766),
        .B2(ciphertext3[92]), .ZN(inst3_n2768) );
  AOI22_X1 inst3_U1140 ( .A1(inst3_n2789), .A2(inst3_n2765), .B1(inst3_n2764),
        .B2(inst3_n2788), .ZN(inst3_n2769) );
  OAI22_X1 inst3_U1139 ( .A1(inst3_n1080), .A2(inst3_n2763), .B1(inst3_n718),
        .B2(inst3_n2762), .ZN(inst3_calcRCon_n45) );
  OAI21_X1 inst3_U1138 ( .B1(inst3_n499), .B2(inst3_n2762), .A(inst3_n2761),
        .ZN(inst3_calcRCon_n50) );
  OAI221_X1 inst3_U1137 ( .B1(inst3_n1071), .B2(inst3_n444), .C1(inst3_n2803),
        .C2(inst3_n2839), .A(inst3_n2794), .ZN(inst3_n2761) );
  OAI22_X1 inst3_U1136 ( .A1(inst3_n1080), .A2(inst3_n2762), .B1(inst3_n1081),
        .B2(inst3_n2760), .ZN(inst3_calcRCon_n46) );
  OAI21_X1 inst3_U1135 ( .B1(inst3_n1081), .B2(inst3_n2762), .A(inst3_n2759),
        .ZN(inst3_calcRCon_n47) );
  OAI221_X1 inst3_U1134 ( .B1(inst3_n706), .B2(inst3_n1071), .C1(inst3_n2813),
        .C2(inst3_n2803), .A(inst3_n2794), .ZN(inst3_n2759) );
  NAND2_X1 inst3_U1133 ( .A1(inst3_n6), .A2(inst3_n2760), .ZN(inst3_n2762) );
  OAI211_X1 inst3_U1132 ( .C1(inst3_n1233), .C2(inst3_n2763), .A(inst3_n2758),
        .B(inst3_n2757), .ZN(inst3_stateArray_S20reg_gff_1_SFF_0_n5) );
  NAND2_X1 inst3_U1131 ( .A1(inst3_n2753), .A2(ciphertext3[48]), .ZN(
        inst3_n2757) );
  AOI22_X1 inst3_U1130 ( .A1(ciphertext3[56]), .A2(inst3_n2756), .B1(
        plaintext3[56]), .B2(inst3_n2806), .ZN(inst3_n2758) );
  OAI211_X1 inst3_U1129 ( .C1(inst3_n1232), .C2(inst3_n2763), .A(inst3_n2755),
        .B(inst3_n2754), .ZN(inst3_stateArray_S20reg_gff_1_SFF_1_n5) );
  NAND2_X1 inst3_U1128 ( .A1(inst3_n2753), .A2(ciphertext3[49]), .ZN(
        inst3_n2754) );
  AOI22_X1 inst3_U1127 ( .A1(ciphertext3[57]), .A2(inst3_n2756), .B1(
        plaintext3[57]), .B2(inst3_n2806), .ZN(inst3_n2755) );
  OAI211_X1 inst3_U1126 ( .C1(inst3_n1231), .C2(inst3_n2763), .A(inst3_n2752),
        .B(inst3_n2751), .ZN(inst3_stateArray_S20reg_gff_1_SFF_2_n5) );
  NAND2_X1 inst3_U1125 ( .A1(inst3_n2753), .A2(ciphertext3[50]), .ZN(
        inst3_n2751) );
  AOI22_X1 inst3_U1124 ( .A1(inst3_n2750), .A2(ciphertext3[58]), .B1(
        plaintext3[58]), .B2(inst3_n2806), .ZN(inst3_n2752) );
  OAI211_X1 inst3_U1123 ( .C1(inst3_n1230), .C2(inst3_n2763), .A(inst3_n2749),
        .B(inst3_n2748), .ZN(inst3_stateArray_S20reg_gff_1_SFF_3_n5) );
  NAND2_X1 inst3_U1122 ( .A1(inst3_n2753), .A2(ciphertext3[51]), .ZN(
        inst3_n2748) );
  AOI22_X1 inst3_U1121 ( .A1(inst3_n2756), .A2(ciphertext3[59]), .B1(
        plaintext3[59]), .B2(inst3_n2806), .ZN(inst3_n2749) );
  OAI211_X1 inst3_U1120 ( .C1(inst3_n1229), .C2(inst3_n2763), .A(inst3_n2747),
        .B(inst3_n2746), .ZN(inst3_stateArray_S20reg_gff_1_SFF_4_n5) );
  NAND2_X1 inst3_U1119 ( .A1(inst3_n2753), .A2(ciphertext3[52]), .ZN(
        inst3_n2746) );
  AOI22_X1 inst3_U1118 ( .A1(ciphertext3[60]), .A2(inst3_n2750), .B1(
        plaintext3[60]), .B2(inst3_n2806), .ZN(inst3_n2747) );
  OAI211_X1 inst3_U1117 ( .C1(inst3_n1228), .C2(inst3_n2760), .A(inst3_n2745),
        .B(inst3_n2744), .ZN(inst3_stateArray_S20reg_gff_1_SFF_5_n5) );
  NAND2_X1 inst3_U1116 ( .A1(inst3_n2753), .A2(ciphertext3[53]), .ZN(
        inst3_n2744) );
  AOI22_X1 inst3_U1115 ( .A1(ciphertext3[61]), .A2(inst3_n2750), .B1(
        plaintext3[61]), .B2(inst3_n2806), .ZN(inst3_n2745) );
  OAI211_X1 inst3_U1114 ( .C1(inst3_n1227), .C2(inst3_n2763), .A(inst3_n2743),
        .B(inst3_n2742), .ZN(inst3_stateArray_S20reg_gff_1_SFF_6_n5) );
  NAND2_X1 inst3_U1113 ( .A1(inst3_n2753), .A2(ciphertext3[54]), .ZN(
        inst3_n2742) );
  AOI22_X1 inst3_U1112 ( .A1(ciphertext3[62]), .A2(inst3_n2750), .B1(
        plaintext3[62]), .B2(inst3_n2806), .ZN(inst3_n2743) );
  OAI211_X1 inst3_U1111 ( .C1(inst3_n1226), .C2(inst3_n2760), .A(inst3_n2741),
        .B(inst3_n2740), .ZN(inst3_stateArray_S20reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst3_U1110 ( .A1(inst3_n1919), .A2(ciphertext3[55]), .ZN(
        inst3_n2740) );
  AOI22_X1 inst3_U1109 ( .A1(inst3_n2750), .A2(ciphertext3[63]), .B1(
        plaintext3[63]), .B2(inst3_n2806), .ZN(inst3_n2741) );
  OAI211_X1 inst3_U1108 ( .C1(inst3_n1233), .C2(inst3_n2775), .A(inst3_n2739),
        .B(inst3_n2738), .ZN(inst3_stateArray_S21reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst3_U1107 ( .A1(plaintext3[48]), .A2(inst3_n2774), .ZN(
        inst3_n2738) );
  AOI22_X1 inst3_U1106 ( .A1(inst3_n2750), .A2(ciphertext3[48]), .B1(
        inst3_n2794), .B2(ciphertext3[32]), .ZN(inst3_n2739) );
  OAI211_X1 inst3_U1105 ( .C1(inst3_n1232), .C2(inst3_n2775), .A(inst3_n2737),
        .B(inst3_n2736), .ZN(inst3_stateArray_S21reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst3_U1104 ( .A1(plaintext3[49]), .A2(inst3_n2774), .ZN(
        inst3_n2736) );
  AOI22_X1 inst3_U1103 ( .A1(inst3_n1914), .A2(ciphertext3[49]), .B1(
        inst3_n2794), .B2(ciphertext3[33]), .ZN(inst3_n2737) );
  OAI211_X1 inst3_U1102 ( .C1(inst3_n1231), .C2(inst3_n2775), .A(inst3_n2735),
        .B(inst3_n2734), .ZN(inst3_stateArray_S21reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst3_U1101 ( .A1(plaintext3[50]), .A2(inst3_n2774), .ZN(
        inst3_n2734) );
  AOI22_X1 inst3_U1100 ( .A1(inst3_n2750), .A2(ciphertext3[50]), .B1(
        inst3_n2794), .B2(ciphertext3[34]), .ZN(inst3_n2735) );
  OAI211_X1 inst3_U1099 ( .C1(inst3_n1230), .C2(inst3_n2775), .A(inst3_n2733),
        .B(inst3_n2732), .ZN(inst3_stateArray_S21reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst3_U1098 ( .A1(plaintext3[51]), .A2(inst3_n2774), .ZN(
        inst3_n2732) );
  AOI22_X1 inst3_U1097 ( .A1(done3), .A2(ciphertext3[51]), .B1(inst3_n2794),
        .B2(ciphertext3[35]), .ZN(inst3_n2733) );
  OAI211_X1 inst3_U1096 ( .C1(inst3_n1229), .C2(inst3_n2775), .A(inst3_n2731),
        .B(inst3_n2730), .ZN(inst3_stateArray_S21reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst3_U1095 ( .A1(plaintext3[52]), .A2(inst3_n2774), .ZN(
        inst3_n2730) );
  AOI22_X1 inst3_U1094 ( .A1(inst3_n2750), .A2(ciphertext3[52]), .B1(
        inst3_n2794), .B2(ciphertext3[36]), .ZN(inst3_n2731) );
  OAI211_X1 inst3_U1093 ( .C1(inst3_n1228), .C2(inst3_n2775), .A(inst3_n2729),
        .B(inst3_n2728), .ZN(inst3_stateArray_S21reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst3_U1092 ( .A1(plaintext3[53]), .A2(inst3_n2727), .ZN(
        inst3_n2728) );
  AOI22_X1 inst3_U1091 ( .A1(done3), .A2(ciphertext3[53]), .B1(inst3_n2794),
        .B2(ciphertext3[37]), .ZN(inst3_n2729) );
  OAI211_X1 inst3_U1090 ( .C1(inst3_n1227), .C2(inst3_n2775), .A(inst3_n2726),
        .B(inst3_n2725), .ZN(inst3_stateArray_S21reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst3_U1089 ( .A1(plaintext3[54]), .A2(inst3_n2774), .ZN(
        inst3_n2725) );
  AOI22_X1 inst3_U1088 ( .A1(inst3_n2750), .A2(ciphertext3[54]), .B1(
        inst3_n2794), .B2(ciphertext3[38]), .ZN(inst3_n2726) );
  OAI211_X1 inst3_U1087 ( .C1(inst3_n1226), .C2(inst3_n2775), .A(inst3_n2724),
        .B(inst3_n2723), .ZN(inst3_stateArray_S21reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst3_U1086 ( .A1(plaintext3[55]), .A2(inst3_n2727), .ZN(
        inst3_n2723) );
  AOI22_X1 inst3_U1085 ( .A1(done3), .A2(ciphertext3[55]), .B1(inst3_n2794),
        .B2(ciphertext3[39]), .ZN(inst3_n2724) );
  OAI21_X1 inst3_U1084 ( .B1(inst3_n1221), .B2(inst3_n2775), .A(inst3_n2722),
        .ZN(inst3_stateArray_S22reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst3_U1083 ( .B1(plaintext3[44]), .B2(inst3_n2774), .A(inst3_n2721), .ZN(inst3_n2722) );
  OAI22_X1 inst3_U1082 ( .A1(inst3_n1229), .A2(inst3_n2720), .B1(inst3_n2763),
        .B2(inst3_n2822), .ZN(inst3_n2721) );
  OAI21_X1 inst3_U1081 ( .B1(inst3_n2775), .B2(inst3_n2836), .A(inst3_n2719),
        .ZN(inst3_stateArray_S30reg_gff_1_SFF_0_n5) );
  AOI21_X1 inst3_U1080 ( .B1(plaintext3[24]), .B2(inst3_n2506), .A(inst3_n2718), .ZN(inst3_n2719) );
  OAI22_X1 inst3_U1079 ( .A1(inst3_n199), .A2(inst3_n2720), .B1(inst3_n1201),
        .B2(inst3_n2760), .ZN(inst3_n2718) );
  OAI21_X1 inst3_U1078 ( .B1(inst3_n2775), .B2(inst3_n2835), .A(inst3_n2717),
        .ZN(inst3_stateArray_S30reg_gff_1_SFF_1_n5) );
  AOI21_X1 inst3_U1077 ( .B1(plaintext3[25]), .B2(inst3_n2527), .A(inst3_n2716), .ZN(inst3_n2717) );
  OAI22_X1 inst3_U1076 ( .A1(inst3_n191), .A2(inst3_n2715), .B1(inst3_n1200),
        .B2(inst3_n2760), .ZN(inst3_n2716) );
  OAI21_X1 inst3_U1075 ( .B1(inst3_n2775), .B2(inst3_n2834), .A(inst3_n2714),
        .ZN(inst3_stateArray_S30reg_gff_1_SFF_2_n5) );
  AOI21_X1 inst3_U1074 ( .B1(plaintext3[26]), .B2(inst3_n2713), .A(inst3_n2712), .ZN(inst3_n2714) );
  OAI22_X1 inst3_U1073 ( .A1(inst3_n203), .A2(inst3_n2720), .B1(inst3_n1199),
        .B2(inst3_n2760), .ZN(inst3_n2712) );
  OAI21_X1 inst3_U1072 ( .B1(inst3_n2775), .B2(inst3_n2833), .A(inst3_n2711),
        .ZN(inst3_stateArray_S30reg_gff_1_SFF_3_n5) );
  AOI21_X1 inst3_U1071 ( .B1(plaintext3[27]), .B2(inst3_n2710), .A(inst3_n2709), .ZN(inst3_n2711) );
  OAI22_X1 inst3_U1070 ( .A1(inst3_n1198), .A2(inst3_n2763), .B1(inst3_n2708),
        .B2(inst3_n2821), .ZN(inst3_n2709) );
  OAI21_X1 inst3_U1069 ( .B1(inst3_n2775), .B2(inst3_n2832), .A(inst3_n2707),
        .ZN(inst3_stateArray_S30reg_gff_1_SFF_4_n5) );
  AOI21_X1 inst3_U1068 ( .B1(plaintext3[28]), .B2(inst3_n2713), .A(inst3_n2706), .ZN(inst3_n2707) );
  OAI22_X1 inst3_U1067 ( .A1(inst3_n207), .A2(inst3_n2715), .B1(inst3_n1197),
        .B2(inst3_n2760), .ZN(inst3_n2706) );
  OAI21_X1 inst3_U1066 ( .B1(inst3_n2775), .B2(inst3_n2831), .A(inst3_n2705),
        .ZN(inst3_stateArray_S30reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst3_U1065 ( .B1(plaintext3[29]), .B2(inst3_n2710), .A(inst3_n2704), .ZN(inst3_n2705) );
  OAI22_X1 inst3_U1064 ( .A1(inst3_n1196), .A2(inst3_n2763), .B1(inst3_n2708),
        .B2(inst3_n2807), .ZN(inst3_n2704) );
  OAI21_X1 inst3_U1063 ( .B1(inst3_n2775), .B2(inst3_n2829), .A(inst3_n2703),
        .ZN(inst3_stateArray_S30reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst3_U1062 ( .B1(plaintext3[30]), .B2(inst3_n2506), .A(inst3_n2702), .ZN(inst3_n2703) );
  OAI22_X1 inst3_U1061 ( .A1(inst3_n215), .A2(inst3_n2720), .B1(inst3_n1195),
        .B2(inst3_n2760), .ZN(inst3_n2702) );
  OAI21_X1 inst3_U1060 ( .B1(inst3_n2775), .B2(inst3_n2830), .A(inst3_n2701),
        .ZN(inst3_stateArray_S30reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst3_U1059 ( .B1(plaintext3[31]), .B2(inst3_n2710), .A(inst3_n2700), .ZN(inst3_n2701) );
  OAI22_X1 inst3_U1058 ( .A1(inst3_n1194), .A2(inst3_n2763), .B1(inst3_n2708),
        .B2(inst3_n2808), .ZN(inst3_n2700) );
  OAI21_X1 inst3_U1057 ( .B1(inst3_n1201), .B2(inst3_n2775), .A(inst3_n2699),
        .ZN(inst3_stateArray_S32reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst3_U1056 ( .B1(plaintext3[8]), .B2(inst3_n2655), .A(inst3_n2698),
        .ZN(inst3_n2699) );
  OAI22_X1 inst3_U1055 ( .A1(inst3_n1209), .A2(inst3_n2715), .B1(inst3_n2763),
        .B2(inst3_n2836), .ZN(inst3_n2698) );
  OAI21_X1 inst3_U1054 ( .B1(inst3_n1200), .B2(inst3_n2775), .A(inst3_n2697),
        .ZN(inst3_stateArray_S32reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst3_U1053 ( .B1(plaintext3[9]), .B2(inst3_n2710), .A(inst3_n2696),
        .ZN(inst3_n2697) );
  OAI22_X1 inst3_U1052 ( .A1(inst3_n1208), .A2(inst3_n2715), .B1(inst3_n2760),
        .B2(inst3_n2835), .ZN(inst3_n2696) );
  OAI21_X1 inst3_U1051 ( .B1(inst3_n1199), .B2(inst3_n2775), .A(inst3_n2695),
        .ZN(inst3_stateArray_S32reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst3_U1050 ( .B1(plaintext3[10]), .B2(inst3_n2713), .A(inst3_n2694), .ZN(inst3_n2695) );
  OAI22_X1 inst3_U1049 ( .A1(inst3_n1207), .A2(inst3_n2715), .B1(inst3_n2760),
        .B2(inst3_n2834), .ZN(inst3_n2694) );
  OAI21_X1 inst3_U1048 ( .B1(inst3_n1198), .B2(inst3_n2775), .A(inst3_n2693),
        .ZN(inst3_stateArray_S32reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst3_U1047 ( .B1(plaintext3[11]), .B2(inst3_n2710), .A(inst3_n2692), .ZN(inst3_n2693) );
  OAI22_X1 inst3_U1046 ( .A1(inst3_n1206), .A2(inst3_n2715), .B1(inst3_n2760),
        .B2(inst3_n2833), .ZN(inst3_n2692) );
  OAI21_X1 inst3_U1045 ( .B1(inst3_n1197), .B2(inst3_n2775), .A(inst3_n2691),
        .ZN(inst3_stateArray_S32reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst3_U1044 ( .B1(plaintext3[12]), .B2(inst3_n2710), .A(inst3_n2690), .ZN(inst3_n2691) );
  OAI22_X1 inst3_U1043 ( .A1(inst3_n1205), .A2(inst3_n2715), .B1(inst3_n2760),
        .B2(inst3_n2832), .ZN(inst3_n2690) );
  OAI21_X1 inst3_U1042 ( .B1(inst3_n1196), .B2(inst3_n2775), .A(inst3_n2689),
        .ZN(inst3_stateArray_S32reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst3_U1041 ( .B1(plaintext3[13]), .B2(inst3_n2710), .A(inst3_n2688), .ZN(inst3_n2689) );
  OAI22_X1 inst3_U1040 ( .A1(inst3_n1204), .A2(inst3_n2715), .B1(inst3_n2763),
        .B2(inst3_n2831), .ZN(inst3_n2688) );
  OAI21_X1 inst3_U1039 ( .B1(inst3_n1195), .B2(inst3_n2775), .A(inst3_n2687),
        .ZN(inst3_stateArray_S32reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst3_U1038 ( .B1(plaintext3[14]), .B2(inst3_n2710), .A(inst3_n2686), .ZN(inst3_n2687) );
  OAI22_X1 inst3_U1037 ( .A1(inst3_n1203), .A2(inst3_n2708), .B1(inst3_n2760),
        .B2(inst3_n2829), .ZN(inst3_n2686) );
  OAI21_X1 inst3_U1036 ( .B1(inst3_n1194), .B2(inst3_n2775), .A(inst3_n2685),
        .ZN(inst3_stateArray_S32reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst3_U1035 ( .B1(plaintext3[15]), .B2(inst3_n2710), .A(inst3_n2684), .ZN(inst3_n2685) );
  OAI22_X1 inst3_U1034 ( .A1(inst3_n1202), .A2(inst3_n2715), .B1(inst3_n2760),
        .B2(inst3_n2830), .ZN(inst3_n2684) );
  INV_X1 inst3_U1033 ( .A(inst3_n2756), .ZN(inst3_n2715) );
  OAI211_X1 inst3_U1032 ( .C1(inst3_n706), .C2(inst3_n2794), .A(inst3_n6), .B(
        inst3_n2683), .ZN(inst3_calcRCon_n48) );
  OAI221_X1 inst3_U1031 ( .B1(inst3_n581), .B2(inst3_n1071), .C1(inst3_n2838),
        .C2(inst3_n2803), .A(inst3_n2794), .ZN(inst3_n2683) );
  OAI21_X1 inst3_U1030 ( .B1(inst3_n1225), .B2(inst3_n2775), .A(inst3_n2682),
        .ZN(inst3_stateArray_S22reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst3_U1029 ( .B1(plaintext3[40]), .B2(inst3_n2710), .A(inst3_n2681), .ZN(inst3_n2682) );
  OAI22_X1 inst3_U1028 ( .A1(inst3_n1233), .A2(inst3_n2720), .B1(inst3_n2760),
        .B2(inst3_n2810), .ZN(inst3_n2681) );
  OAI211_X1 inst3_U1027 ( .C1(inst3_n1204), .C2(inst3_n2775), .A(inst3_n2680),
        .B(inst3_n2679), .ZN(inst3_stateArray_S31reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst3_U1026 ( .A1(plaintext3[21]), .A2(inst3_n2774), .ZN(
        inst3_n2679) );
  AOI22_X1 inst3_U1025 ( .A1(inst3_n2750), .A2(ciphertext3[21]), .B1(
        inst3_n2794), .B2(ciphertext3[29]), .ZN(inst3_n2680) );
  OAI21_X1 inst3_U1024 ( .B1(inst3_n1224), .B2(inst3_n2775), .A(inst3_n2678),
        .ZN(inst3_stateArray_S22reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst3_U1023 ( .B1(plaintext3[41]), .B2(inst3_n2710), .A(inst3_n2677), .ZN(inst3_n2678) );
  OAI22_X1 inst3_U1022 ( .A1(inst3_n1232), .A2(inst3_n2720), .B1(inst3_n2763),
        .B2(inst3_n2811), .ZN(inst3_n2677) );
  OAI21_X1 inst3_U1021 ( .B1(inst3_n1223), .B2(inst3_n2775), .A(inst3_n2676),
        .ZN(inst3_stateArray_S22reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst3_U1020 ( .B1(plaintext3[42]), .B2(inst3_n2710), .A(inst3_n2675), .ZN(inst3_n2676) );
  OAI22_X1 inst3_U1019 ( .A1(inst3_n193), .A2(inst3_n2763), .B1(inst3_n1231),
        .B2(inst3_n2720), .ZN(inst3_n2675) );
  OAI21_X1 inst3_U1018 ( .B1(inst3_n1222), .B2(inst3_n2775), .A(inst3_n2674),
        .ZN(inst3_stateArray_S22reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst3_U1017 ( .B1(plaintext3[43]), .B2(inst3_n2713), .A(inst3_n2673), .ZN(inst3_n2674) );
  OAI22_X1 inst3_U1016 ( .A1(inst3_n196), .A2(inst3_n2763), .B1(inst3_n1230),
        .B2(inst3_n2720), .ZN(inst3_n2673) );
  OAI21_X1 inst3_U1015 ( .B1(inst3_n1219), .B2(inst3_n2775), .A(inst3_n2672),
        .ZN(inst3_stateArray_S22reg_gff_1_SFF_6_n6) );
  AOI21_X1 inst3_U1014 ( .B1(plaintext3[46]), .B2(inst3_n2713), .A(inst3_n2671), .ZN(inst3_n2672) );
  OAI22_X1 inst3_U1013 ( .A1(inst3_n1227), .A2(inst3_n2720), .B1(inst3_n2760),
        .B2(inst3_n2809), .ZN(inst3_n2671) );
  OAI21_X1 inst3_U1012 ( .B1(inst3_n1218), .B2(inst3_n2775), .A(inst3_n2670),
        .ZN(inst3_stateArray_S22reg_gff_1_SFF_7_n6) );
  AOI21_X1 inst3_U1011 ( .B1(plaintext3[47]), .B2(inst3_n2713), .A(inst3_n2669), .ZN(inst3_n2670) );
  OAI22_X1 inst3_U1010 ( .A1(inst3_n219), .A2(inst3_n2763), .B1(inst3_n1226),
        .B2(inst3_n2720), .ZN(inst3_n2669) );
  OAI211_X1 inst3_U1009 ( .C1(inst3_n1184), .C2(inst3_n2668), .A(inst3_n2667),
        .B(inst3_n2666), .ZN(inst3_KeyArray_S01reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst3_U1008 ( .A1(inst3_n2665), .A2(inst3_n137), .ZN(inst3_n2666)
         );
  AOI22_X1 inst3_U1007 ( .A1(inst3_n2584), .A2(inst3_n2841), .B1(key3[113]),
        .B2(inst3_n2806), .ZN(inst3_n2667) );
  OAI211_X1 inst3_U1006 ( .C1(inst3_n1183), .C2(inst3_n2668), .A(inst3_n2664),
        .B(inst3_n2663), .ZN(inst3_KeyArray_S01reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst3_U1005 ( .A1(inst3_n2662), .A2(inst3_n136), .ZN(inst3_n2663)
         );
  AOI22_X1 inst3_U1004 ( .A1(inst3_n2538), .A2(inst3_n2828), .B1(key3[114]),
        .B2(inst3_n2806), .ZN(inst3_n2664) );
  OAI211_X1 inst3_U1003 ( .C1(inst3_n1182), .C2(inst3_n2668), .A(inst3_n2661),
        .B(inst3_n2660), .ZN(inst3_KeyArray_S01reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst3_U1002 ( .A1(inst3_n2665), .A2(inst3_n135), .ZN(inst3_n2660)
         );
  AOI22_X1 inst3_U1001 ( .A1(inst3_n2543), .A2(inst3_n2827), .B1(key3[115]),
        .B2(inst3_n2806), .ZN(inst3_n2661) );
  OAI211_X1 inst3_U1000 ( .C1(inst3_n1181), .C2(inst3_n2668), .A(inst3_n2659),
        .B(inst3_n2658), .ZN(inst3_KeyArray_S01reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst3_U999 ( .A1(inst3_n2665), .A2(inst3_n134), .ZN(inst3_n2658) );
  AOI22_X1 inst3_U998 ( .A1(inst3_n2487), .A2(inst3_n2840), .B1(key3[116]),
        .B2(inst3_n2806), .ZN(inst3_n2659) );
  OAI211_X1 inst3_U997 ( .C1(inst3_n1180), .C2(inst3_n2668), .A(inst3_n2657),
        .B(inst3_n2656), .ZN(inst3_KeyArray_S01reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst3_U996 ( .A1(inst3_n2665), .A2(inst3_n133), .ZN(inst3_n2656) );
  AOI22_X1 inst3_U995 ( .A1(inst3_n2538), .A2(inst3_n2826), .B1(key3[117]),
        .B2(inst3_n2655), .ZN(inst3_n2657) );
  OAI211_X1 inst3_U994 ( .C1(inst3_n1179), .C2(inst3_n2668), .A(inst3_n2654),
        .B(inst3_n2653), .ZN(inst3_KeyArray_S01reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst3_U993 ( .A1(inst3_n2665), .A2(inst3_n132), .ZN(inst3_n2653) );
  AOI22_X1 inst3_U992 ( .A1(inst3_n2543), .A2(inst3_n2825), .B1(key3[118]),
        .B2(inst3_n2655), .ZN(inst3_n2654) );
  OAI211_X1 inst3_U991 ( .C1(inst3_n1178), .C2(inst3_n2668), .A(inst3_n2652),
        .B(inst3_n2651), .ZN(inst3_KeyArray_S01reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst3_U990 ( .A1(inst3_n2665), .A2(inst3_n131), .ZN(inst3_n2651) );
  AOI22_X1 inst3_U989 ( .A1(inst3_n2487), .A2(inst3_n2824), .B1(key3[119]),
        .B2(inst3_n2655), .ZN(inst3_n2652) );
  OAI21_X1 inst3_U988 ( .B1(inst3_n2648), .B2(inst3_n2873), .A(inst3_n2650),
        .ZN(inst3_KeyArray_S02reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst3_U987 ( .B1(key3[104]), .B2(inst3_n2713), .A(inst3_n2649),
        .ZN(inst3_n2650) );
  OAI22_X1 inst3_U986 ( .A1(inst3_n1177), .A2(inst3_n2780), .B1(inst3_n1185),
        .B2(inst3_n2799), .ZN(inst3_n2649) );
  OAI21_X1 inst3_U985 ( .B1(inst3_n2648), .B2(inst3_n2872), .A(inst3_n2647),
        .ZN(inst3_KeyArray_S02reg_gff_1_SFF_1_n6) );
  AOI21_X1 inst3_U984 ( .B1(key3[105]), .B2(inst3_n2713), .A(inst3_n2646),
        .ZN(inst3_n2647) );
  OAI22_X1 inst3_U983 ( .A1(inst3_n1176), .A2(inst3_n2780), .B1(inst3_n1184),
        .B2(inst3_n2799), .ZN(inst3_n2646) );
  OAI21_X1 inst3_U982 ( .B1(inst3_n2648), .B2(inst3_n2871), .A(inst3_n2645),
        .ZN(inst3_KeyArray_S02reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst3_U981 ( .B1(key3[106]), .B2(inst3_n2713), .A(inst3_n2644),
        .ZN(inst3_n2645) );
  OAI22_X1 inst3_U980 ( .A1(inst3_n1175), .A2(inst3_n2780), .B1(inst3_n1183),
        .B2(inst3_n2799), .ZN(inst3_n2644) );
  OAI21_X1 inst3_U979 ( .B1(inst3_n2648), .B2(inst3_n2870), .A(inst3_n2643),
        .ZN(inst3_KeyArray_S02reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst3_U978 ( .B1(key3[107]), .B2(inst3_n2713), .A(inst3_n2642),
        .ZN(inst3_n2643) );
  OAI22_X1 inst3_U977 ( .A1(inst3_n1174), .A2(inst3_n2780), .B1(inst3_n1182),
        .B2(inst3_n2799), .ZN(inst3_n2642) );
  OAI21_X1 inst3_U976 ( .B1(inst3_n2648), .B2(inst3_n2869), .A(inst3_n2641),
        .ZN(inst3_KeyArray_S02reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst3_U975 ( .B1(key3[108]), .B2(inst3_n2713), .A(inst3_n2640),
        .ZN(inst3_n2641) );
  OAI22_X1 inst3_U974 ( .A1(inst3_n1173), .A2(inst3_n2780), .B1(inst3_n1181),
        .B2(inst3_n2799), .ZN(inst3_n2640) );
  OAI21_X1 inst3_U973 ( .B1(inst3_n2648), .B2(inst3_n2868), .A(inst3_n2639),
        .ZN(inst3_KeyArray_S02reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst3_U972 ( .B1(key3[109]), .B2(inst3_n2713), .A(inst3_n2638),
        .ZN(inst3_n2639) );
  OAI22_X1 inst3_U971 ( .A1(inst3_n1172), .A2(inst3_n2780), .B1(inst3_n1180),
        .B2(inst3_n2799), .ZN(inst3_n2638) );
  OAI21_X1 inst3_U970 ( .B1(inst3_n2648), .B2(inst3_n2867), .A(inst3_n2637),
        .ZN(inst3_KeyArray_S02reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst3_U969 ( .B1(key3[110]), .B2(inst3_n2713), .A(inst3_n2636),
        .ZN(inst3_n2637) );
  OAI22_X1 inst3_U968 ( .A1(inst3_n1171), .A2(inst3_n2780), .B1(inst3_n1179),
        .B2(inst3_n2799), .ZN(inst3_n2636) );
  OAI21_X1 inst3_U967 ( .B1(inst3_n2648), .B2(inst3_n2866), .A(inst3_n2635),
        .ZN(inst3_KeyArray_S02reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst3_U966 ( .B1(key3[111]), .B2(inst3_n2713), .A(inst3_n2634),
        .ZN(inst3_n2635) );
  OAI22_X1 inst3_U965 ( .A1(inst3_n1170), .A2(inst3_n2780), .B1(inst3_n1178),
        .B2(inst3_n2799), .ZN(inst3_n2634) );
  INV_X2 inst3_U964 ( .A(inst3_n6), .ZN(inst3_n2713) );
  OAI21_X1 inst3_U963 ( .B1(inst3_n2648), .B2(inst3_n2857), .A(inst3_n2633),
        .ZN(inst3_KeyArray_S03reg_gff_1_SFF_0_n5) );
  AOI21_X1 inst3_U962 ( .B1(key3[96]), .B2(inst3_n2710), .A(inst3_n2632), .ZN(
        inst3_n2633) );
  OAI22_X1 inst3_U961 ( .A1(inst3_n1169), .A2(inst3_n2780), .B1(inst3_n1177),
        .B2(inst3_n2799), .ZN(inst3_n2632) );
  OAI21_X1 inst3_U960 ( .B1(inst3_n2648), .B2(inst3_n2856), .A(inst3_n2631),
        .ZN(inst3_KeyArray_S03reg_gff_1_SFF_1_n5) );
  AOI21_X1 inst3_U959 ( .B1(key3[97]), .B2(inst3_n2713), .A(inst3_n2630), .ZN(
        inst3_n2631) );
  OAI22_X1 inst3_U958 ( .A1(inst3_n1168), .A2(inst3_n2780), .B1(inst3_n1176),
        .B2(inst3_n2799), .ZN(inst3_n2630) );
  OAI21_X1 inst3_U957 ( .B1(inst3_n2648), .B2(inst3_n2855), .A(inst3_n2629),
        .ZN(inst3_KeyArray_S03reg_gff_1_SFF_2_n5) );
  AOI21_X1 inst3_U956 ( .B1(key3[98]), .B2(inst3_n2713), .A(inst3_n2628), .ZN(
        inst3_n2629) );
  OAI22_X1 inst3_U955 ( .A1(inst3_n1167), .A2(inst3_n2461), .B1(inst3_n1175),
        .B2(inst3_n2799), .ZN(inst3_n2628) );
  OAI21_X1 inst3_U954 ( .B1(inst3_n2648), .B2(inst3_n2854), .A(inst3_n2627),
        .ZN(inst3_KeyArray_S03reg_gff_1_SFF_3_n5) );
  AOI21_X1 inst3_U953 ( .B1(key3[99]), .B2(inst3_n2727), .A(inst3_n2626), .ZN(
        inst3_n2627) );
  OAI22_X1 inst3_U952 ( .A1(inst3_n1166), .A2(inst3_n2461), .B1(inst3_n1174),
        .B2(inst3_n2799), .ZN(inst3_n2626) );
  OAI21_X1 inst3_U951 ( .B1(inst3_n2648), .B2(inst3_n2853), .A(inst3_n2625),
        .ZN(inst3_KeyArray_S03reg_gff_1_SFF_4_n5) );
  AOI21_X1 inst3_U950 ( .B1(key3[100]), .B2(inst3_n2774), .A(inst3_n2624),
        .ZN(inst3_n2625) );
  OAI22_X1 inst3_U949 ( .A1(inst3_n1165), .A2(inst3_n2461), .B1(inst3_n1173),
        .B2(inst3_n2799), .ZN(inst3_n2624) );
  OAI21_X1 inst3_U948 ( .B1(inst3_n2648), .B2(inst3_n2852), .A(inst3_n2623),
        .ZN(inst3_KeyArray_S03reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst3_U947 ( .B1(key3[101]), .B2(inst3_n2593), .A(inst3_n2622),
        .ZN(inst3_n2623) );
  OAI22_X1 inst3_U946 ( .A1(inst3_n1164), .A2(inst3_n2461), .B1(inst3_n1172),
        .B2(inst3_n2799), .ZN(inst3_n2622) );
  OAI21_X1 inst3_U945 ( .B1(inst3_n2648), .B2(inst3_n2851), .A(inst3_n2621),
        .ZN(inst3_KeyArray_S03reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst3_U944 ( .B1(key3[102]), .B2(inst3_n2593), .A(inst3_n2620),
        .ZN(inst3_n2621) );
  OAI22_X1 inst3_U943 ( .A1(inst3_n1163), .A2(inst3_n2780), .B1(inst3_n1171),
        .B2(inst3_n2799), .ZN(inst3_n2620) );
  OAI21_X1 inst3_U942 ( .B1(inst3_n2648), .B2(inst3_n2850), .A(inst3_n2619),
        .ZN(inst3_KeyArray_S03reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst3_U941 ( .B1(key3[103]), .B2(inst3_n2593), .A(inst3_n2618),
        .ZN(inst3_n2619) );
  OAI22_X1 inst3_U940 ( .A1(inst3_n1162), .A2(inst3_n2668), .B1(inst3_n1170),
        .B2(inst3_n2799), .ZN(inst3_n2618) );
  OAI21_X1 inst3_U939 ( .B1(inst3_n2648), .B2(inst3_n2865), .A(inst3_n2617),
        .ZN(inst3_KeyArray_S10reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst3_U938 ( .B1(key3[88]), .B2(inst3_n2713), .A(inst3_n2616), .ZN(
        inst3_n2617) );
  OAI22_X1 inst3_U937 ( .A1(inst3_n1169), .A2(inst3_n2799), .B1(inst3_n1161),
        .B2(inst3_n2780), .ZN(inst3_n2616) );
  OAI211_X1 inst3_U936 ( .C1(inst3_n1168), .C2(inst3_n2799), .A(inst3_n2615),
        .B(inst3_n2614), .ZN(inst3_KeyArray_S10reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst3_U935 ( .A1(inst3_n2665), .A2(inst3_n121), .ZN(inst3_n2614) );
  AOI22_X1 inst3_U934 ( .A1(inst3_n137), .A2(inst3_n2613), .B1(key3[89]), .B2(
        inst3_n2655), .ZN(inst3_n2615) );
  OAI211_X1 inst3_U933 ( .C1(inst3_n1167), .C2(inst3_n2799), .A(inst3_n2612),
        .B(inst3_n2611), .ZN(inst3_KeyArray_S10reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst3_U932 ( .A1(inst3_n2665), .A2(inst3_n120), .ZN(inst3_n2611) );
  AOI22_X1 inst3_U931 ( .A1(inst3_n136), .A2(inst3_n2610), .B1(key3[90]), .B2(
        inst3_n2655), .ZN(inst3_n2612) );
  OAI211_X1 inst3_U930 ( .C1(inst3_n1166), .C2(inst3_n2799), .A(inst3_n2609),
        .B(inst3_n2608), .ZN(inst3_KeyArray_S10reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst3_U929 ( .A1(inst3_n2662), .A2(inst3_n119), .ZN(inst3_n2608) );
  AOI22_X1 inst3_U928 ( .A1(inst3_n135), .A2(inst3_n2610), .B1(key3[91]), .B2(
        inst3_n2655), .ZN(inst3_n2609) );
  OAI211_X1 inst3_U927 ( .C1(inst3_n1165), .C2(inst3_n2799), .A(inst3_n2607),
        .B(inst3_n2606), .ZN(inst3_KeyArray_S10reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst3_U926 ( .A1(inst3_n2662), .A2(inst3_n118), .ZN(inst3_n2606) );
  AOI22_X1 inst3_U925 ( .A1(inst3_n134), .A2(inst3_n2610), .B1(key3[92]), .B2(
        inst3_n2655), .ZN(inst3_n2607) );
  OAI211_X1 inst3_U924 ( .C1(inst3_n1164), .C2(inst3_n2799), .A(inst3_n2605),
        .B(inst3_n2604), .ZN(inst3_KeyArray_S10reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst3_U923 ( .A1(inst3_n2662), .A2(inst3_n117), .ZN(inst3_n2604) );
  AOI22_X1 inst3_U922 ( .A1(inst3_n133), .A2(inst3_n2610), .B1(key3[93]), .B2(
        inst3_n2655), .ZN(inst3_n2605) );
  OAI211_X1 inst3_U921 ( .C1(inst3_n1163), .C2(inst3_n2799), .A(inst3_n2603),
        .B(inst3_n2602), .ZN(inst3_KeyArray_S10reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst3_U920 ( .A1(inst3_n2662), .A2(inst3_n116), .ZN(inst3_n2602) );
  AOI22_X1 inst3_U919 ( .A1(inst3_n132), .A2(inst3_n2610), .B1(key3[94]), .B2(
        inst3_n2655), .ZN(inst3_n2603) );
  OAI211_X1 inst3_U918 ( .C1(inst3_n1162), .C2(inst3_n2799), .A(inst3_n2601),
        .B(inst3_n2600), .ZN(inst3_KeyArray_S10reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst3_U917 ( .A1(inst3_n2662), .A2(inst3_n115), .ZN(inst3_n2600) );
  AOI22_X1 inst3_U916 ( .A1(inst3_n131), .A2(inst3_n2613), .B1(key3[95]), .B2(
        inst3_n2655), .ZN(inst3_n2601) );
  OAI211_X1 inst3_U915 ( .C1(inst3_n1161), .C2(inst3_n2799), .A(inst3_n2599),
        .B(inst3_n2598), .ZN(inst3_KeyArray_S11reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst3_U914 ( .A1(inst3_n2662), .A2(inst3_n114), .ZN(inst3_n2598) );
  AOI22_X1 inst3_U913 ( .A1(inst3_n130), .A2(inst3_n2613), .B1(key3[80]), .B2(
        inst3_n2655), .ZN(inst3_n2599) );
  NAND2_X1 inst3_U912 ( .A1(inst3_n2597), .A2(inst3_n2596), .ZN(
        inst3_KeyArray_S11reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U911 ( .A1(inst3_n2584), .A2(inst3_n137), .B1(inst3_n2665),
        .B2(inst3_n113), .ZN(inst3_n2596) );
  AOI22_X1 inst3_U910 ( .A1(inst3_n129), .A2(inst3_n2613), .B1(key3[81]), .B2(
        inst3_n2655), .ZN(inst3_n2597) );
  INV_X1 inst3_U909 ( .A(inst3_n6), .ZN(inst3_n2655) );
  NAND2_X1 inst3_U908 ( .A1(inst3_n2595), .A2(inst3_n2594), .ZN(
        inst3_KeyArray_S11reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U907 ( .A1(inst3_n2538), .A2(inst3_n136), .B1(inst3_n2665),
        .B2(inst3_n112), .ZN(inst3_n2594) );
  AOI22_X1 inst3_U906 ( .A1(inst3_n128), .A2(inst3_n2613), .B1(key3[82]), .B2(
        inst3_n2593), .ZN(inst3_n2595) );
  NAND2_X1 inst3_U905 ( .A1(inst3_n2592), .A2(inst3_n2591), .ZN(
        inst3_KeyArray_S11reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U904 ( .A1(inst3_n2543), .A2(inst3_n135), .B1(inst3_n2665),
        .B2(inst3_n111), .ZN(inst3_n2591) );
  AOI22_X1 inst3_U903 ( .A1(inst3_n127), .A2(inst3_n2613), .B1(key3[83]), .B2(
        inst3_n2593), .ZN(inst3_n2592) );
  NAND2_X1 inst3_U902 ( .A1(inst3_n2590), .A2(inst3_n2589), .ZN(
        inst3_KeyArray_S11reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U901 ( .A1(inst3_n2487), .A2(inst3_n134), .B1(inst3_n2665),
        .B2(inst3_n110), .ZN(inst3_n2589) );
  AOI22_X1 inst3_U900 ( .A1(inst3_n126), .A2(inst3_n2613), .B1(key3[84]), .B2(
        inst3_n2593), .ZN(inst3_n2590) );
  NAND2_X1 inst3_U899 ( .A1(inst3_n2588), .A2(inst3_n2587), .ZN(
        inst3_KeyArray_S11reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst3_U898 ( .A1(inst3_n2584), .A2(inst3_n133), .B1(inst3_n2662),
        .B2(inst3_n109), .ZN(inst3_n2587) );
  AOI22_X1 inst3_U897 ( .A1(inst3_n125), .A2(inst3_n2613), .B1(key3[85]), .B2(
        inst3_n2593), .ZN(inst3_n2588) );
  NAND2_X1 inst3_U896 ( .A1(inst3_n2586), .A2(inst3_n2585), .ZN(
        inst3_KeyArray_S11reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst3_U895 ( .A1(inst3_n2584), .A2(inst3_n132), .B1(inst3_n2665),
        .B2(inst3_n108), .ZN(inst3_n2585) );
  AOI22_X1 inst3_U894 ( .A1(inst3_n124), .A2(inst3_n2613), .B1(key3[86]), .B2(
        inst3_n2593), .ZN(inst3_n2586) );
  NAND2_X1 inst3_U893 ( .A1(inst3_n2583), .A2(inst3_n2582), .ZN(
        inst3_KeyArray_S11reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst3_U892 ( .A1(inst3_n2584), .A2(inst3_n131), .B1(inst3_n2665),
        .B2(inst3_n107), .ZN(inst3_n2582) );
  AOI22_X1 inst3_U891 ( .A1(inst3_n123), .A2(inst3_n2613), .B1(key3[87]), .B2(
        inst3_n2593), .ZN(inst3_n2583) );
  OAI21_X1 inst3_U890 ( .B1(inst3_n1185), .B2(inst3_n2648), .A(inst3_n2581),
        .ZN(inst3_KeyArray_S32reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst3_U889 ( .B1(key3[8]), .B2(inst3_n2593), .A(inst3_n2580), .ZN(
        inst3_n2581) );
  OAI22_X1 inst3_U888 ( .A1(inst3_n1089), .A2(inst3_n2668), .B1(inst3_n1097),
        .B2(inst3_n2799), .ZN(inst3_n2580) );
  OAI21_X1 inst3_U887 ( .B1(inst3_n1183), .B2(inst3_n2648), .A(inst3_n2579),
        .ZN(inst3_KeyArray_S32reg_gff_1_SFF_2_n6) );
  AOI21_X1 inst3_U886 ( .B1(key3[10]), .B2(inst3_n2593), .A(inst3_n2578), .ZN(
        inst3_n2579) );
  OAI22_X1 inst3_U885 ( .A1(inst3_n1087), .A2(inst3_n2780), .B1(inst3_n1095),
        .B2(inst3_n2799), .ZN(inst3_n2578) );
  OAI21_X1 inst3_U884 ( .B1(inst3_n1182), .B2(inst3_n2648), .A(inst3_n2577),
        .ZN(inst3_KeyArray_S32reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst3_U883 ( .B1(key3[11]), .B2(inst3_n2655), .A(inst3_n2576), .ZN(
        inst3_n2577) );
  OAI22_X1 inst3_U882 ( .A1(inst3_n1086), .A2(inst3_n2668), .B1(inst3_n1094),
        .B2(inst3_n2799), .ZN(inst3_n2576) );
  OAI21_X1 inst3_U881 ( .B1(inst3_n1181), .B2(inst3_n2648), .A(inst3_n2575),
        .ZN(inst3_KeyArray_S32reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst3_U880 ( .B1(key3[12]), .B2(inst3_n2713), .A(inst3_n2574), .ZN(
        inst3_n2575) );
  OAI22_X1 inst3_U879 ( .A1(inst3_n1085), .A2(inst3_n2461), .B1(inst3_n1093),
        .B2(inst3_n2799), .ZN(inst3_n2574) );
  OAI21_X1 inst3_U878 ( .B1(inst3_n1180), .B2(inst3_n2648), .A(inst3_n2573),
        .ZN(inst3_KeyArray_S32reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst3_U877 ( .B1(key3[13]), .B2(inst3_n2527), .A(inst3_n2572), .ZN(
        inst3_n2573) );
  OAI22_X1 inst3_U876 ( .A1(inst3_n1084), .A2(inst3_n2668), .B1(inst3_n1092),
        .B2(inst3_n2799), .ZN(inst3_n2572) );
  OAI21_X1 inst3_U875 ( .B1(inst3_n1179), .B2(inst3_n2648), .A(inst3_n2571),
        .ZN(inst3_KeyArray_S32reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst3_U874 ( .B1(key3[14]), .B2(inst3_n2710), .A(inst3_n2570), .ZN(
        inst3_n2571) );
  OAI22_X1 inst3_U873 ( .A1(inst3_n1083), .A2(inst3_n2780), .B1(inst3_n1091),
        .B2(inst3_n2799), .ZN(inst3_n2570) );
  OAI21_X1 inst3_U872 ( .B1(inst3_n1178), .B2(inst3_n2648), .A(inst3_n2569),
        .ZN(inst3_KeyArray_S32reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst3_U871 ( .B1(key3[15]), .B2(inst3_n2506), .A(inst3_n2568), .ZN(
        inst3_n2569) );
  OAI22_X1 inst3_U870 ( .A1(inst3_n1082), .A2(inst3_n2668), .B1(inst3_n1090),
        .B2(inst3_n2799), .ZN(inst3_n2568) );
  OAI21_X1 inst3_U869 ( .B1(inst3_n1161), .B2(inst3_n2648), .A(inst3_n2567),
        .ZN(inst3_KeyArray_S01reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst3_U868 ( .B1(key3[112]), .B2(inst3_n2593), .A(inst3_n2566),
        .ZN(inst3_n2567) );
  OAI22_X1 inst3_U867 ( .A1(inst3_n1193), .A2(inst3_n2799), .B1(inst3_n1185),
        .B2(inst3_n2780), .ZN(inst3_n2566) );
  NAND2_X1 inst3_U866 ( .A1(inst3_n2565), .A2(inst3_n2564), .ZN(
        inst3_KeyArray_S12reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst3_U865 ( .A1(inst3_n2584), .A2(inst3_n130), .B1(inst3_n2662),
        .B2(inst3_n98), .ZN(inst3_n2564) );
  AOI22_X1 inst3_U864 ( .A1(inst3_n22), .A2(inst3_n2613), .B1(key3[72]), .B2(
        inst3_n2593), .ZN(inst3_n2565) );
  NAND2_X1 inst3_U863 ( .A1(inst3_n2563), .A2(inst3_n2562), .ZN(
        inst3_KeyArray_S12reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U862 ( .A1(inst3_n2584), .A2(inst3_n129), .B1(inst3_n2662),
        .B2(inst3_n97), .ZN(inst3_n2562) );
  AOI22_X1 inst3_U861 ( .A1(inst3_n17), .A2(inst3_n2613), .B1(key3[73]), .B2(
        inst3_n2593), .ZN(inst3_n2563) );
  NAND2_X1 inst3_U860 ( .A1(inst3_n2561), .A2(inst3_n2560), .ZN(
        inst3_KeyArray_S12reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U859 ( .A1(inst3_n2584), .A2(inst3_n128), .B1(inst3_n2665),
        .B2(inst3_n96), .ZN(inst3_n2560) );
  AOI22_X1 inst3_U858 ( .A1(inst3_n14), .A2(inst3_n2613), .B1(key3[74]), .B2(
        inst3_n2593), .ZN(inst3_n2561) );
  NAND2_X1 inst3_U857 ( .A1(inst3_n2559), .A2(inst3_n2558), .ZN(
        inst3_KeyArray_S12reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U856 ( .A1(inst3_n2584), .A2(inst3_n127), .B1(inst3_n2662),
        .B2(inst3_n95), .ZN(inst3_n2558) );
  AOI22_X1 inst3_U855 ( .A1(inst3_n12), .A2(inst3_n2613), .B1(key3[75]), .B2(
        inst3_n2593), .ZN(inst3_n2559) );
  NAND2_X1 inst3_U854 ( .A1(inst3_n2557), .A2(inst3_n2556), .ZN(
        inst3_KeyArray_S12reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U853 ( .A1(inst3_n2584), .A2(inst3_n126), .B1(inst3_n2662),
        .B2(inst3_n94), .ZN(inst3_n2556) );
  AOI22_X1 inst3_U852 ( .A1(inst3_n11), .A2(inst3_n2555), .B1(key3[76]), .B2(
        inst3_n2593), .ZN(inst3_n2557) );
  NAND2_X1 inst3_U851 ( .A1(inst3_n2554), .A2(inst3_n2553), .ZN(
        inst3_KeyArray_S12reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst3_U850 ( .A1(inst3_n2584), .A2(inst3_n125), .B1(inst3_n2662),
        .B2(inst3_n93), .ZN(inst3_n2553) );
  AOI22_X1 inst3_U849 ( .A1(inst3_n10), .A2(inst3_n2552), .B1(key3[77]), .B2(
        inst3_n2593), .ZN(inst3_n2554) );
  INV_X1 inst3_U848 ( .A(inst3_n6), .ZN(inst3_n2593) );
  NAND2_X1 inst3_U847 ( .A1(inst3_n2551), .A2(inst3_n2550), .ZN(
        inst3_KeyArray_S12reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst3_U846 ( .A1(inst3_n2584), .A2(inst3_n124), .B1(inst3_n2662),
        .B2(inst3_n92), .ZN(inst3_n2550) );
  AOI22_X1 inst3_U845 ( .A1(inst3_n24), .A2(inst3_n2613), .B1(key3[78]), .B2(
        inst3_n2713), .ZN(inst3_n2551) );
  NAND2_X1 inst3_U844 ( .A1(inst3_n2549), .A2(inst3_n2548), .ZN(
        inst3_KeyArray_S12reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst3_U843 ( .A1(inst3_n2584), .A2(inst3_n123), .B1(inst3_n2662),
        .B2(inst3_n91), .ZN(inst3_n2548) );
  AOI22_X1 inst3_U842 ( .A1(inst3_n9), .A2(inst3_n2555), .B1(key3[79]), .B2(
        inst3_n2713), .ZN(inst3_n2549) );
  NAND2_X1 inst3_U841 ( .A1(inst3_n2547), .A2(inst3_n2546), .ZN(
        inst3_KeyArray_S13reg_gff_1_SFF_0_n5) );
  AOI22_X1 inst3_U840 ( .A1(inst3_n2584), .A2(inst3_n22), .B1(inst3_n2662),
        .B2(inst3_n90), .ZN(inst3_n2546) );
  AOI22_X1 inst3_U839 ( .A1(inst3_n122), .A2(inst3_n2552), .B1(key3[64]), .B2(
        inst3_n2506), .ZN(inst3_n2547) );
  NAND2_X1 inst3_U838 ( .A1(inst3_n2545), .A2(inst3_n2544), .ZN(
        inst3_KeyArray_S13reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst3_U837 ( .A1(inst3_n2543), .A2(inst3_n17), .B1(inst3_n2662),
        .B2(inst3_n89), .ZN(inst3_n2544) );
  AOI22_X1 inst3_U836 ( .A1(inst3_n121), .A2(inst3_n2613), .B1(key3[65]), .B2(
        inst3_n2527), .ZN(inst3_n2545) );
  NAND2_X1 inst3_U835 ( .A1(inst3_n2542), .A2(inst3_n2541), .ZN(
        inst3_KeyArray_S13reg_gff_1_SFF_2_n5) );
  AOI22_X1 inst3_U834 ( .A1(inst3_n2584), .A2(inst3_n14), .B1(inst3_n2662),
        .B2(inst3_n88), .ZN(inst3_n2541) );
  INV_X1 inst3_U833 ( .A(inst3_n2799), .ZN(inst3_n2584) );
  AOI22_X1 inst3_U832 ( .A1(inst3_n120), .A2(inst3_n2555), .B1(key3[66]), .B2(
        inst3_n2713), .ZN(inst3_n2542) );
  NAND2_X1 inst3_U831 ( .A1(inst3_n2540), .A2(inst3_n2539), .ZN(
        inst3_KeyArray_S13reg_gff_1_SFF_3_n5) );
  AOI22_X1 inst3_U830 ( .A1(inst3_n2538), .A2(inst3_n12), .B1(inst3_n2662),
        .B2(inst3_n87), .ZN(inst3_n2539) );
  AOI22_X1 inst3_U829 ( .A1(inst3_n119), .A2(inst3_n2552), .B1(key3[67]), .B2(
        inst3_n2593), .ZN(inst3_n2540) );
  NAND2_X1 inst3_U828 ( .A1(inst3_n2537), .A2(inst3_n2536), .ZN(
        inst3_KeyArray_S13reg_gff_1_SFF_4_n5) );
  AOI22_X1 inst3_U827 ( .A1(inst3_n2538), .A2(inst3_n11), .B1(inst3_n2662),
        .B2(inst3_n86), .ZN(inst3_n2536) );
  AOI22_X1 inst3_U826 ( .A1(inst3_n118), .A2(inst3_n2613), .B1(key3[68]), .B2(
        inst3_n2713), .ZN(inst3_n2537) );
  NAND2_X1 inst3_U825 ( .A1(inst3_n2535), .A2(inst3_n2534), .ZN(
        inst3_KeyArray_S13reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst3_U824 ( .A1(inst3_n2538), .A2(inst3_n10), .B1(inst3_n2662),
        .B2(inst3_n85), .ZN(inst3_n2534) );
  AOI22_X1 inst3_U823 ( .A1(inst3_n117), .A2(inst3_n2552), .B1(key3[69]), .B2(
        inst3_n2593), .ZN(inst3_n2535) );
  NAND2_X1 inst3_U822 ( .A1(inst3_n2533), .A2(inst3_n2532), .ZN(
        inst3_KeyArray_S13reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst3_U821 ( .A1(inst3_n2538), .A2(inst3_n24), .B1(inst3_n2662),
        .B2(inst3_n84), .ZN(inst3_n2532) );
  AOI22_X1 inst3_U820 ( .A1(inst3_n116), .A2(inst3_n2613), .B1(key3[70]), .B2(
        inst3_n2710), .ZN(inst3_n2533) );
  NAND2_X1 inst3_U819 ( .A1(inst3_n2531), .A2(inst3_n2530), .ZN(
        inst3_KeyArray_S13reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst3_U818 ( .A1(inst3_n2538), .A2(inst3_n9), .B1(inst3_n2662),
        .B2(inst3_n83), .ZN(inst3_n2530) );
  AOI22_X1 inst3_U817 ( .A1(inst3_n115), .A2(inst3_n2610), .B1(key3[71]), .B2(
        inst3_n2713), .ZN(inst3_n2531) );
  NAND2_X1 inst3_U816 ( .A1(inst3_n2529), .A2(inst3_n2528), .ZN(
        inst3_KeyArray_S20reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst3_U815 ( .A1(inst3_n2538), .A2(inst3_n122), .B1(inst3_n2662),
        .B2(inst3_n82), .ZN(inst3_n2528) );
  AOI22_X1 inst3_U814 ( .A1(inst3_n114), .A2(inst3_n2552), .B1(key3[56]), .B2(
        inst3_n2527), .ZN(inst3_n2529) );
  NAND2_X1 inst3_U813 ( .A1(inst3_n2526), .A2(inst3_n2525), .ZN(
        inst3_KeyArray_S20reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U812 ( .A1(inst3_n2538), .A2(inst3_n121), .B1(inst3_n2662),
        .B2(inst3_n81), .ZN(inst3_n2525) );
  AOI22_X1 inst3_U811 ( .A1(inst3_n113), .A2(inst3_n2552), .B1(key3[57]), .B2(
        inst3_n2727), .ZN(inst3_n2526) );
  NAND2_X1 inst3_U810 ( .A1(inst3_n2524), .A2(inst3_n2523), .ZN(
        inst3_KeyArray_S20reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U809 ( .A1(inst3_n2538), .A2(inst3_n120), .B1(inst3_n2662),
        .B2(inst3_n80), .ZN(inst3_n2523) );
  AOI22_X1 inst3_U808 ( .A1(inst3_n112), .A2(inst3_n2610), .B1(key3[58]), .B2(
        inst3_n2527), .ZN(inst3_n2524) );
  NAND2_X1 inst3_U807 ( .A1(inst3_n2522), .A2(inst3_n2521), .ZN(
        inst3_KeyArray_S20reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U806 ( .A1(inst3_n2538), .A2(inst3_n119), .B1(inst3_n2662),
        .B2(inst3_n79), .ZN(inst3_n2521) );
  AOI22_X1 inst3_U805 ( .A1(inst3_n111), .A2(inst3_n2555), .B1(key3[59]), .B2(
        inst3_n2527), .ZN(inst3_n2522) );
  NAND2_X1 inst3_U804 ( .A1(inst3_n2520), .A2(inst3_n2519), .ZN(
        inst3_KeyArray_S20reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U803 ( .A1(inst3_n2538), .A2(inst3_n118), .B1(inst3_n78),
        .B2(inst3_n2662), .ZN(inst3_n2519) );
  AOI22_X1 inst3_U802 ( .A1(inst3_n110), .A2(inst3_n2555), .B1(key3[60]), .B2(
        inst3_n2527), .ZN(inst3_n2520) );
  NAND2_X1 inst3_U801 ( .A1(inst3_n2518), .A2(inst3_n2517), .ZN(
        inst3_KeyArray_S20reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst3_U800 ( .A1(inst3_n2538), .A2(inst3_n117), .B1(inst3_n2662),
        .B2(inst3_n77), .ZN(inst3_n2517) );
  AOI22_X1 inst3_U799 ( .A1(inst3_n109), .A2(inst3_n2610), .B1(key3[61]), .B2(
        inst3_n2527), .ZN(inst3_n2518) );
  NAND2_X1 inst3_U798 ( .A1(inst3_n2516), .A2(inst3_n2515), .ZN(
        inst3_KeyArray_S20reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst3_U797 ( .A1(inst3_n2538), .A2(inst3_n116), .B1(inst3_n2662),
        .B2(inst3_n76), .ZN(inst3_n2515) );
  INV_X1 inst3_U796 ( .A(inst3_n2799), .ZN(inst3_n2538) );
  AOI22_X1 inst3_U795 ( .A1(inst3_n108), .A2(inst3_n2610), .B1(key3[62]), .B2(
        inst3_n2527), .ZN(inst3_n2516) );
  NAND2_X1 inst3_U794 ( .A1(inst3_n2514), .A2(inst3_n2513), .ZN(
        inst3_KeyArray_S20reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst3_U793 ( .A1(inst3_n2543), .A2(inst3_n115), .B1(inst3_n2662),
        .B2(inst3_n75), .ZN(inst3_n2513) );
  AOI22_X1 inst3_U792 ( .A1(inst3_n107), .A2(inst3_n2555), .B1(key3[63]), .B2(
        inst3_n2527), .ZN(inst3_n2514) );
  NAND2_X1 inst3_U791 ( .A1(inst3_n2512), .A2(inst3_n2511), .ZN(
        inst3_KeyArray_S21reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst3_U790 ( .A1(inst3_n2543), .A2(inst3_n114), .B1(inst3_n2662),
        .B2(inst3_n74), .ZN(inst3_n2511) );
  AOI22_X1 inst3_U789 ( .A1(inst3_n98), .A2(inst3_n2555), .B1(key3[48]), .B2(
        inst3_n2527), .ZN(inst3_n2512) );
  NAND2_X1 inst3_U788 ( .A1(inst3_n2510), .A2(inst3_n2509), .ZN(
        inst3_KeyArray_S21reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U787 ( .A1(inst3_n2543), .A2(inst3_n113), .B1(inst3_n2662),
        .B2(inst3_n73), .ZN(inst3_n2509) );
  AOI22_X1 inst3_U786 ( .A1(inst3_n97), .A2(inst3_n2613), .B1(key3[49]), .B2(
        inst3_n2527), .ZN(inst3_n2510) );
  NAND2_X1 inst3_U785 ( .A1(inst3_n2508), .A2(inst3_n2507), .ZN(
        inst3_KeyArray_S21reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U784 ( .A1(inst3_n2543), .A2(inst3_n112), .B1(inst3_n2662),
        .B2(inst3_n72), .ZN(inst3_n2507) );
  AOI22_X1 inst3_U783 ( .A1(inst3_n96), .A2(inst3_n2552), .B1(key3[50]), .B2(
        inst3_n2506), .ZN(inst3_n2508) );
  NAND2_X1 inst3_U782 ( .A1(inst3_n2505), .A2(inst3_n2504), .ZN(
        inst3_KeyArray_S21reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U781 ( .A1(inst3_n2543), .A2(inst3_n111), .B1(inst3_n2662),
        .B2(inst3_n71), .ZN(inst3_n2504) );
  AOI22_X1 inst3_U780 ( .A1(inst3_n95), .A2(inst3_n2552), .B1(key3[51]), .B2(
        inst3_n2527), .ZN(inst3_n2505) );
  NAND2_X1 inst3_U779 ( .A1(inst3_n2503), .A2(inst3_n2502), .ZN(
        inst3_KeyArray_S21reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U778 ( .A1(inst3_n2543), .A2(inst3_n110), .B1(inst3_n70),
        .B2(inst3_n2662), .ZN(inst3_n2502) );
  AOI22_X1 inst3_U777 ( .A1(inst3_n94), .A2(inst3_n2552), .B1(key3[52]), .B2(
        inst3_n2506), .ZN(inst3_n2503) );
  NAND2_X1 inst3_U776 ( .A1(inst3_n2501), .A2(inst3_n2500), .ZN(
        inst3_KeyArray_S21reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst3_U775 ( .A1(inst3_n2543), .A2(inst3_n109), .B1(inst3_n2662),
        .B2(inst3_n69), .ZN(inst3_n2500) );
  AOI22_X1 inst3_U774 ( .A1(inst3_n93), .A2(inst3_n2552), .B1(key3[53]), .B2(
        inst3_n2527), .ZN(inst3_n2501) );
  NAND2_X1 inst3_U773 ( .A1(inst3_n2499), .A2(inst3_n2498), .ZN(
        inst3_KeyArray_S21reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst3_U772 ( .A1(inst3_n2543), .A2(inst3_n108), .B1(inst3_n2662),
        .B2(inst3_n68), .ZN(inst3_n2498) );
  AOI22_X1 inst3_U771 ( .A1(inst3_n92), .A2(inst3_n2552), .B1(key3[54]), .B2(
        inst3_n2506), .ZN(inst3_n2499) );
  NAND2_X1 inst3_U770 ( .A1(inst3_n2497), .A2(inst3_n2496), .ZN(
        inst3_KeyArray_S21reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst3_U769 ( .A1(inst3_n2543), .A2(inst3_n107), .B1(inst3_n2662),
        .B2(inst3_n67), .ZN(inst3_n2496) );
  AOI22_X1 inst3_U768 ( .A1(inst3_n91), .A2(inst3_n2552), .B1(key3[55]), .B2(
        inst3_n2506), .ZN(inst3_n2497) );
  OAI211_X1 inst3_U767 ( .C1(inst3_n1097), .C2(inst3_n2648), .A(inst3_n2495),
        .B(inst3_n2494), .ZN(inst3_KeyArray_S22reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst3_U766 ( .A1(inst3_n2487), .A2(inst3_n98), .ZN(inst3_n2494) );
  AOI22_X1 inst3_U765 ( .A1(inst3_n90), .A2(inst3_n2552), .B1(key3[40]), .B2(
        inst3_n2527), .ZN(inst3_n2495) );
  INV_X1 inst3_U764 ( .A(inst3_n6), .ZN(inst3_n2527) );
  NAND2_X1 inst3_U763 ( .A1(inst3_n2493), .A2(inst3_n2492), .ZN(
        inst3_KeyArray_S22reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U762 ( .A1(inst3_n2543), .A2(inst3_n97), .B1(inst3_n2662),
        .B2(inst3_n65), .ZN(inst3_n2492) );
  AOI22_X1 inst3_U761 ( .A1(inst3_n89), .A2(inst3_n2552), .B1(key3[41]), .B2(
        inst3_n2506), .ZN(inst3_n2493) );
  OAI211_X1 inst3_U760 ( .C1(inst3_n1095), .C2(inst3_n2648), .A(inst3_n2491),
        .B(inst3_n2490), .ZN(inst3_KeyArray_S22reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst3_U759 ( .A1(inst3_n2584), .A2(inst3_n96), .ZN(inst3_n2490) );
  AOI22_X1 inst3_U758 ( .A1(inst3_n88), .A2(inst3_n2552), .B1(key3[42]), .B2(
        inst3_n2506), .ZN(inst3_n2491) );
  OAI211_X1 inst3_U757 ( .C1(inst3_n1094), .C2(inst3_n2648), .A(inst3_n2489),
        .B(inst3_n2488), .ZN(inst3_KeyArray_S22reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst3_U756 ( .A1(inst3_n2487), .A2(inst3_n95), .ZN(inst3_n2488) );
  AOI22_X1 inst3_U755 ( .A1(inst3_n87), .A2(inst3_n2552), .B1(key3[43]), .B2(
        inst3_n2506), .ZN(inst3_n2489) );
  OAI211_X1 inst3_U754 ( .C1(inst3_n1093), .C2(inst3_n2648), .A(inst3_n2486),
        .B(inst3_n2485), .ZN(inst3_KeyArray_S22reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst3_U753 ( .A1(inst3_n2487), .A2(inst3_n94), .ZN(inst3_n2485) );
  AOI22_X1 inst3_U752 ( .A1(inst3_n86), .A2(inst3_n2552), .B1(key3[44]), .B2(
        inst3_n2506), .ZN(inst3_n2486) );
  OAI211_X1 inst3_U751 ( .C1(inst3_n1092), .C2(inst3_n2648), .A(inst3_n2484),
        .B(inst3_n2483), .ZN(inst3_KeyArray_S22reg_gff_1_SFF_5_n5) );
  NAND2_X1 inst3_U750 ( .A1(inst3_n2487), .A2(inst3_n93), .ZN(inst3_n2483) );
  AOI22_X1 inst3_U749 ( .A1(inst3_n85), .A2(inst3_n2552), .B1(key3[45]), .B2(
        inst3_n2527), .ZN(inst3_n2484) );
  OAI211_X1 inst3_U748 ( .C1(inst3_n1091), .C2(inst3_n2648), .A(inst3_n2482),
        .B(inst3_n2481), .ZN(inst3_KeyArray_S22reg_gff_1_SFF_6_n5) );
  NAND2_X1 inst3_U747 ( .A1(inst3_n2538), .A2(inst3_n92), .ZN(inst3_n2481) );
  AOI22_X1 inst3_U746 ( .A1(inst3_n84), .A2(inst3_n2613), .B1(key3[46]), .B2(
        inst3_n2506), .ZN(inst3_n2482) );
  OAI211_X1 inst3_U745 ( .C1(inst3_n1090), .C2(inst3_n2648), .A(inst3_n2480),
        .B(inst3_n2479), .ZN(inst3_KeyArray_S22reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst3_U744 ( .A1(inst3_n2487), .A2(inst3_n91), .ZN(inst3_n2479) );
  AOI22_X1 inst3_U743 ( .A1(inst3_n83), .A2(inst3_n2552), .B1(key3[47]), .B2(
        inst3_n2655), .ZN(inst3_n2480) );
  OAI211_X1 inst3_U742 ( .C1(inst3_n1089), .C2(inst3_n2648), .A(inst3_n2478),
        .B(inst3_n2477), .ZN(inst3_KeyArray_S23reg_gff_1_SFF_0_n5) );
  NAND2_X1 inst3_U741 ( .A1(inst3_n2543), .A2(inst3_n90), .ZN(inst3_n2477) );
  AOI22_X1 inst3_U740 ( .A1(inst3_n82), .A2(inst3_n2552), .B1(key3[32]), .B2(
        inst3_n2506), .ZN(inst3_n2478) );
  NAND2_X1 inst3_U739 ( .A1(inst3_n2476), .A2(inst3_n2475), .ZN(
        inst3_KeyArray_S23reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst3_U738 ( .A1(inst3_n2474), .A2(inst3_n89), .B1(inst3_n2662),
        .B2(inst3_n57), .ZN(inst3_n2475) );
  AOI22_X1 inst3_U737 ( .A1(inst3_n81), .A2(inst3_n2613), .B1(key3[33]), .B2(
        inst3_n2506), .ZN(inst3_n2476) );
  OAI211_X1 inst3_U736 ( .C1(inst3_n1087), .C2(inst3_n2648), .A(inst3_n2473),
        .B(inst3_n2472), .ZN(inst3_KeyArray_S23reg_gff_1_SFF_2_n5) );
  NAND2_X1 inst3_U735 ( .A1(inst3_n2487), .A2(inst3_n88), .ZN(inst3_n2472) );
  AOI22_X1 inst3_U734 ( .A1(inst3_n80), .A2(inst3_n2610), .B1(key3[34]), .B2(
        inst3_n2506), .ZN(inst3_n2473) );
  INV_X1 inst3_U733 ( .A(inst3_n6), .ZN(inst3_n2506) );
  OAI211_X1 inst3_U732 ( .C1(inst3_n1086), .C2(inst3_n2648), .A(inst3_n2471),
        .B(inst3_n2470), .ZN(inst3_KeyArray_S23reg_gff_1_SFF_3_n5) );
  NAND2_X1 inst3_U731 ( .A1(inst3_n2487), .A2(inst3_n87), .ZN(inst3_n2470) );
  AOI22_X1 inst3_U730 ( .A1(inst3_n79), .A2(inst3_n2555), .B1(key3[35]), .B2(
        inst3_n2655), .ZN(inst3_n2471) );
  OAI211_X1 inst3_U729 ( .C1(inst3_n1085), .C2(inst3_n2648), .A(inst3_n2469),
        .B(inst3_n2468), .ZN(inst3_KeyArray_S23reg_gff_1_SFF_4_n5) );
  NAND2_X1 inst3_U728 ( .A1(inst3_n2487), .A2(inst3_n86), .ZN(inst3_n2468) );
  AOI22_X1 inst3_U727 ( .A1(inst3_n2555), .A2(inst3_n78), .B1(key3[36]), .B2(
        inst3_n2727), .ZN(inst3_n2469) );
  OAI211_X1 inst3_U726 ( .C1(inst3_n1084), .C2(inst3_n2648), .A(inst3_n2467),
        .B(inst3_n2466), .ZN(inst3_KeyArray_S23reg_gff_1_SFF_5_n5) );
  NAND2_X1 inst3_U725 ( .A1(inst3_n2487), .A2(inst3_n85), .ZN(inst3_n2466) );
  AOI22_X1 inst3_U724 ( .A1(inst3_n77), .A2(inst3_n2610), .B1(key3[37]), .B2(
        inst3_n2655), .ZN(inst3_n2467) );
  OAI211_X1 inst3_U723 ( .C1(inst3_n1083), .C2(inst3_n2648), .A(inst3_n2465),
        .B(inst3_n2464), .ZN(inst3_KeyArray_S23reg_gff_1_SFF_6_n5) );
  NAND2_X1 inst3_U722 ( .A1(inst3_n2487), .A2(inst3_n84), .ZN(inst3_n2464) );
  AOI22_X1 inst3_U721 ( .A1(inst3_n76), .A2(inst3_n2613), .B1(key3[38]), .B2(
        inst3_n2774), .ZN(inst3_n2465) );
  OAI211_X1 inst3_U720 ( .C1(inst3_n1082), .C2(inst3_n2648), .A(inst3_n2463),
        .B(inst3_n2462), .ZN(inst3_KeyArray_S23reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst3_U719 ( .A1(inst3_n2487), .A2(inst3_n83), .ZN(inst3_n2462) );
  AOI22_X1 inst3_U718 ( .A1(inst3_n75), .A2(inst3_n2552), .B1(key3[39]), .B2(
        inst3_n2527), .ZN(inst3_n2463) );
  OAI211_X1 inst3_U717 ( .C1(inst3_n1097), .C2(inst3_n2461), .A(inst3_n2460),
        .B(inst3_n2459), .ZN(inst3_KeyArray_S31reg_gff_1_SFF_0_n6) );
  OR2_X1 inst3_U716 ( .A1(inst3_n2648), .A2(inst3_n1193), .ZN(inst3_n2459) );
  AOI22_X1 inst3_U715 ( .A1(inst3_n74), .A2(inst3_n2538), .B1(key3[16]), .B2(
        inst3_n2727), .ZN(inst3_n2460) );
  OAI211_X1 inst3_U714 ( .C1(inst3_n1192), .C2(inst3_n2648), .A(inst3_n2458),
        .B(inst3_n2457), .ZN(inst3_KeyArray_S31reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst3_U713 ( .A1(inst3_n2487), .A2(inst3_n73), .ZN(inst3_n2457) );
  AOI22_X1 inst3_U712 ( .A1(inst3_n65), .A2(inst3_n2555), .B1(key3[17]), .B2(
        inst3_n2506), .ZN(inst3_n2458) );
  OAI211_X1 inst3_U711 ( .C1(inst3_n1095), .C2(inst3_n2668), .A(inst3_n2456),
        .B(inst3_n2455), .ZN(inst3_KeyArray_S31reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst3_U710 ( .A1(inst3_n2665), .A2(inst3_n2828), .ZN(inst3_n2455)
         );
  AOI22_X1 inst3_U709 ( .A1(inst3_n72), .A2(inst3_n2474), .B1(key3[18]), .B2(
        inst3_n2727), .ZN(inst3_n2456) );
  OAI211_X1 inst3_U708 ( .C1(inst3_n1094), .C2(inst3_n2668), .A(inst3_n2454),
        .B(inst3_n2453), .ZN(inst3_KeyArray_S31reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst3_U707 ( .A1(inst3_n2665), .A2(inst3_n2827), .ZN(inst3_n2453)
         );
  AOI22_X1 inst3_U706 ( .A1(inst3_n71), .A2(inst3_n2543), .B1(key3[19]), .B2(
        inst3_n2655), .ZN(inst3_n2454) );
  OAI21_X1 inst3_U705 ( .B1(inst3_n1189), .B2(inst3_n2648), .A(inst3_n2452),
        .ZN(inst3_KeyArray_S31reg_gff_1_SFF_4_n6) );
  AOI21_X1 inst3_U704 ( .B1(key3[20]), .B2(inst3_n2593), .A(inst3_n2451), .ZN(
        inst3_n2452) );
  OAI22_X1 inst3_U703 ( .A1(inst3_n1093), .A2(inst3_n2461), .B1(inst3_n2799),
        .B2(inst3_n2837), .ZN(inst3_n2451) );
  OAI211_X1 inst3_U702 ( .C1(inst3_n1092), .C2(inst3_n2668), .A(inst3_n2450),
        .B(inst3_n2449), .ZN(inst3_KeyArray_S31reg_gff_1_SFF_5_n6) );
  NAND2_X1 inst3_U701 ( .A1(inst3_n2665), .A2(inst3_n2826), .ZN(inst3_n2449)
         );
  AOI22_X1 inst3_U700 ( .A1(inst3_n69), .A2(inst3_n2584), .B1(key3[21]), .B2(
        inst3_n2727), .ZN(inst3_n2450) );
  OAI211_X1 inst3_U699 ( .C1(inst3_n1091), .C2(inst3_n2668), .A(inst3_n2448),
        .B(inst3_n2447), .ZN(inst3_KeyArray_S31reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst3_U698 ( .A1(inst3_n2662), .A2(inst3_n2825), .ZN(inst3_n2447)
         );
  AOI22_X1 inst3_U697 ( .A1(inst3_n68), .A2(inst3_n2538), .B1(key3[22]), .B2(
        inst3_n2774), .ZN(inst3_n2448) );
  OAI211_X1 inst3_U696 ( .C1(inst3_n1090), .C2(inst3_n2668), .A(inst3_n2446),
        .B(inst3_n2445), .ZN(inst3_KeyArray_S31reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst3_U695 ( .A1(inst3_n2665), .A2(inst3_n2824), .ZN(inst3_n2445)
         );
  AOI22_X1 inst3_U694 ( .A1(inst3_n67), .A2(inst3_n2584), .B1(key3[23]), .B2(
        inst3_n2727), .ZN(inst3_n2446) );
  OAI211_X1 inst3_U693 ( .C1(inst3_n1184), .C2(inst3_n2648), .A(inst3_n2444),
        .B(inst3_n2443), .ZN(inst3_KeyArray_S32reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst3_U692 ( .A1(inst3_n2487), .A2(inst3_n65), .ZN(inst3_n2443) );
  AOI22_X1 inst3_U691 ( .A1(inst3_n57), .A2(inst3_n2610), .B1(key3[9]), .B2(
        inst3_n2713), .ZN(inst3_n2444) );
  OAI21_X1 inst3_U690 ( .B1(inst3_n1265), .B2(inst3_n2442), .A(inst3_n2441),
        .ZN(inst3_stateArray_S10reg_gff_1_SFF_0_n5) );
  AOI22_X1 inst3_U689 ( .A1(inst3_n2756), .A2(ciphertext3[88]), .B1(
        plaintext3[88]), .B2(inst3_n2710), .ZN(inst3_n2441) );
  OAI21_X1 inst3_U688 ( .B1(inst3_n1264), .B2(inst3_n2442), .A(inst3_n2440),
        .ZN(inst3_stateArray_S10reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst3_U687 ( .A1(inst3_n2756), .A2(ciphertext3[89]), .B1(
        plaintext3[89]), .B2(inst3_n2710), .ZN(inst3_n2440) );
  OAI21_X1 inst3_U686 ( .B1(inst3_n1263), .B2(inst3_n2442), .A(inst3_n2439),
        .ZN(inst3_stateArray_S10reg_gff_1_SFF_2_n5) );
  AOI22_X1 inst3_U685 ( .A1(done3), .A2(ciphertext3[90]), .B1(plaintext3[90]),
        .B2(inst3_n2527), .ZN(inst3_n2439) );
  OAI21_X1 inst3_U684 ( .B1(inst3_n1262), .B2(inst3_n2442), .A(inst3_n2438),
        .ZN(inst3_stateArray_S10reg_gff_1_SFF_3_n5) );
  AOI22_X1 inst3_U683 ( .A1(inst3_n2756), .A2(ciphertext3[91]), .B1(
        plaintext3[91]), .B2(inst3_n2713), .ZN(inst3_n2438) );
  OAI21_X1 inst3_U682 ( .B1(inst3_n1261), .B2(inst3_n2442), .A(inst3_n2437),
        .ZN(inst3_stateArray_S10reg_gff_1_SFF_4_n5) );
  AOI22_X1 inst3_U681 ( .A1(done3), .A2(ciphertext3[92]), .B1(plaintext3[92]),
        .B2(inst3_n2506), .ZN(inst3_n2437) );
  OAI21_X1 inst3_U680 ( .B1(inst3_n1260), .B2(inst3_n2442), .A(inst3_n2436),
        .ZN(inst3_stateArray_S10reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst3_U679 ( .A1(inst3_n2756), .A2(ciphertext3[93]), .B1(
        plaintext3[93]), .B2(inst3_n2727), .ZN(inst3_n2436) );
  OAI21_X1 inst3_U678 ( .B1(inst3_n1259), .B2(inst3_n2442), .A(inst3_n2435),
        .ZN(inst3_stateArray_S10reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst3_U677 ( .A1(inst3_n1914), .A2(ciphertext3[94]), .B1(
        plaintext3[94]), .B2(inst3_n2713), .ZN(inst3_n2435) );
  OAI21_X1 inst3_U676 ( .B1(inst3_n1258), .B2(inst3_n2442), .A(inst3_n2434),
        .ZN(inst3_stateArray_S10reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst3_U675 ( .A1(inst3_n1914), .A2(ciphertext3[95]), .B1(
        plaintext3[95]), .B2(inst3_n2655), .ZN(inst3_n2434) );
  INV_X1 inst3_U674 ( .A(inst3_n2433), .ZN(inst3_n2442) );
  OAI21_X1 inst3_U673 ( .B1(inst3_n1265), .B2(inst3_n2708), .A(inst3_n2432),
        .ZN(inst3_stateArray_S11reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst3_U672 ( .A1(inst3_n2433), .A2(ciphertext3[72]), .B1(
        plaintext3[80]), .B2(inst3_n2527), .ZN(inst3_n2432) );
  OAI21_X1 inst3_U671 ( .B1(inst3_n1264), .B2(inst3_n2708), .A(inst3_n2431),
        .ZN(inst3_stateArray_S11reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U670 ( .A1(inst3_n2433), .A2(ciphertext3[73]), .B1(
        plaintext3[81]), .B2(inst3_n2713), .ZN(inst3_n2431) );
  OAI21_X1 inst3_U669 ( .B1(inst3_n1263), .B2(inst3_n2708), .A(inst3_n2430),
        .ZN(inst3_stateArray_S11reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U668 ( .A1(inst3_n2433), .A2(ciphertext3[74]), .B1(
        plaintext3[82]), .B2(inst3_n2710), .ZN(inst3_n2430) );
  OAI21_X1 inst3_U667 ( .B1(inst3_n1262), .B2(inst3_n2708), .A(inst3_n2429),
        .ZN(inst3_stateArray_S11reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U666 ( .A1(inst3_n2433), .A2(ciphertext3[75]), .B1(
        plaintext3[83]), .B2(inst3_n2527), .ZN(inst3_n2429) );
  OAI21_X1 inst3_U665 ( .B1(inst3_n1250), .B2(inst3_n2708), .A(inst3_n2428),
        .ZN(inst3_stateArray_S12reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst3_U664 ( .A1(inst3_n2433), .A2(ciphertext3[71]), .B1(
        plaintext3[79]), .B2(inst3_n2713), .ZN(inst3_n2428) );
  OAI21_X1 inst3_U663 ( .B1(inst3_n1261), .B2(inst3_n2708), .A(inst3_n2427),
        .ZN(inst3_stateArray_S11reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U662 ( .A1(inst3_n2433), .A2(ciphertext3[76]), .B1(
        plaintext3[84]), .B2(inst3_n2774), .ZN(inst3_n2427) );
  OAI21_X1 inst3_U661 ( .B1(inst3_n1260), .B2(inst3_n2708), .A(inst3_n2426),
        .ZN(inst3_stateArray_S11reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst3_U660 ( .A1(inst3_n2433), .A2(ciphertext3[77]), .B1(
        plaintext3[85]), .B2(inst3_n2713), .ZN(inst3_n2426) );
  OAI21_X1 inst3_U659 ( .B1(inst3_n1259), .B2(inst3_n2708), .A(inst3_n2425),
        .ZN(inst3_stateArray_S11reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst3_U658 ( .A1(inst3_n2433), .A2(ciphertext3[78]), .B1(
        plaintext3[86]), .B2(inst3_n2506), .ZN(inst3_n2425) );
  OAI21_X1 inst3_U657 ( .B1(inst3_n1258), .B2(inst3_n2708), .A(inst3_n2424),
        .ZN(inst3_stateArray_S11reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst3_U656 ( .A1(inst3_n2433), .A2(ciphertext3[79]), .B1(
        plaintext3[87]), .B2(inst3_n2727), .ZN(inst3_n2424) );
  OAI21_X1 inst3_U655 ( .B1(inst3_n1257), .B2(inst3_n2708), .A(inst3_n2423),
        .ZN(inst3_stateArray_S12reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst3_U654 ( .A1(inst3_n2433), .A2(ciphertext3[64]), .B1(
        plaintext3[72]), .B2(inst3_n2710), .ZN(inst3_n2423) );
  OAI21_X1 inst3_U653 ( .B1(inst3_n1256), .B2(inst3_n2708), .A(inst3_n2422),
        .ZN(inst3_stateArray_S12reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U652 ( .A1(inst3_n2433), .A2(ciphertext3[65]), .B1(
        plaintext3[73]), .B2(inst3_n2774), .ZN(inst3_n2422) );
  OAI21_X1 inst3_U651 ( .B1(inst3_n1255), .B2(inst3_n2708), .A(inst3_n2421),
        .ZN(inst3_stateArray_S12reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U650 ( .A1(inst3_n2433), .A2(ciphertext3[66]), .B1(
        plaintext3[74]), .B2(inst3_n2727), .ZN(inst3_n2421) );
  OAI21_X1 inst3_U649 ( .B1(inst3_n1254), .B2(inst3_n2708), .A(inst3_n2420),
        .ZN(inst3_stateArray_S12reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U648 ( .A1(inst3_n2433), .A2(ciphertext3[67]), .B1(
        plaintext3[75]), .B2(inst3_n2713), .ZN(inst3_n2420) );
  OAI21_X1 inst3_U647 ( .B1(inst3_n1253), .B2(inst3_n2708), .A(inst3_n2419),
        .ZN(inst3_stateArray_S12reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U646 ( .A1(inst3_n2433), .A2(ciphertext3[68]), .B1(
        plaintext3[76]), .B2(inst3_n2655), .ZN(inst3_n2419) );
  OAI21_X1 inst3_U645 ( .B1(inst3_n1252), .B2(inst3_n2708), .A(inst3_n2418),
        .ZN(inst3_stateArray_S12reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst3_U644 ( .A1(inst3_n2433), .A2(ciphertext3[69]), .B1(
        plaintext3[77]), .B2(inst3_n2710), .ZN(inst3_n2418) );
  OAI21_X1 inst3_U643 ( .B1(inst3_n1251), .B2(inst3_n2708), .A(inst3_n2417),
        .ZN(inst3_stateArray_S12reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst3_U642 ( .A1(inst3_n2433), .A2(ciphertext3[70]), .B1(
        plaintext3[78]), .B2(inst3_n2506), .ZN(inst3_n2417) );
  NOR2_X2 inst3_U641 ( .A1(inst3_n2756), .A2(inst3_n2774), .ZN(inst3_n2433) );
  OAI211_X1 inst3_U640 ( .C1(inst3_n1176), .C2(inst3_n2648), .A(inst3_n2416),
        .B(inst3_n2415), .ZN(inst3_KeyArray_S33reg_gff_1_SFF_1_n5) );
  NAND2_X1 inst3_U639 ( .A1(inst3_n2487), .A2(inst3_n57), .ZN(inst3_n2415) );
  INV_X1 inst3_U638 ( .A(inst3_n2799), .ZN(inst3_n2487) );
  AOI22_X1 inst3_U637 ( .A1(inst3_n2610), .A2(inst3_n2814), .B1(key3[1]), .B2(
        inst3_n2727), .ZN(inst3_n2416) );
  OAI21_X1 inst3_U636 ( .B1(inst3_n1175), .B2(inst3_n2648), .A(inst3_n2414),
        .ZN(inst3_KeyArray_S33reg_gff_1_SFF_2_n5) );
  AOI21_X1 inst3_U635 ( .B1(key3[2]), .B2(inst3_n2727), .A(inst3_n2413), .ZN(
        inst3_n2414) );
  OAI22_X1 inst3_U634 ( .A1(inst3_n225), .A2(inst3_n2461), .B1(inst3_n1087),
        .B2(inst3_n2799), .ZN(inst3_n2413) );
  OAI21_X1 inst3_U633 ( .B1(inst3_n1174), .B2(inst3_n2648), .A(inst3_n2412),
        .ZN(inst3_KeyArray_S33reg_gff_1_SFF_3_n5) );
  AOI21_X1 inst3_U632 ( .B1(key3[3]), .B2(inst3_n2713), .A(inst3_n2411), .ZN(
        inst3_n2412) );
  OAI22_X1 inst3_U631 ( .A1(inst3_n224), .A2(inst3_n2461), .B1(inst3_n1086),
        .B2(inst3_n2799), .ZN(inst3_n2411) );
  OAI211_X1 inst3_U630 ( .C1(inst3_n1203), .C2(inst3_n2775), .A(inst3_n2410),
        .B(inst3_n2409), .ZN(inst3_stateArray_S31reg_gff_1_SFF_6_n6) );
  NAND2_X1 inst3_U629 ( .A1(plaintext3[22]), .A2(inst3_n2727), .ZN(inst3_n2409) );
  AOI22_X1 inst3_U628 ( .A1(ciphertext3[22]), .A2(inst3_n2750), .B1(
        inst3_n2794), .B2(ciphertext3[30]), .ZN(inst3_n2410) );
  OAI211_X1 inst3_U627 ( .C1(inst3_n1202), .C2(inst3_n2775), .A(inst3_n2408),
        .B(inst3_n2407), .ZN(inst3_stateArray_S31reg_gff_1_SFF_7_n6) );
  NAND2_X1 inst3_U626 ( .A1(plaintext3[23]), .A2(inst3_n2774), .ZN(inst3_n2407) );
  AOI22_X1 inst3_U625 ( .A1(done3), .A2(ciphertext3[23]), .B1(inst3_n2794),
        .B2(ciphertext3[31]), .ZN(inst3_n2408) );
  OAI21_X1 inst3_U624 ( .B1(inst3_n1220), .B2(inst3_n2775), .A(inst3_n2406),
        .ZN(inst3_stateArray_S22reg_gff_1_SFF_5_n6) );
  AOI21_X1 inst3_U623 ( .B1(plaintext3[45]), .B2(inst3_n2713), .A(inst3_n2405),
        .ZN(inst3_n2406) );
  OAI22_X1 inst3_U622 ( .A1(inst3_n1228), .A2(inst3_n2708), .B1(inst3_n2760),
        .B2(inst3_n2823), .ZN(inst3_n2405) );
  OAI21_X1 inst3_U621 ( .B1(inst3_n1177), .B2(inst3_n2648), .A(inst3_n2404),
        .ZN(inst3_KeyArray_S33reg_gff_1_SFF_0_n5) );
  AOI21_X1 inst3_U620 ( .B1(key3[0]), .B2(inst3_n2710), .A(inst3_n2403), .ZN(
        inst3_n2404) );
  OAI22_X1 inst3_U619 ( .A1(inst3_n227), .A2(inst3_n2461), .B1(inst3_n1089),
        .B2(inst3_n2799), .ZN(inst3_n2403) );
  OAI21_X1 inst3_U618 ( .B1(inst3_n1173), .B2(inst3_n2648), .A(inst3_n2402),
        .ZN(inst3_KeyArray_S33reg_gff_1_SFF_4_n5) );
  AOI21_X1 inst3_U617 ( .B1(key3[4]), .B2(inst3_n2713), .A(inst3_n2401), .ZN(
        inst3_n2402) );
  OAI22_X1 inst3_U616 ( .A1(inst3_n223), .A2(inst3_n2461), .B1(inst3_n1085),
        .B2(inst3_n2799), .ZN(inst3_n2401) );
  OAI21_X1 inst3_U615 ( .B1(inst3_n1172), .B2(inst3_n2648), .A(inst3_n2400),
        .ZN(inst3_KeyArray_S33reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst3_U614 ( .B1(key3[5]), .B2(inst3_n2593), .A(inst3_n2399), .ZN(
        inst3_n2400) );
  OAI22_X1 inst3_U613 ( .A1(inst3_n228), .A2(inst3_n2461), .B1(inst3_n1084),
        .B2(inst3_n2799), .ZN(inst3_n2399) );
  OAI21_X1 inst3_U612 ( .B1(inst3_n1171), .B2(inst3_n2648), .A(inst3_n2398),
        .ZN(inst3_KeyArray_S33reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst3_U611 ( .B1(key3[6]), .B2(inst3_n2713), .A(inst3_n2397), .ZN(
        inst3_n2398) );
  OAI22_X1 inst3_U610 ( .A1(inst3_n222), .A2(inst3_n2461), .B1(inst3_n1083),
        .B2(inst3_n2799), .ZN(inst3_n2397) );
  OAI21_X1 inst3_U609 ( .B1(inst3_n1170), .B2(inst3_n2648), .A(inst3_n2396),
        .ZN(inst3_KeyArray_S33reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst3_U608 ( .B1(key3[7]), .B2(inst3_n2713), .A(inst3_n2395), .ZN(
        inst3_n2396) );
  OAI22_X1 inst3_U607 ( .A1(inst3_n221), .A2(inst3_n2461), .B1(inst3_n1082),
        .B2(inst3_n2799), .ZN(inst3_n2395) );
  OAI211_X1 inst3_U606 ( .C1(inst3_n210), .C2(inst3_n2792), .A(inst3_n2394),
        .B(inst3_n2393), .ZN(inst3_stateArray_S03reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst3_U605 ( .A1(inst3_n2555), .A2(ciphertext3[88]), .B1(
        inst3_n2392), .B2(inst3_n2391), .ZN(inst3_n2393) );
  XNOR2_X1 inst3_U604 ( .A(inst3_n2786), .B(inst3_n2390), .ZN(inst3_n2391) );
  AOI22_X1 inst3_U603 ( .A1(inst3_n2389), .A2(ciphertext3[88]), .B1(inst3_n209), .B2(inst3_n2388), .ZN(inst3_n2390) );
  AOI22_X1 inst3_U602 ( .A1(inst3_n2474), .A2(ciphertext3[96]), .B1(
        plaintext3[96]), .B2(inst3_n2713), .ZN(inst3_n2394) );
  OAI211_X1 inst3_U601 ( .C1(inst3_n1169), .C2(inst3_n2648), .A(inst3_n2387),
        .B(inst3_n2386), .ZN(inst3_KeyArray_S00reg_gff_1_SFF_0_n6) );
  OAI21_X1 inst3_U600 ( .B1(inst3_n1193), .B2(inst3_n2385), .A(inst3_n2384),
        .ZN(inst3_n2386) );
  AOI21_X1 inst3_U599 ( .B1(inst3_n1193), .B2(inst3_n2385), .A(inst3_n2780),
        .ZN(inst3_n2384) );
  NAND2_X1 inst3_U598 ( .A1(inst3_n2383), .A2(inst3_n2820), .ZN(inst3_n2385)
         );
  AOI22_X1 inst3_U597 ( .A1(inst3_n2474), .A2(inst3_n2820), .B1(key3[120]),
        .B2(inst3_n2713), .ZN(inst3_n2387) );
  OAI211_X1 inst3_U596 ( .C1(inst3_n1168), .C2(inst3_n2648), .A(inst3_n2382),
        .B(inst3_n2381), .ZN(inst3_KeyArray_S00reg_gff_1_SFF_1_n6) );
  OAI21_X1 inst3_U595 ( .B1(inst3_n1192), .B2(inst3_n2380), .A(inst3_n2379),
        .ZN(inst3_n2381) );
  AOI21_X1 inst3_U594 ( .B1(inst3_n1192), .B2(inst3_n2380), .A(inst3_n2780),
        .ZN(inst3_n2379) );
  NAND2_X1 inst3_U593 ( .A1(inst3_n2383), .A2(inst3_n2814), .ZN(inst3_n2380)
         );
  AOI22_X1 inst3_U592 ( .A1(inst3_n2474), .A2(inst3_n2814), .B1(key3[121]),
        .B2(inst3_n2506), .ZN(inst3_n2382) );
  OAI211_X1 inst3_U591 ( .C1(inst3_n1167), .C2(inst3_n2648), .A(inst3_n2378),
        .B(inst3_n2377), .ZN(inst3_KeyArray_S00reg_gff_1_SFF_2_n6) );
  OAI21_X1 inst3_U590 ( .B1(inst3_n1191), .B2(inst3_n2376), .A(inst3_n2375),
        .ZN(inst3_n2377) );
  AOI21_X1 inst3_U589 ( .B1(inst3_n1191), .B2(inst3_n2376), .A(inst3_n2780),
        .ZN(inst3_n2375) );
  INV_X1 inst3_U588 ( .A(inst3_n2555), .ZN(inst3_n2780) );
  NAND2_X1 inst3_U587 ( .A1(inst3_n2383), .A2(inst3_n2815), .ZN(inst3_n2376)
         );
  AOI22_X1 inst3_U586 ( .A1(inst3_n2474), .A2(inst3_n2815), .B1(key3[122]),
        .B2(inst3_n2806), .ZN(inst3_n2378) );
  OAI211_X1 inst3_U585 ( .C1(inst3_n1166), .C2(inst3_n2648), .A(inst3_n2374),
        .B(inst3_n2373), .ZN(inst3_KeyArray_S00reg_gff_1_SFF_3_n6) );
  OAI21_X1 inst3_U584 ( .B1(inst3_n1190), .B2(inst3_n2372), .A(inst3_n2371),
        .ZN(inst3_n2373) );
  AOI21_X1 inst3_U583 ( .B1(inst3_n1190), .B2(inst3_n2372), .A(inst3_n2461),
        .ZN(inst3_n2371) );
  NAND2_X1 inst3_U582 ( .A1(inst3_n2383), .A2(inst3_n2819), .ZN(inst3_n2372)
         );
  AOI22_X1 inst3_U581 ( .A1(inst3_n2474), .A2(inst3_n2819), .B1(key3[123]),
        .B2(inst3_n2806), .ZN(inst3_n2374) );
  OAI211_X1 inst3_U580 ( .C1(inst3_n1165), .C2(inst3_n2648), .A(inst3_n2370),
        .B(inst3_n2369), .ZN(inst3_KeyArray_S00reg_gff_1_SFF_4_n6) );
  OAI21_X1 inst3_U579 ( .B1(inst3_n1189), .B2(inst3_n2368), .A(inst3_n2367),
        .ZN(inst3_n2369) );
  AOI21_X1 inst3_U578 ( .B1(inst3_n1189), .B2(inst3_n2368), .A(inst3_n2461),
        .ZN(inst3_n2367) );
  NAND2_X1 inst3_U577 ( .A1(inst3_n2383), .A2(inst3_n2818), .ZN(inst3_n2368)
         );
  AOI22_X1 inst3_U576 ( .A1(inst3_n2543), .A2(inst3_n2818), .B1(key3[124]),
        .B2(inst3_n2806), .ZN(inst3_n2370) );
  INV_X1 inst3_U575 ( .A(inst3_n2799), .ZN(inst3_n2543) );
  OAI211_X1 inst3_U574 ( .C1(inst3_n1164), .C2(inst3_n2648), .A(inst3_n2366),
        .B(inst3_n2365), .ZN(inst3_KeyArray_S00reg_gff_1_SFF_5_n6) );
  OAI21_X1 inst3_U573 ( .B1(inst3_n1188), .B2(inst3_n2364), .A(inst3_n2363),
        .ZN(inst3_n2365) );
  AOI21_X1 inst3_U572 ( .B1(inst3_n1188), .B2(inst3_n2364), .A(inst3_n2461),
        .ZN(inst3_n2363) );
  NAND2_X1 inst3_U571 ( .A1(inst3_n2383), .A2(inst3_n2817), .ZN(inst3_n2364)
         );
  AOI22_X1 inst3_U570 ( .A1(inst3_n2474), .A2(inst3_n2817), .B1(key3[125]),
        .B2(inst3_n2806), .ZN(inst3_n2366) );
  OAI211_X1 inst3_U569 ( .C1(inst3_n1163), .C2(inst3_n2648), .A(inst3_n2362),
        .B(inst3_n2361), .ZN(inst3_KeyArray_S00reg_gff_1_SFF_6_n6) );
  OAI21_X1 inst3_U568 ( .B1(inst3_n1187), .B2(inst3_n2360), .A(inst3_n2359),
        .ZN(inst3_n2361) );
  AOI21_X1 inst3_U567 ( .B1(inst3_n1187), .B2(inst3_n2360), .A(inst3_n2780),
        .ZN(inst3_n2359) );
  NAND2_X1 inst3_U566 ( .A1(inst3_n2383), .A2(inst3_n2816), .ZN(inst3_n2360)
         );
  AOI22_X1 inst3_U565 ( .A1(inst3_n2474), .A2(inst3_n2816), .B1(key3[126]),
        .B2(inst3_n2806), .ZN(inst3_n2362) );
  OAI211_X1 inst3_U564 ( .C1(inst3_n1162), .C2(inst3_n2648), .A(inst3_n2358),
        .B(inst3_n2357), .ZN(inst3_KeyArray_S00reg_gff_1_SFF_7_n6) );
  OAI21_X1 inst3_U563 ( .B1(inst3_n1186), .B2(inst3_n2356), .A(inst3_n2355),
        .ZN(inst3_n2357) );
  AOI21_X1 inst3_U562 ( .B1(inst3_n1186), .B2(inst3_n2356), .A(inst3_n2780),
        .ZN(inst3_n2355) );
  NAND2_X1 inst3_U561 ( .A1(inst3_n2383), .A2(inst3_n2804), .ZN(inst3_n2356)
         );
  AOI21_X1 inst3_U560 ( .B1(inst3_n2354), .B2(inst3_n2353), .A(inst3_n2801),
        .ZN(inst3_n2383) );
  NOR2_X1 inst3_U559 ( .A1(inst3_n143), .A2(inst3_n25), .ZN(inst3_n2801) );
  AND4_X1 inst3_U558 ( .A1(inst3_n2838), .A2(inst3_n499), .A3(inst3_n1081),
        .A4(inst3_n1080), .ZN(inst3_n2353) );
  AND4_X1 inst3_U557 ( .A1(inst3_n2803), .A2(inst3_n2813), .A3(inst3_n2839),
        .A4(inst3_n718), .ZN(inst3_n2354) );
  AOI22_X1 inst3_U556 ( .A1(inst3_n2474), .A2(inst3_n2804), .B1(key3[127]),
        .B2(inst3_n2806), .ZN(inst3_n2358) );
  INV_X4 inst3_U555 ( .A(inst3_n2662), .ZN(inst3_n2648) );
  OAI211_X1 inst3_U554 ( .C1(inst3_n1206), .C2(inst3_n2775), .A(inst3_n2352),
        .B(inst3_n2351), .ZN(inst3_stateArray_S31reg_gff_1_SFF_3_n6) );
  NAND2_X1 inst3_U553 ( .A1(plaintext3[19]), .A2(inst3_n2727), .ZN(inst3_n2351) );
  AOI22_X1 inst3_U552 ( .A1(done3), .A2(ciphertext3[19]), .B1(inst3_n2794),
        .B2(ciphertext3[27]), .ZN(inst3_n2352) );
  OAI211_X1 inst3_U551 ( .C1(inst3_n198), .C2(inst3_n2792), .A(inst3_n2350),
        .B(inst3_n2349), .ZN(inst3_stateArray_S03reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U550 ( .A1(inst3_n2610), .A2(ciphertext3[89]), .B1(
        inst3_n2392), .B2(inst3_n2348), .ZN(inst3_n2349) );
  XNOR2_X1 inst3_U549 ( .A(inst3_n2347), .B(inst3_n2346), .ZN(inst3_n2348) );
  AOI22_X1 inst3_U548 ( .A1(inst3_n2389), .A2(ciphertext3[89]), .B1(inst3_n197), .B2(inst3_n2388), .ZN(inst3_n2346) );
  AOI22_X1 inst3_U547 ( .A1(inst3_n2345), .A2(inst3_n2776), .B1(inst3_n2777),
        .B2(inst3_n2344), .ZN(inst3_n2347) );
  INV_X1 inst3_U546 ( .A(inst3_n2345), .ZN(inst3_n2344) );
  INV_X1 inst3_U545 ( .A(inst3_n2776), .ZN(inst3_n2777) );
  AOI22_X1 inst3_U544 ( .A1(inst3_n2474), .A2(ciphertext3[97]), .B1(
        plaintext3[97]), .B2(inst3_n2806), .ZN(inst3_n2350) );
  OAI211_X1 inst3_U543 ( .C1(inst3_n202), .C2(inst3_n2792), .A(inst3_n2343),
        .B(inst3_n2342), .ZN(inst3_stateArray_S03reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U542 ( .A1(inst3_n2555), .A2(ciphertext3[91]), .B1(
        inst3_n2392), .B2(inst3_n2341), .ZN(inst3_n2342) );
  XNOR2_X1 inst3_U541 ( .A(inst3_n2340), .B(inst3_n2339), .ZN(inst3_n2341) );
  AOI22_X1 inst3_U540 ( .A1(inst3_n201), .A2(inst3_n2389), .B1(inst3_n2388),
        .B2(ciphertext3[91]), .ZN(inst3_n2339) );
  AOI22_X1 inst3_U539 ( .A1(inst3_n2779), .A2(inst3_n2765), .B1(inst3_n2764),
        .B2(inst3_n2338), .ZN(inst3_n2340) );
  INV_X1 inst3_U538 ( .A(inst3_n2779), .ZN(inst3_n2338) );
  INV_X1 inst3_U537 ( .A(inst3_n2765), .ZN(inst3_n2764) );
  AOI22_X1 inst3_U536 ( .A1(inst3_n2487), .A2(ciphertext3[99]), .B1(
        plaintext3[99]), .B2(inst3_n2806), .ZN(inst3_n2343) );
  OAI211_X1 inst3_U535 ( .C1(inst3_n216), .C2(inst3_n2792), .A(inst3_n2337),
        .B(inst3_n2336), .ZN(inst3_stateArray_S03reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst3_U534 ( .A1(inst3_n2610), .A2(ciphertext3[94]), .B1(
        inst3_n2392), .B2(inst3_n2335), .ZN(inst3_n2336) );
  XNOR2_X1 inst3_U533 ( .A(inst3_n2334), .B(inst3_n2333), .ZN(inst3_n2335) );
  AOI22_X1 inst3_U532 ( .A1(inst3_n214), .A2(ciphertext3[30]), .B1(inst3_n215),
        .B2(ciphertext3[125]), .ZN(inst3_n2333) );
  AOI22_X1 inst3_U531 ( .A1(inst3_n2332), .A2(inst3_n190), .B1(ciphertext3[93]), .B2(inst3_n2331), .ZN(inst3_n2334) );
  INV_X1 inst3_U530 ( .A(inst3_n2332), .ZN(inst3_n2331) );
  AOI22_X1 inst3_U529 ( .A1(inst3_n2474), .A2(ciphertext3[102]), .B1(
        plaintext3[102]), .B2(inst3_n2806), .ZN(inst3_n2337) );
  OAI211_X1 inst3_U528 ( .C1(inst3_n2805), .C2(inst3_n2792), .A(inst3_n2330),
        .B(inst3_n2329), .ZN(inst3_stateArray_S03reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U527 ( .A1(inst3_n2610), .A2(ciphertext3[90]), .B1(
        inst3_n2392), .B2(inst3_n2328), .ZN(inst3_n2329) );
  XNOR2_X1 inst3_U526 ( .A(inst3_n2327), .B(inst3_n2326), .ZN(inst3_n2328) );
  AOI22_X1 inst3_U525 ( .A1(inst3_n203), .A2(inst3_n2787), .B1(inst3_n2325),
        .B2(ciphertext3[26]), .ZN(inst3_n2326) );
  INV_X1 inst3_U524 ( .A(inst3_n2787), .ZN(inst3_n2325) );
  AOI22_X1 inst3_U523 ( .A1(inst3_n2543), .A2(ciphertext3[98]), .B1(
        plaintext3[98]), .B2(inst3_n2806), .ZN(inst3_n2330) );
  OAI211_X1 inst3_U522 ( .C1(inst3_n214), .C2(inst3_n2792), .A(inst3_n2324),
        .B(inst3_n2323), .ZN(inst3_stateArray_S03reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst3_U521 ( .A1(inst3_n2610), .A2(ciphertext3[93]), .B1(
        inst3_n2392), .B2(inst3_n2322), .ZN(inst3_n2323) );
  XNOR2_X1 inst3_U520 ( .A(inst3_n2321), .B(inst3_n2320), .ZN(inst3_n2322) );
  AOI22_X1 inst3_U519 ( .A1(ciphertext3[124]), .A2(inst3_n2807), .B1(
        ciphertext3[29]), .B2(inst3_n2802), .ZN(inst3_n2320) );
  AOI22_X1 inst3_U518 ( .A1(inst3_n212), .A2(inst3_n2319), .B1(inst3_n2318),
        .B2(ciphertext3[92]), .ZN(inst3_n2321) );
  INV_X1 inst3_U517 ( .A(inst3_n2319), .ZN(inst3_n2318) );
  AOI22_X1 inst3_U516 ( .A1(inst3_n2474), .A2(ciphertext3[101]), .B1(
        plaintext3[101]), .B2(inst3_n2806), .ZN(inst3_n2324) );
  OAI211_X1 inst3_U515 ( .C1(inst3_n2802), .C2(inst3_n2792), .A(inst3_n2317),
        .B(inst3_n2316), .ZN(inst3_stateArray_S03reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U514 ( .A1(inst3_n2555), .A2(ciphertext3[92]), .B1(
        inst3_n2392), .B2(inst3_n2315), .ZN(inst3_n2316) );
  XNOR2_X1 inst3_U513 ( .A(inst3_n2314), .B(inst3_n2313), .ZN(inst3_n2315) );
  AOI22_X1 inst3_U512 ( .A1(inst3_n207), .A2(inst3_n2312), .B1(inst3_n2311),
        .B2(ciphertext3[28]), .ZN(inst3_n2313) );
  INV_X1 inst3_U511 ( .A(inst3_n2311), .ZN(inst3_n2312) );
  AOI22_X1 inst3_U510 ( .A1(inst3_n2310), .A2(inst3_n2389), .B1(inst3_n2388),
        .B2(inst3_n2309), .ZN(inst3_n2314) );
  AOI22_X1 inst3_U509 ( .A1(inst3_n2487), .A2(ciphertext3[100]), .B1(
        plaintext3[100]), .B2(inst3_n2713), .ZN(inst3_n2317) );
  OAI211_X1 inst3_U508 ( .C1(inst3_n1208), .C2(inst3_n2775), .A(inst3_n2308),
        .B(inst3_n2307), .ZN(inst3_stateArray_S31reg_gff_1_SFF_1_n6) );
  NAND2_X1 inst3_U507 ( .A1(plaintext3[17]), .A2(inst3_n2727), .ZN(inst3_n2307) );
  AOI22_X1 inst3_U506 ( .A1(done3), .A2(ciphertext3[17]), .B1(inst3_n2794),
        .B2(ciphertext3[25]), .ZN(inst3_n2308) );
  OAI211_X1 inst3_U505 ( .C1(inst3_n1209), .C2(inst3_n2775), .A(inst3_n2306),
        .B(inst3_n2305), .ZN(inst3_stateArray_S31reg_gff_1_SFF_0_n6) );
  NAND2_X1 inst3_U504 ( .A1(plaintext3[16]), .A2(inst3_n2727), .ZN(inst3_n2305) );
  AOI22_X1 inst3_U503 ( .A1(done3), .A2(ciphertext3[16]), .B1(inst3_n2794),
        .B2(ciphertext3[24]), .ZN(inst3_n2306) );
  OAI211_X1 inst3_U502 ( .C1(inst3_n218), .C2(inst3_n2792), .A(inst3_n2304),
        .B(inst3_n2303), .ZN(inst3_stateArray_S03reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst3_U501 ( .A1(inst3_n2610), .A2(ciphertext3[95]), .B1(
        inst3_n2392), .B2(inst3_n2302), .ZN(inst3_n2303) );
  XNOR2_X1 inst3_U500 ( .A(inst3_n2301), .B(inst3_n2300), .ZN(inst3_n2302) );
  AOI22_X1 inst3_U499 ( .A1(inst3_n216), .A2(ciphertext3[94]), .B1(inst3_n206),
        .B2(ciphertext3[126]), .ZN(inst3_n2300) );
  AOI22_X1 inst3_U498 ( .A1(inst3_n220), .A2(inst3_n2789), .B1(inst3_n2788),
        .B2(ciphertext3[95]), .ZN(inst3_n2301) );
  AOI22_X1 inst3_U497 ( .A1(inst3_n2474), .A2(ciphertext3[103]), .B1(
        plaintext3[103]), .B2(inst3_n2655), .ZN(inst3_n2304) );
  INV_X1 inst3_U496 ( .A(inst3_n2799), .ZN(inst3_n2474) );
  OAI211_X1 inst3_U495 ( .C1(inst3_n1207), .C2(inst3_n2775), .A(inst3_n2299),
        .B(inst3_n2298), .ZN(inst3_stateArray_S31reg_gff_1_SFF_2_n6) );
  NAND2_X1 inst3_U494 ( .A1(plaintext3[18]), .A2(inst3_n2727), .ZN(inst3_n2298) );
  AOI22_X1 inst3_U493 ( .A1(inst3_n2756), .A2(ciphertext3[18]), .B1(
        inst3_n2794), .B2(ciphertext3[26]), .ZN(inst3_n2299) );
  OAI211_X1 inst3_U492 ( .C1(inst3_n1205), .C2(inst3_n2775), .A(inst3_n2297),
        .B(inst3_n2296), .ZN(inst3_stateArray_S31reg_gff_1_SFF_4_n6) );
  NAND2_X1 inst3_U491 ( .A1(plaintext3[20]), .A2(inst3_n2727), .ZN(inst3_n2296) );
  AOI22_X1 inst3_U490 ( .A1(inst3_n2750), .A2(ciphertext3[20]), .B1(
        inst3_n2794), .B2(ciphertext3[28]), .ZN(inst3_n2297) );
  OAI211_X1 inst3_U489 ( .C1(inst3_n2797), .C2(inst3_n2295), .A(inst3_n2294),
        .B(inst3_n2293), .ZN(inst3_stateArray_S13reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst3_U488 ( .A1(inst3_n2555), .A2(ciphertext3[56]), .B1(
        ciphertext3[88]), .B2(inst3_n2292), .ZN(inst3_n2293) );
  AOI22_X1 inst3_U487 ( .A1(done3), .A2(ciphertext3[64]), .B1(plaintext3[64]),
        .B2(inst3_n2727), .ZN(inst3_n2294) );
  XNOR2_X1 inst3_U486 ( .A(inst3_n2786), .B(inst3_n2291), .ZN(inst3_n2295) );
  AOI22_X1 inst3_U485 ( .A1(inst3_n210), .A2(inst3_n2290), .B1(inst3_n2289),
        .B2(ciphertext3[120]), .ZN(inst3_n2291) );
  AOI22_X1 inst3_U484 ( .A1(inst3_n199), .A2(ciphertext3[56]), .B1(inst3_n2810), .B2(ciphertext3[24]), .ZN(inst3_n2786) );
  OAI211_X1 inst3_U483 ( .C1(inst3_n2288), .C2(inst3_n2784), .A(inst3_n2287),
        .B(inst3_n2286), .ZN(inst3_stateArray_S13reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U482 ( .A1(inst3_n2555), .A2(ciphertext3[57]), .B1(
        ciphertext3[89]), .B2(inst3_n2292), .ZN(inst3_n2286) );
  AOI22_X1 inst3_U481 ( .A1(inst3_n2750), .A2(ciphertext3[65]), .B1(
        plaintext3[65]), .B2(inst3_n2710), .ZN(inst3_n2287) );
  XNOR2_X1 inst3_U480 ( .A(inst3_n2285), .B(inst3_n2284), .ZN(inst3_n2288) );
  AOI22_X1 inst3_U479 ( .A1(inst3_n209), .A2(inst3_n2290), .B1(inst3_n2289),
        .B2(ciphertext3[88]), .ZN(inst3_n2284) );
  XNOR2_X1 inst3_U478 ( .A(inst3_n2776), .B(inst3_n2283), .ZN(inst3_n2285) );
  AOI22_X1 inst3_U477 ( .A1(inst3_n198), .A2(ciphertext3[56]), .B1(inst3_n2810), .B2(ciphertext3[121]), .ZN(inst3_n2283) );
  AOI22_X1 inst3_U476 ( .A1(inst3_n191), .A2(ciphertext3[57]), .B1(inst3_n2811), .B2(ciphertext3[25]), .ZN(inst3_n2776) );
  OAI211_X1 inst3_U475 ( .C1(inst3_n2282), .C2(inst3_n2784), .A(inst3_n2281),
        .B(inst3_n2280), .ZN(inst3_stateArray_S13reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U474 ( .A1(inst3_n2555), .A2(ciphertext3[58]), .B1(
        ciphertext3[90]), .B2(inst3_n2292), .ZN(inst3_n2280) );
  AOI22_X1 inst3_U473 ( .A1(inst3_n2750), .A2(ciphertext3[66]), .B1(
        plaintext3[66]), .B2(inst3_n2774), .ZN(inst3_n2281) );
  XNOR2_X1 inst3_U472 ( .A(inst3_n2279), .B(inst3_n2278), .ZN(inst3_n2282) );
  AOI22_X1 inst3_U471 ( .A1(inst3_n197), .A2(ciphertext3[57]), .B1(inst3_n2811), .B2(ciphertext3[89]), .ZN(inst3_n2278) );
  XNOR2_X1 inst3_U470 ( .A(inst3_n2277), .B(inst3_n193), .ZN(inst3_n2279) );
  OAI211_X1 inst3_U469 ( .C1(inst3_n2797), .C2(inst3_n2276), .A(inst3_n2275),
        .B(inst3_n2274), .ZN(inst3_stateArray_S13reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U468 ( .A1(inst3_n2555), .A2(ciphertext3[59]), .B1(
        ciphertext3[91]), .B2(inst3_n2292), .ZN(inst3_n2274) );
  AOI22_X1 inst3_U467 ( .A1(inst3_n2756), .A2(ciphertext3[67]), .B1(
        plaintext3[67]), .B2(inst3_n2713), .ZN(inst3_n2275) );
  XNOR2_X1 inst3_U466 ( .A(inst3_n2273), .B(inst3_n2272), .ZN(inst3_n2276) );
  AOI22_X1 inst3_U465 ( .A1(inst3_n202), .A2(inst3_n2289), .B1(inst3_n2290),
        .B2(ciphertext3[123]), .ZN(inst3_n2272) );
  INV_X1 inst3_U464 ( .A(inst3_n2290), .ZN(inst3_n2289) );
  XNOR2_X1 inst3_U463 ( .A(inst3_n2765), .B(inst3_n2327), .ZN(inst3_n2273) );
  AOI22_X1 inst3_U462 ( .A1(inst3_n194), .A2(inst3_n193), .B1(ciphertext3[58]),
        .B2(ciphertext3[90]), .ZN(inst3_n2327) );
  AOI22_X1 inst3_U461 ( .A1(ciphertext3[27]), .A2(inst3_n196), .B1(
        ciphertext3[59]), .B2(inst3_n2821), .ZN(inst3_n2765) );
  OAI211_X1 inst3_U460 ( .C1(inst3_n2271), .C2(inst3_n2797), .A(inst3_n2270),
        .B(inst3_n2269), .ZN(inst3_stateArray_S13reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U459 ( .A1(inst3_n2555), .A2(ciphertext3[60]), .B1(
        ciphertext3[92]), .B2(inst3_n2292), .ZN(inst3_n2269) );
  AOI22_X1 inst3_U458 ( .A1(inst3_n2750), .A2(ciphertext3[68]), .B1(
        plaintext3[68]), .B2(inst3_n2527), .ZN(inst3_n2270) );
  XNOR2_X1 inst3_U457 ( .A(inst3_n2268), .B(inst3_n2267), .ZN(inst3_n2271) );
  AOI22_X1 inst3_U456 ( .A1(inst3_n201), .A2(inst3_n2767), .B1(inst3_n2766),
        .B2(ciphertext3[91]), .ZN(inst3_n2267) );
  INV_X1 inst3_U455 ( .A(inst3_n2767), .ZN(inst3_n2766) );
  XNOR2_X1 inst3_U454 ( .A(inst3_n2290), .B(inst3_n2266), .ZN(inst3_n2268) );
  AOI22_X1 inst3_U453 ( .A1(ciphertext3[60]), .A2(inst3_n196), .B1(
        ciphertext3[59]), .B2(inst3_n2822), .ZN(inst3_n2266) );
  AOI22_X1 inst3_U452 ( .A1(inst3_n219), .A2(inst3_n220), .B1(ciphertext3[95]),
        .B2(ciphertext3[63]), .ZN(inst3_n2290) );
  OAI211_X1 inst3_U451 ( .C1(inst3_n2797), .C2(inst3_n2265), .A(inst3_n2264),
        .B(inst3_n2263), .ZN(inst3_stateArray_S13reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst3_U450 ( .A1(inst3_n2555), .A2(ciphertext3[61]), .B1(
        ciphertext3[93]), .B2(inst3_n2292), .ZN(inst3_n2263) );
  AOI22_X1 inst3_U449 ( .A1(inst3_n2750), .A2(ciphertext3[69]), .B1(
        plaintext3[69]), .B2(inst3_n2713), .ZN(inst3_n2264) );
  XNOR2_X1 inst3_U448 ( .A(inst3_n2311), .B(inst3_n2262), .ZN(inst3_n2265) );
  AOI22_X1 inst3_U447 ( .A1(inst3_n2261), .A2(ciphertext3[61]), .B1(
        inst3_n2823), .B2(inst3_n2260), .ZN(inst3_n2262) );
  OAI211_X1 inst3_U446 ( .C1(inst3_n2259), .C2(inst3_n2797), .A(inst3_n2258),
        .B(inst3_n2257), .ZN(inst3_stateArray_S13reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst3_U445 ( .A1(inst3_n2555), .A2(ciphertext3[62]), .B1(
        ciphertext3[94]), .B2(inst3_n2292), .ZN(inst3_n2257) );
  AOI22_X1 inst3_U444 ( .A1(inst3_n2750), .A2(ciphertext3[70]), .B1(
        plaintext3[70]), .B2(inst3_n2527), .ZN(inst3_n2258) );
  XNOR2_X1 inst3_U443 ( .A(inst3_n2319), .B(inst3_n2256), .ZN(inst3_n2259) );
  AOI22_X1 inst3_U442 ( .A1(ciphertext3[62]), .A2(inst3_n2255), .B1(
        inst3_n2254), .B2(inst3_n2809), .ZN(inst3_n2256) );
  OAI211_X1 inst3_U441 ( .C1(inst3_n2253), .C2(inst3_n2797), .A(inst3_n2252),
        .B(inst3_n2251), .ZN(inst3_stateArray_S13reg_gff_1_SFF_7_n5) );
  AOI22_X1 inst3_U440 ( .A1(inst3_n2555), .A2(ciphertext3[63]), .B1(
        ciphertext3[95]), .B2(inst3_n2292), .ZN(inst3_n2251) );
  NAND2_X1 inst3_U439 ( .A1(inst3_n2792), .A2(inst3_n2763), .ZN(inst3_n2292)
         );
  AOI22_X1 inst3_U438 ( .A1(inst3_n2750), .A2(ciphertext3[71]), .B1(
        plaintext3[71]), .B2(inst3_n2506), .ZN(inst3_n2252) );
  XNOR2_X1 inst3_U437 ( .A(inst3_n2332), .B(inst3_n2250), .ZN(inst3_n2253) );
  AOI22_X1 inst3_U436 ( .A1(inst3_n218), .A2(inst3_n2788), .B1(inst3_n2789),
        .B2(ciphertext3[127]), .ZN(inst3_n2250) );
  OAI211_X1 inst3_U435 ( .C1(inst3_n2794), .C2(inst3_n444), .A(inst3_n6), .B(
        inst3_n2249), .ZN(inst3_calcRCon_n51) );
  NAND2_X1 inst3_U434 ( .A1(inst3_n2794), .A2(inst3_n2803), .ZN(inst3_n2249)
         );
  OAI221_X1 inst3_U433 ( .B1(inst3_n2794), .B2(inst3_n581), .C1(inst3_n2763),
        .C2(inst3_n499), .A(inst3_n6), .ZN(inst3_calcRCon_n49) );
  OAI221_X1 inst3_U432 ( .B1(inst3_n2794), .B2(inst3_n1071), .C1(inst3_n2760),
        .C2(inst3_n718), .A(inst3_n6), .ZN(inst3_calcRCon_n44) );
  OAI21_X1 inst3_U431 ( .B1(inst3_n210), .B2(inst3_n2799), .A(inst3_n2248),
        .ZN(inst3_stateArray_S00reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst3_U430 ( .A1(ciphertext3[112]), .A2(inst3_n2753), .B1(
        plaintext3[120]), .B2(inst3_n2593), .ZN(inst3_n2248) );
  OAI21_X1 inst3_U429 ( .B1(inst3_n198), .B2(inst3_n2799), .A(inst3_n2247),
        .ZN(inst3_stateArray_S00reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U428 ( .A1(ciphertext3[113]), .A2(inst3_n2753), .B1(
        plaintext3[121]), .B2(inst3_n2710), .ZN(inst3_n2247) );
  OAI21_X1 inst3_U427 ( .B1(inst3_n2799), .B2(inst3_n2805), .A(inst3_n2246),
        .ZN(inst3_stateArray_S00reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U426 ( .A1(ciphertext3[114]), .A2(inst3_n1919), .B1(
        plaintext3[122]), .B2(inst3_n2713), .ZN(inst3_n2246) );
  OAI21_X1 inst3_U425 ( .B1(inst3_n202), .B2(inst3_n2799), .A(inst3_n2245),
        .ZN(inst3_stateArray_S00reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U424 ( .A1(ciphertext3[115]), .A2(inst3_n2753), .B1(
        plaintext3[123]), .B2(inst3_n2506), .ZN(inst3_n2245) );
  OAI21_X1 inst3_U423 ( .B1(inst3_n2799), .B2(inst3_n2802), .A(inst3_n2244),
        .ZN(inst3_stateArray_S00reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U422 ( .A1(ciphertext3[116]), .A2(inst3_n2753), .B1(
        plaintext3[124]), .B2(inst3_n2713), .ZN(inst3_n2244) );
  OAI21_X1 inst3_U421 ( .B1(inst3_n214), .B2(inst3_n2799), .A(inst3_n2243),
        .ZN(inst3_stateArray_S00reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst3_U420 ( .A1(ciphertext3[117]), .A2(inst3_n2753), .B1(
        plaintext3[125]), .B2(inst3_n2710), .ZN(inst3_n2243) );
  OAI21_X1 inst3_U419 ( .B1(inst3_n216), .B2(inst3_n2799), .A(inst3_n2242),
        .ZN(inst3_stateArray_S00reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst3_U418 ( .A1(ciphertext3[118]), .A2(inst3_n2753), .B1(
        plaintext3[126]), .B2(inst3_n2655), .ZN(inst3_n2242) );
  OAI21_X1 inst3_U417 ( .B1(inst3_n218), .B2(inst3_n2799), .A(inst3_n2241),
        .ZN(inst3_stateArray_S00reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst3_U416 ( .A1(ciphertext3[119]), .A2(inst3_n2753), .B1(
        plaintext3[127]), .B2(inst3_n2774), .ZN(inst3_n2241) );
  OAI21_X1 inst3_U415 ( .B1(inst3_n2799), .B2(inst3_n2849), .A(inst3_n2240),
        .ZN(inst3_stateArray_S01reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst3_U414 ( .A1(ciphertext3[104]), .A2(inst3_n2753), .B1(
        plaintext3[112]), .B2(inst3_n2774), .ZN(inst3_n2240) );
  OAI21_X1 inst3_U413 ( .B1(inst3_n2799), .B2(inst3_n2848), .A(inst3_n2239),
        .ZN(inst3_stateArray_S01reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U412 ( .A1(ciphertext3[105]), .A2(inst3_n2753), .B1(
        plaintext3[113]), .B2(inst3_n2655), .ZN(inst3_n2239) );
  OAI21_X1 inst3_U411 ( .B1(inst3_n2799), .B2(inst3_n2847), .A(inst3_n2238),
        .ZN(inst3_stateArray_S01reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U410 ( .A1(ciphertext3[106]), .A2(inst3_n2753), .B1(
        plaintext3[114]), .B2(inst3_n2713), .ZN(inst3_n2238) );
  OAI21_X1 inst3_U409 ( .B1(inst3_n2799), .B2(inst3_n2846), .A(inst3_n2237),
        .ZN(inst3_stateArray_S01reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U408 ( .A1(ciphertext3[107]), .A2(inst3_n2753), .B1(
        plaintext3[115]), .B2(inst3_n2727), .ZN(inst3_n2237) );
  OAI21_X1 inst3_U407 ( .B1(inst3_n2799), .B2(inst3_n2845), .A(inst3_n2236),
        .ZN(inst3_stateArray_S01reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U406 ( .A1(ciphertext3[108]), .A2(inst3_n2753), .B1(
        plaintext3[116]), .B2(inst3_n2713), .ZN(inst3_n2236) );
  OAI21_X1 inst3_U405 ( .B1(inst3_n2799), .B2(inst3_n2844), .A(inst3_n2235),
        .ZN(inst3_stateArray_S01reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst3_U404 ( .A1(ciphertext3[109]), .A2(inst3_n2753), .B1(
        plaintext3[117]), .B2(inst3_n2527), .ZN(inst3_n2235) );
  OAI21_X1 inst3_U403 ( .B1(inst3_n2799), .B2(inst3_n2843), .A(inst3_n2234),
        .ZN(inst3_stateArray_S01reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst3_U402 ( .A1(ciphertext3[110]), .A2(inst3_n2753), .B1(
        plaintext3[118]), .B2(inst3_n2774), .ZN(inst3_n2234) );
  OAI21_X1 inst3_U401 ( .B1(inst3_n2799), .B2(inst3_n2842), .A(inst3_n2233),
        .ZN(inst3_stateArray_S01reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst3_U400 ( .A1(ciphertext3[111]), .A2(inst3_n2753), .B1(
        plaintext3[119]), .B2(inst3_n2774), .ZN(inst3_n2233) );
  OAI21_X1 inst3_U399 ( .B1(inst3_n1273), .B2(inst3_n2775), .A(inst3_n2232),
        .ZN(inst3_stateArray_S02reg_gff_1_SFF_0_n6) );
  AOI22_X1 inst3_U398 ( .A1(ciphertext3[104]), .A2(inst3_n2543), .B1(
        plaintext3[104]), .B2(inst3_n2774), .ZN(inst3_n2232) );
  OAI21_X1 inst3_U397 ( .B1(inst3_n1272), .B2(inst3_n2775), .A(inst3_n2231),
        .ZN(inst3_stateArray_S02reg_gff_1_SFF_1_n6) );
  AOI22_X1 inst3_U396 ( .A1(ciphertext3[105]), .A2(inst3_n2584), .B1(
        plaintext3[105]), .B2(inst3_n2774), .ZN(inst3_n2231) );
  OAI21_X1 inst3_U395 ( .B1(inst3_n1271), .B2(inst3_n2775), .A(inst3_n2230),
        .ZN(inst3_stateArray_S02reg_gff_1_SFF_2_n6) );
  AOI22_X1 inst3_U394 ( .A1(ciphertext3[106]), .A2(inst3_n2474), .B1(
        plaintext3[106]), .B2(inst3_n2774), .ZN(inst3_n2230) );
  OAI21_X1 inst3_U393 ( .B1(inst3_n1270), .B2(inst3_n2775), .A(inst3_n2229),
        .ZN(inst3_stateArray_S02reg_gff_1_SFF_3_n6) );
  AOI22_X1 inst3_U392 ( .A1(ciphertext3[107]), .A2(inst3_n2487), .B1(
        plaintext3[107]), .B2(inst3_n2774), .ZN(inst3_n2229) );
  OAI21_X1 inst3_U391 ( .B1(inst3_n1269), .B2(inst3_n2775), .A(inst3_n2228),
        .ZN(inst3_stateArray_S02reg_gff_1_SFF_4_n6) );
  AOI22_X1 inst3_U390 ( .A1(ciphertext3[108]), .A2(inst3_n2584), .B1(
        plaintext3[108]), .B2(inst3_n2774), .ZN(inst3_n2228) );
  OAI21_X1 inst3_U389 ( .B1(inst3_n1268), .B2(inst3_n2775), .A(inst3_n2227),
        .ZN(inst3_stateArray_S02reg_gff_1_SFF_5_n6) );
  AOI22_X1 inst3_U388 ( .A1(ciphertext3[109]), .A2(inst3_n2538), .B1(
        plaintext3[109]), .B2(inst3_n2774), .ZN(inst3_n2227) );
  OAI21_X1 inst3_U387 ( .B1(inst3_n1267), .B2(inst3_n2775), .A(inst3_n2226),
        .ZN(inst3_stateArray_S02reg_gff_1_SFF_6_n6) );
  AOI22_X1 inst3_U386 ( .A1(ciphertext3[110]), .A2(inst3_n2538), .B1(
        plaintext3[110]), .B2(inst3_n2774), .ZN(inst3_n2226) );
  OAI21_X1 inst3_U385 ( .B1(inst3_n1266), .B2(inst3_n2775), .A(inst3_n2225),
        .ZN(inst3_stateArray_S02reg_gff_1_SFF_7_n6) );
  AOI22_X1 inst3_U384 ( .A1(ciphertext3[111]), .A2(inst3_n2487), .B1(
        plaintext3[111]), .B2(inst3_n2713), .ZN(inst3_n2225) );
  OAI211_X1 inst3_U383 ( .C1(inst3_n2797), .C2(inst3_n2224), .A(inst3_n2223),
        .B(inst3_n2222), .ZN(inst3_stateArray_S23reg_gff_1_SFF_0_n6) );
  AOI21_X1 inst3_U382 ( .B1(inst3_n2794), .B2(ciphertext3[48]), .A(inst3_n2221), .ZN(inst3_n2222) );
  OAI22_X1 inst3_U381 ( .A1(inst3_n199), .A2(inst3_n2461), .B1(inst3_n2792),
        .B2(inst3_n2810), .ZN(inst3_n2221) );
  AOI22_X1 inst3_U380 ( .A1(inst3_n2750), .A2(ciphertext3[32]), .B1(
        plaintext3[32]), .B2(inst3_n2774), .ZN(inst3_n2223) );
  XNOR2_X1 inst3_U379 ( .A(inst3_n2345), .B(inst3_n2220), .ZN(inst3_n2224) );
  AOI22_X1 inst3_U378 ( .A1(inst3_n199), .A2(inst3_n2789), .B1(inst3_n2788),
        .B2(ciphertext3[24]), .ZN(inst3_n2220) );
  INV_X1 inst3_U377 ( .A(inst3_n2789), .ZN(inst3_n2788) );
  OAI211_X1 inst3_U376 ( .C1(inst3_n2219), .C2(inst3_n2797), .A(inst3_n2218),
        .B(inst3_n2217), .ZN(inst3_stateArray_S23reg_gff_1_SFF_5_n5) );
  AOI21_X1 inst3_U375 ( .B1(inst3_n2794), .B2(ciphertext3[53]), .A(inst3_n2216), .ZN(inst3_n2217) );
  OAI22_X1 inst3_U374 ( .A1(inst3_n2461), .A2(inst3_n2807), .B1(inst3_n2792),
        .B2(inst3_n2823), .ZN(inst3_n2216) );
  AOI22_X1 inst3_U373 ( .A1(inst3_n2750), .A2(ciphertext3[37]), .B1(
        plaintext3[37]), .B2(inst3_n2806), .ZN(inst3_n2218) );
  XNOR2_X1 inst3_U372 ( .A(inst3_n2215), .B(inst3_n2214), .ZN(inst3_n2219) );
  AOI22_X1 inst3_U371 ( .A1(inst3_n2261), .A2(ciphertext3[28]), .B1(inst3_n207), .B2(inst3_n2260), .ZN(inst3_n2214) );
  INV_X1 inst3_U370 ( .A(inst3_n2261), .ZN(inst3_n2260) );
  AOI22_X1 inst3_U369 ( .A1(ciphertext3[60]), .A2(inst3_n190), .B1(
        ciphertext3[93]), .B2(inst3_n2822), .ZN(inst3_n2215) );
  OAI211_X1 inst3_U368 ( .C1(inst3_n2213), .C2(inst3_n2784), .A(inst3_n2212),
        .B(inst3_n2211), .ZN(inst3_stateArray_S23reg_gff_1_SFF_6_n5) );
  AOI21_X1 inst3_U367 ( .B1(inst3_n2794), .B2(ciphertext3[54]), .A(inst3_n2210), .ZN(inst3_n2211) );
  OAI22_X1 inst3_U366 ( .A1(inst3_n215), .A2(inst3_n2461), .B1(inst3_n2792),
        .B2(inst3_n2809), .ZN(inst3_n2210) );
  AOI22_X1 inst3_U365 ( .A1(inst3_n2750), .A2(ciphertext3[38]), .B1(
        plaintext3[38]), .B2(inst3_n2806), .ZN(inst3_n2212) );
  XNOR2_X1 inst3_U364 ( .A(inst3_n2209), .B(inst3_n2208), .ZN(inst3_n2213) );
  AOI22_X1 inst3_U363 ( .A1(inst3_n206), .A2(inst3_n2807), .B1(ciphertext3[29]), .B2(ciphertext3[94]), .ZN(inst3_n2208) );
  AOI22_X1 inst3_U362 ( .A1(inst3_n2254), .A2(ciphertext3[61]), .B1(
        inst3_n2823), .B2(inst3_n2255), .ZN(inst3_n2209) );
  INV_X1 inst3_U361 ( .A(inst3_n2254), .ZN(inst3_n2255) );
  OAI211_X1 inst3_U360 ( .C1(inst3_n2207), .C2(inst3_n2797), .A(inst3_n2206),
        .B(inst3_n2205), .ZN(inst3_stateArray_S23reg_gff_1_SFF_7_n5) );
  AOI21_X1 inst3_U359 ( .B1(inst3_n2794), .B2(ciphertext3[55]), .A(inst3_n2204), .ZN(inst3_n2205) );
  OAI22_X1 inst3_U358 ( .A1(inst3_n219), .A2(inst3_n2792), .B1(inst3_n2461),
        .B2(inst3_n2808), .ZN(inst3_n2204) );
  AOI22_X1 inst3_U357 ( .A1(inst3_n2750), .A2(ciphertext3[39]), .B1(
        plaintext3[39]), .B2(inst3_n2806), .ZN(inst3_n2206) );
  XNOR2_X1 inst3_U356 ( .A(inst3_n2203), .B(inst3_n2202), .ZN(inst3_n2207) );
  AOI22_X1 inst3_U355 ( .A1(inst3_n215), .A2(inst3_n2809), .B1(ciphertext3[62]), .B2(ciphertext3[30]), .ZN(inst3_n2202) );
  AOI22_X1 inst3_U354 ( .A1(ciphertext3[31]), .A2(inst3_n2389), .B1(
        inst3_n2388), .B2(inst3_n2808), .ZN(inst3_n2203) );
  INV_X1 inst3_U353 ( .A(inst3_n2389), .ZN(inst3_n2388) );
  OAI211_X1 inst3_U352 ( .C1(inst3_n2201), .C2(inst3_n2784), .A(inst3_n2200),
        .B(inst3_n2199), .ZN(inst3_stateArray_S23reg_gff_1_SFF_3_n6) );
  AOI21_X1 inst3_U351 ( .B1(inst3_n2794), .B2(ciphertext3[51]), .A(inst3_n2198), .ZN(inst3_n2199) );
  OAI22_X1 inst3_U350 ( .A1(inst3_n196), .A2(inst3_n2792), .B1(inst3_n2461),
        .B2(inst3_n2821), .ZN(inst3_n2198) );
  AOI22_X1 inst3_U349 ( .A1(inst3_n2750), .A2(ciphertext3[35]), .B1(
        plaintext3[35]), .B2(inst3_n2806), .ZN(inst3_n2200) );
  INV_X1 inst3_U348 ( .A(inst3_n2720), .ZN(inst3_n2750) );
  XNOR2_X1 inst3_U347 ( .A(inst3_n2197), .B(inst3_n2196), .ZN(inst3_n2201) );
  AOI22_X1 inst3_U346 ( .A1(ciphertext3[27]), .A2(inst3_n2310), .B1(
        inst3_n2309), .B2(inst3_n2821), .ZN(inst3_n2196) );
  INV_X1 inst3_U345 ( .A(inst3_n2310), .ZN(inst3_n2309) );
  XNOR2_X1 inst3_U344 ( .A(inst3_n2789), .B(inst3_n2195), .ZN(inst3_n2197) );
  AOI22_X1 inst3_U343 ( .A1(inst3_n203), .A2(inst3_n193), .B1(ciphertext3[58]),
        .B2(ciphertext3[26]), .ZN(inst3_n2195) );
  AOI22_X1 inst3_U342 ( .A1(ciphertext3[31]), .A2(inst3_n219), .B1(
        ciphertext3[63]), .B2(inst3_n2808), .ZN(inst3_n2789) );
  NAND2_X1 inst3_U341 ( .A1(inst3_n2194), .A2(inst3_n2193), .ZN(
        inst3_stateArray_S33reg_gff_1_SFF_0_n5) );
  AOI22_X1 inst3_U340 ( .A1(inst3_n2192), .A2(inst3_n2191), .B1(inst3_n2190),
        .B2(inst3_n2189), .ZN(inst3_n2193) );
  AOI211_X1 inst3_U339 ( .C1(plaintext3[0]), .C2(inst3_n2806), .A(inst3_n2188),
        .B(inst3_n2187), .ZN(inst3_n2194) );
  OAI22_X1 inst3_U338 ( .A1(inst3_n2186), .A2(inst3_n2784), .B1(inst3_n1201),
        .B2(inst3_n2720), .ZN(inst3_n2187) );
  XNOR2_X1 inst3_U337 ( .A(inst3_n2345), .B(inst3_n2185), .ZN(inst3_n2186) );
  AOI22_X1 inst3_U336 ( .A1(inst3_n2184), .A2(inst3_n2810), .B1(
        ciphertext3[56]), .B2(inst3_n2183), .ZN(inst3_n2185) );
  AOI22_X1 inst3_U335 ( .A1(inst3_n210), .A2(inst3_n209), .B1(ciphertext3[88]),
        .B2(ciphertext3[120]), .ZN(inst3_n2345) );
  OAI22_X1 inst3_U334 ( .A1(inst3_n199), .A2(inst3_n2792), .B1(inst3_n1209),
        .B2(inst3_n2760), .ZN(inst3_n2188) );
  NAND2_X1 inst3_U333 ( .A1(inst3_n2182), .A2(inst3_n2181), .ZN(
        inst3_stateArray_S33reg_gff_1_SFF_1_n5) );
  AOI22_X1 inst3_U332 ( .A1(inst3_n2180), .A2(inst3_n2191), .B1(inst3_n2190),
        .B2(inst3_n2179), .ZN(inst3_n2181) );
  AOI211_X1 inst3_U331 ( .C1(plaintext3[1]), .C2(inst3_n2806), .A(inst3_n2178),
        .B(inst3_n2177), .ZN(inst3_n2182) );
  OAI22_X1 inst3_U330 ( .A1(inst3_n2176), .A2(inst3_n2784), .B1(inst3_n1200),
        .B2(inst3_n2720), .ZN(inst3_n2177) );
  XNOR2_X1 inst3_U329 ( .A(inst3_n2175), .B(inst3_n2174), .ZN(inst3_n2176) );
  AOI22_X1 inst3_U328 ( .A1(inst3_n210), .A2(inst3_n2184), .B1(inst3_n2183),
        .B2(ciphertext3[120]), .ZN(inst3_n2174) );
  XNOR2_X1 inst3_U327 ( .A(inst3_n2787), .B(inst3_n2173), .ZN(inst3_n2175) );
  AOI22_X1 inst3_U326 ( .A1(inst3_n199), .A2(ciphertext3[57]), .B1(inst3_n2811), .B2(ciphertext3[24]), .ZN(inst3_n2173) );
  AOI22_X1 inst3_U325 ( .A1(inst3_n198), .A2(inst3_n197), .B1(ciphertext3[89]),
        .B2(ciphertext3[121]), .ZN(inst3_n2787) );
  OAI22_X1 inst3_U324 ( .A1(inst3_n191), .A2(inst3_n2792), .B1(inst3_n1208),
        .B2(inst3_n2760), .ZN(inst3_n2178) );
  NAND2_X1 inst3_U323 ( .A1(inst3_n2172), .A2(inst3_n2171), .ZN(
        inst3_stateArray_S33reg_gff_1_SFF_2_n5) );
  AOI22_X1 inst3_U322 ( .A1(inst3_n2170), .A2(inst3_n2190), .B1(inst3_n2191),
        .B2(inst3_n2169), .ZN(inst3_n2171) );
  AOI211_X1 inst3_U321 ( .C1(plaintext3[2]), .C2(inst3_n2806), .A(inst3_n2168),
        .B(inst3_n2167), .ZN(inst3_n2172) );
  OAI22_X1 inst3_U320 ( .A1(inst3_n1199), .A2(inst3_n2720), .B1(inst3_n2784),
        .B2(inst3_n2166), .ZN(inst3_n2167) );
  XNOR2_X1 inst3_U319 ( .A(inst3_n2165), .B(inst3_n2164), .ZN(inst3_n2166) );
  AOI22_X1 inst3_U318 ( .A1(inst3_n198), .A2(ciphertext3[58]), .B1(inst3_n193),
        .B2(ciphertext3[121]), .ZN(inst3_n2164) );
  XNOR2_X1 inst3_U317 ( .A(inst3_n191), .B(inst3_n2779), .ZN(inst3_n2165) );
  AOI22_X1 inst3_U316 ( .A1(ciphertext3[122]), .A2(inst3_n194), .B1(
        ciphertext3[90]), .B2(inst3_n2805), .ZN(inst3_n2779) );
  OAI22_X1 inst3_U315 ( .A1(inst3_n203), .A2(inst3_n2792), .B1(inst3_n1207),
        .B2(inst3_n2760), .ZN(inst3_n2168) );
  NAND2_X1 inst3_U314 ( .A1(inst3_n2163), .A2(inst3_n2162), .ZN(
        inst3_stateArray_S33reg_gff_1_SFF_3_n5) );
  AOI22_X1 inst3_U313 ( .A1(inst3_n2161), .A2(inst3_n2191), .B1(inst3_n2160),
        .B2(inst3_n2190), .ZN(inst3_n2162) );
  AOI211_X1 inst3_U312 ( .C1(plaintext3[3]), .C2(inst3_n2806), .A(inst3_n2159),
        .B(inst3_n2158), .ZN(inst3_n2163) );
  OAI22_X1 inst3_U311 ( .A1(inst3_n2157), .A2(inst3_n2784), .B1(inst3_n1198),
        .B2(inst3_n2720), .ZN(inst3_n2158) );
  XNOR2_X1 inst3_U310 ( .A(inst3_n2156), .B(inst3_n2155), .ZN(inst3_n2157) );
  AOI22_X1 inst3_U309 ( .A1(inst3_n2184), .A2(inst3_n196), .B1(ciphertext3[59]), .B2(inst3_n2183), .ZN(inst3_n2155) );
  INV_X1 inst3_U308 ( .A(inst3_n2184), .ZN(inst3_n2183) );
  XNOR2_X1 inst3_U307 ( .A(inst3_n2310), .B(inst3_n2277), .ZN(inst3_n2156) );
  AOI22_X1 inst3_U306 ( .A1(ciphertext3[122]), .A2(inst3_n203), .B1(
        ciphertext3[26]), .B2(inst3_n2805), .ZN(inst3_n2277) );
  AOI22_X1 inst3_U305 ( .A1(inst3_n202), .A2(inst3_n201), .B1(ciphertext3[91]),
        .B2(ciphertext3[123]), .ZN(inst3_n2310) );
  OAI22_X1 inst3_U304 ( .A1(inst3_n1206), .A2(inst3_n2763), .B1(inst3_n2792),
        .B2(inst3_n2821), .ZN(inst3_n2159) );
  NAND2_X1 inst3_U303 ( .A1(inst3_n2154), .A2(inst3_n2153), .ZN(
        inst3_stateArray_S33reg_gff_1_SFF_4_n5) );
  AOI22_X1 inst3_U302 ( .A1(inst3_n2190), .A2(inst3_n2152), .B1(inst3_n2191),
        .B2(inst3_n2151), .ZN(inst3_n2153) );
  AOI211_X1 inst3_U301 ( .C1(plaintext3[4]), .C2(inst3_n2806), .A(inst3_n2150),
        .B(inst3_n2149), .ZN(inst3_n2154) );
  OAI22_X1 inst3_U300 ( .A1(inst3_n2148), .A2(inst3_n2784), .B1(inst3_n1197),
        .B2(inst3_n2720), .ZN(inst3_n2149) );
  XNOR2_X1 inst3_U299 ( .A(inst3_n2147), .B(inst3_n2146), .ZN(inst3_n2148) );
  XNOR2_X1 inst3_U298 ( .A(inst3_n202), .B(inst3_n2311), .ZN(inst3_n2146) );
  AOI22_X1 inst3_U297 ( .A1(inst3_n212), .A2(ciphertext3[60]), .B1(inst3_n2822), .B2(ciphertext3[92]), .ZN(inst3_n2311) );
  XOR2_X1 inst3_U296 ( .A(inst3_n2145), .B(inst3_n2184), .Z(inst3_n2147) );
  AOI22_X1 inst3_U295 ( .A1(inst3_n218), .A2(ciphertext3[31]), .B1(inst3_n2808), .B2(ciphertext3[127]), .ZN(inst3_n2184) );
  AOI22_X1 inst3_U294 ( .A1(ciphertext3[124]), .A2(ciphertext3[27]), .B1(
        inst3_n2821), .B2(inst3_n2802), .ZN(inst3_n2145) );
  OAI22_X1 inst3_U293 ( .A1(inst3_n207), .A2(inst3_n2792), .B1(inst3_n1205),
        .B2(inst3_n2760), .ZN(inst3_n2150) );
  NAND2_X1 inst3_U292 ( .A1(inst3_n2144), .A2(inst3_n2143), .ZN(
        inst3_stateArray_S33reg_gff_1_SFF_5_n5) );
  AOI22_X1 inst3_U291 ( .A1(inst3_n2142), .A2(inst3_n2191), .B1(inst3_n2190),
        .B2(inst3_n2141), .ZN(inst3_n2143) );
  AOI211_X1 inst3_U290 ( .C1(plaintext3[5]), .C2(inst3_n2806), .A(inst3_n2140),
        .B(inst3_n2139), .ZN(inst3_n2144) );
  OAI22_X1 inst3_U289 ( .A1(inst3_n2138), .A2(inst3_n2784), .B1(inst3_n1196),
        .B2(inst3_n2720), .ZN(inst3_n2139) );
  XNOR2_X1 inst3_U288 ( .A(inst3_n2137), .B(inst3_n2319), .ZN(inst3_n2138) );
  AOI22_X1 inst3_U287 ( .A1(ciphertext3[61]), .A2(inst3_n190), .B1(
        ciphertext3[93]), .B2(inst3_n2823), .ZN(inst3_n2319) );
  XNOR2_X1 inst3_U286 ( .A(inst3_n214), .B(inst3_n2767), .ZN(inst3_n2137) );
  AOI22_X1 inst3_U285 ( .A1(ciphertext3[124]), .A2(inst3_n207), .B1(
        ciphertext3[28]), .B2(inst3_n2802), .ZN(inst3_n2767) );
  OAI22_X1 inst3_U284 ( .A1(inst3_n1204), .A2(inst3_n2763), .B1(inst3_n2792),
        .B2(inst3_n2807), .ZN(inst3_n2140) );
  NAND2_X1 inst3_U283 ( .A1(inst3_n2136), .A2(inst3_n2135), .ZN(
        inst3_stateArray_S33reg_gff_1_SFF_6_n5) );
  AOI22_X1 inst3_U282 ( .A1(inst3_n2134), .A2(inst3_n2191), .B1(inst3_n2190),
        .B2(inst3_n2133), .ZN(inst3_n2135) );
  AOI211_X1 inst3_U281 ( .C1(plaintext3[6]), .C2(inst3_n2806), .A(inst3_n2132),
        .B(inst3_n2131), .ZN(inst3_n2136) );
  OAI22_X1 inst3_U280 ( .A1(inst3_n2130), .A2(inst3_n2784), .B1(inst3_n1195),
        .B2(inst3_n2720), .ZN(inst3_n2131) );
  XNOR2_X1 inst3_U279 ( .A(inst3_n2129), .B(inst3_n2261), .ZN(inst3_n2130) );
  AOI22_X1 inst3_U278 ( .A1(inst3_n214), .A2(ciphertext3[29]), .B1(inst3_n2807), .B2(ciphertext3[125]), .ZN(inst3_n2261) );
  XNOR2_X1 inst3_U277 ( .A(inst3_n216), .B(inst3_n2332), .ZN(inst3_n2129) );
  AOI22_X1 inst3_U276 ( .A1(ciphertext3[62]), .A2(inst3_n206), .B1(
        ciphertext3[94]), .B2(inst3_n2809), .ZN(inst3_n2332) );
  OAI22_X1 inst3_U275 ( .A1(inst3_n215), .A2(inst3_n2792), .B1(inst3_n1203),
        .B2(inst3_n2760), .ZN(inst3_n2132) );
  INV_X1 inst3_U274 ( .A(inst3_n2794), .ZN(inst3_n2760) );
  OAI211_X1 inst3_U273 ( .C1(inst3_n2128), .C2(inst3_n2127), .A(inst3_n2126),
        .B(inst3_n2125), .ZN(inst3_stateArray_S33reg_gff_1_SFF_7_n5) );
  NAND2_X1 inst3_U272 ( .A1(inst3_n2124), .A2(inst3_n2191), .ZN(inst3_n2125)
         );
  NOR2_X1 inst3_U271 ( .A1(inst3_n2461), .A2(inst3_n2123), .ZN(inst3_n2191) );
  INV_X1 inst3_U270 ( .A(inst3_n2610), .ZN(inst3_n2461) );
  AOI211_X1 inst3_U269 ( .C1(plaintext3[7]), .C2(inst3_n2806), .A(inst3_n2122),
        .B(inst3_n2121), .ZN(inst3_n2126) );
  OAI22_X1 inst3_U268 ( .A1(inst3_n2120), .A2(inst3_n2784), .B1(inst3_n1194),
        .B2(inst3_n2720), .ZN(inst3_n2121) );
  INV_X1 inst3_U267 ( .A(inst3_n2392), .ZN(inst3_n2784) );
  INV_X1 inst3_U266 ( .A(inst3_n2797), .ZN(inst3_n2392) );
  NAND2_X1 inst3_U265 ( .A1(inst3_n2665), .A2(inst3_n2123), .ZN(inst3_n2797)
         );
  INV_X1 inst3_U264 ( .A(inst3_n2119), .ZN(inst3_n2665) );
  XNOR2_X1 inst3_U263 ( .A(inst3_n2118), .B(inst3_n2254), .ZN(inst3_n2120) );
  AOI22_X1 inst3_U262 ( .A1(inst3_n216), .A2(inst3_n215), .B1(ciphertext3[30]),
        .B2(ciphertext3[126]), .ZN(inst3_n2254) );
  XNOR2_X1 inst3_U261 ( .A(inst3_n219), .B(inst3_n2389), .ZN(inst3_n2118) );
  AOI22_X1 inst3_U260 ( .A1(inst3_n218), .A2(inst3_n220), .B1(ciphertext3[95]),
        .B2(ciphertext3[127]), .ZN(inst3_n2389) );
  OAI22_X1 inst3_U259 ( .A1(inst3_n1202), .A2(inst3_n2763), .B1(inst3_n2792),
        .B2(inst3_n2808), .ZN(inst3_n2122) );
  AND2_X1 inst3_U258 ( .A1(inst3_n2662), .A2(inst3_n2116), .ZN(inst3_n2117) );
  INV_X1 inst3_U257 ( .A(inst3_n2794), .ZN(inst3_n2763) );
  AND2_X2 inst3_U256 ( .A1(inst3_n2474), .A2(inst3_n2708), .ZN(inst3_n2794) );
  INV_X1 inst3_U255 ( .A(inst3_n2190), .ZN(inst3_n2127) );
  NOR2_X1 inst3_U254 ( .A1(inst3_n2116), .A2(inst3_n2668), .ZN(inst3_n2190) );
  OAI211_X1 inst3_U253 ( .C1(inst3_n2864), .C2(inst3_n2799), .A(inst3_n2115),
        .B(inst3_n2114), .ZN(inst3_KeyArray_S30reg_gff_1_SFF_3_n6) );
  OAI21_X1 inst3_U252 ( .B1(inst3_n224), .B2(inst3_n2113), .A(inst3_n2112),
        .ZN(inst3_n2114) );
  AOI21_X1 inst3_U251 ( .B1(inst3_n224), .B2(inst3_n2113), .A(inst3_n2648),
        .ZN(inst3_n2112) );
  XNOR2_X1 inst3_U250 ( .A(inst3_n2160), .B(inst3_n2111), .ZN(inst3_n2113) );
  NOR2_X1 inst3_U249 ( .A1(inst3_n321), .A2(inst3_n706), .ZN(inst3_n2111) );
  XNOR2_X1 inst3_U248 ( .A(inst3_n2110), .B(inst3_n2109), .ZN(inst3_n2160) );
  XNOR2_X1 inst3_U247 ( .A(inst3_n2108), .B(inst3_n2107), .ZN(inst3_n2110) );
  AOI22_X1 inst3_U246 ( .A1(inst3_n71), .A2(inst3_n2610), .B1(key3[27]), .B2(
        inst3_n2806), .ZN(inst3_n2115) );
  OAI211_X1 inst3_U245 ( .C1(inst3_n2863), .C2(inst3_n2799), .A(inst3_n2106),
        .B(inst3_n2105), .ZN(inst3_KeyArray_S30reg_gff_1_SFF_6_n6) );
  OAI21_X1 inst3_U244 ( .B1(inst3_n222), .B2(inst3_n2104), .A(inst3_n2103),
        .ZN(inst3_n2105) );
  AOI21_X1 inst3_U243 ( .B1(inst3_n222), .B2(inst3_n2104), .A(inst3_n2648),
        .ZN(inst3_n2103) );
  XNOR2_X1 inst3_U242 ( .A(inst3_n2102), .B(inst3_n2133), .ZN(inst3_n2104) );
  XNOR2_X1 inst3_U241 ( .A(inst3_n2101), .B(inst3_n2100), .ZN(inst3_n2133) );
  NOR2_X1 inst3_U240 ( .A1(inst3_n718), .A2(inst3_n321), .ZN(inst3_n2102) );
  AOI22_X1 inst3_U239 ( .A1(inst3_n68), .A2(inst3_n2610), .B1(key3[30]), .B2(
        inst3_n2806), .ZN(inst3_n2106) );
  OAI211_X1 inst3_U238 ( .C1(inst3_n2862), .C2(inst3_n2799), .A(inst3_n2099),
        .B(inst3_n2098), .ZN(inst3_KeyArray_S30reg_gff_1_SFF_1_n6) );
  OAI21_X1 inst3_U237 ( .B1(inst3_n226), .B2(inst3_n2097), .A(inst3_n2096),
        .ZN(inst3_n2098) );
  AOI21_X1 inst3_U236 ( .B1(inst3_n226), .B2(inst3_n2097), .A(inst3_n2648),
        .ZN(inst3_n2096) );
  XNOR2_X1 inst3_U235 ( .A(inst3_n2095), .B(inst3_n2179), .ZN(inst3_n2097) );
  XNOR2_X1 inst3_U234 ( .A(inst3_n2094), .B(inst3_n2093), .ZN(inst3_n2179) );
  XNOR2_X1 inst3_U233 ( .A(inst3_n2109), .B(inst3_n2092), .ZN(inst3_n2094) );
  XNOR2_X1 inst3_U232 ( .A(inst3_n2091), .B(inst3_n2090), .ZN(inst3_n2092) );
  XOR2_X1 inst3_U231 ( .A(inst3_n2089), .B(inst3_n2088), .Z(inst3_n2090) );
  XNOR2_X1 inst3_U230 ( .A(inst3_n2087), .B(inst3_n2086), .ZN(inst3_n2109) );
  NOR2_X1 inst3_U229 ( .A1(inst3_n499), .A2(inst3_n321), .ZN(inst3_n2095) );
  AOI22_X1 inst3_U228 ( .A1(inst3_n73), .A2(inst3_n2613), .B1(key3[25]), .B2(
        inst3_n2806), .ZN(inst3_n2099) );
  INV_X1 inst3_U227 ( .A(inst3_n2668), .ZN(inst3_n2613) );
  OAI211_X1 inst3_U226 ( .C1(inst3_n2861), .C2(inst3_n2799), .A(inst3_n2085),
        .B(inst3_n2084), .ZN(inst3_KeyArray_S30reg_gff_1_SFF_2_n6) );
  OAI21_X1 inst3_U225 ( .B1(inst3_n225), .B2(inst3_n2083), .A(inst3_n2082),
        .ZN(inst3_n2084) );
  AOI21_X1 inst3_U224 ( .B1(inst3_n225), .B2(inst3_n2083), .A(inst3_n2648),
        .ZN(inst3_n2082) );
  XNOR2_X1 inst3_U223 ( .A(inst3_n2081), .B(inst3_n2170), .ZN(inst3_n2083) );
  XNOR2_X1 inst3_U222 ( .A(inst3_n2080), .B(inst3_n2079), .ZN(inst3_n2170) );
  XNOR2_X1 inst3_U221 ( .A(inst3_n2093), .B(inst3_n2078), .ZN(inst3_n2079) );
  XNOR2_X1 inst3_U220 ( .A(inst3_n2077), .B(inst3_n2076), .ZN(inst3_n2080) );
  XOR2_X1 inst3_U219 ( .A(inst3_n2075), .B(inst3_n2074), .Z(inst3_n2076) );
  NOR2_X1 inst3_U218 ( .A1(inst3_n2073), .A2(inst3_n2072), .ZN(inst3_n2077) );
  AOI21_X1 inst3_U217 ( .B1(inst3_n2071), .B2(inst3_n2070), .A(inst3_n2069),
        .ZN(inst3_n2073) );
  NOR2_X1 inst3_U216 ( .A1(inst3_n581), .A2(inst3_n321), .ZN(inst3_n2081) );
  AOI22_X1 inst3_U215 ( .A1(inst3_n72), .A2(inst3_n2552), .B1(key3[26]), .B2(
        inst3_n2806), .ZN(inst3_n2085) );
  INV_X1 inst3_U214 ( .A(inst3_n2668), .ZN(inst3_n2552) );
  OAI211_X1 inst3_U213 ( .C1(inst3_n2837), .C2(inst3_n2668), .A(inst3_n2068),
        .B(inst3_n2067), .ZN(inst3_KeyArray_S30reg_gff_1_SFF_4_n6) );
  OAI21_X1 inst3_U212 ( .B1(inst3_n223), .B2(inst3_n2066), .A(inst3_n2065),
        .ZN(inst3_n2067) );
  AOI21_X1 inst3_U211 ( .B1(inst3_n223), .B2(inst3_n2066), .A(inst3_n2648),
        .ZN(inst3_n2065) );
  XNOR2_X1 inst3_U210 ( .A(inst3_n2064), .B(inst3_n2152), .ZN(inst3_n2066) );
  XNOR2_X1 inst3_U209 ( .A(inst3_n2075), .B(inst3_n2101), .ZN(inst3_n2152) );
  XNOR2_X1 inst3_U208 ( .A(inst3_n2063), .B(inst3_n2108), .ZN(inst3_n2101) );
  XNOR2_X1 inst3_U207 ( .A(inst3_n2062), .B(inst3_n2061), .ZN(inst3_n2108) );
  NAND2_X1 inst3_U206 ( .A1(inst3_n2060), .A2(inst3_n2059), .ZN(inst3_n2062)
         );
  NOR2_X1 inst3_U205 ( .A1(inst3_n321), .A2(inst3_n1081), .ZN(inst3_n2064) );
  AOI22_X1 inst3_U204 ( .A1(inst3_n78), .A2(inst3_n2474), .B1(key3[28]), .B2(
        inst3_n2806), .ZN(inst3_n2068) );
  OAI211_X1 inst3_U203 ( .C1(inst3_n2860), .C2(inst3_n2799), .A(inst3_n2058),
        .B(inst3_n2057), .ZN(inst3_KeyArray_S30reg_gff_1_SFF_7_n6) );
  OAI21_X1 inst3_U202 ( .B1(inst3_n2056), .B2(inst3_n2804), .A(inst3_n2055),
        .ZN(inst3_n2057) );
  AOI21_X1 inst3_U201 ( .B1(inst3_n2056), .B2(inst3_n2804), .A(inst3_n2648),
        .ZN(inst3_n2055) );
  XNOR2_X1 inst3_U200 ( .A(inst3_n2054), .B(inst3_n2128), .ZN(inst3_n2056) );
  XNOR2_X1 inst3_U199 ( .A(inst3_n2053), .B(inst3_n2100), .ZN(inst3_n2128) );
  XNOR2_X1 inst3_U198 ( .A(inst3_n2093), .B(inst3_n2052), .ZN(inst3_n2100) );
  OAI221_X1 inst3_U197 ( .B1(inst3_n2051), .B2(inst3_n2050), .C1(inst3_n2049),
        .C2(inst3_n2048), .A(inst3_n2047), .ZN(inst3_n2093) );
  INV_X1 inst3_U196 ( .A(inst3_n2048), .ZN(inst3_n2050) );
  XNOR2_X1 inst3_U195 ( .A(inst3_n2075), .B(inst3_n2061), .ZN(inst3_n2053) );
  XNOR2_X1 inst3_U194 ( .A(inst3_n2046), .B(inst3_n2074), .ZN(inst3_n2061) );
  XNOR2_X1 inst3_U193 ( .A(inst3_n2045), .B(inst3_n2044), .ZN(inst3_n2074) );
  NAND2_X1 inst3_U192 ( .A1(inst3_n2060), .A2(inst3_n2043), .ZN(inst3_n2045)
         );
  XNOR2_X1 inst3_U191 ( .A(inst3_n2042), .B(inst3_n2041), .ZN(inst3_n2060) );
  XNOR2_X1 inst3_U190 ( .A(inst3_n2040), .B(inst3_n2039), .ZN(inst3_n2042) );
  NAND2_X1 inst3_U189 ( .A1(inst3_n2038), .A2(inst3_n2037), .ZN(inst3_n2046)
         );
  XNOR2_X1 inst3_U188 ( .A(inst3_n2036), .B(inst3_n2086), .ZN(inst3_n2075) );
  NAND2_X1 inst3_U187 ( .A1(inst3_n2035), .A2(inst3_n2034), .ZN(inst3_n2086)
         );
  NOR2_X1 inst3_U186 ( .A1(inst3_n1071), .A2(inst3_n321), .ZN(inst3_n2054) );
  AOI22_X1 inst3_U185 ( .A1(inst3_n67), .A2(inst3_n2610), .B1(key3[31]), .B2(
        inst3_n2806), .ZN(inst3_n2058) );
  OAI211_X1 inst3_U184 ( .C1(inst3_n2859), .C2(inst3_n2799), .A(inst3_n2033),
        .B(inst3_n2032), .ZN(inst3_KeyArray_S30reg_gff_1_SFF_0_n6) );
  OAI21_X1 inst3_U183 ( .B1(inst3_n227), .B2(inst3_n2031), .A(inst3_n2030),
        .ZN(inst3_n2032) );
  AOI21_X1 inst3_U182 ( .B1(inst3_n227), .B2(inst3_n2031), .A(inst3_n2648),
        .ZN(inst3_n2030) );
  XNOR2_X1 inst3_U181 ( .A(inst3_n2029), .B(inst3_n2189), .ZN(inst3_n2031) );
  XNOR2_X1 inst3_U180 ( .A(inst3_n2036), .B(inst3_n2028), .ZN(inst3_n2189) );
  XNOR2_X1 inst3_U179 ( .A(inst3_n2027), .B(inst3_n2091), .ZN(inst3_n2028) );
  XOR2_X1 inst3_U178 ( .A(inst3_n2044), .B(inst3_n2026), .Z(inst3_n2091) );
  OAI211_X1 inst3_U177 ( .C1(inst3_n2025), .C2(inst3_n2024), .A(inst3_n2023),
        .B(inst3_n2034), .ZN(inst3_n2026) );
  MUX2_X1 inst3_U176 ( .A(inst3_n2022), .B(inst3_n2040), .S(inst3_n2021), .Z(
        inst3_n2034) );
  XOR2_X1 inst3_U175 ( .A(inst3_n2020), .B(inst3_n2019), .Z(inst3_n2044) );
  NAND2_X1 inst3_U174 ( .A1(inst3_n2047), .A2(inst3_n2018), .ZN(inst3_n2019)
         );
  XNOR2_X1 inst3_U173 ( .A(inst3_n2017), .B(inst3_n2016), .ZN(inst3_n2047) );
  XNOR2_X1 inst3_U172 ( .A(inst3_n2015), .B(inst3_n2014), .ZN(inst3_n2016) );
  XOR2_X1 inst3_U171 ( .A(inst3_n2013), .B(inst3_n2012), .Z(inst3_n2017) );
  XNOR2_X1 inst3_U170 ( .A(inst3_n2087), .B(inst3_n2011), .ZN(inst3_n2027) );
  NOR2_X1 inst3_U169 ( .A1(inst3_n2010), .A2(inst3_n2009), .ZN(inst3_n2087) );
  AND2_X1 inst3_U168 ( .A1(inst3_n2008), .A2(inst3_n2007), .ZN(inst3_n2036) );
  NOR2_X1 inst3_U167 ( .A1(inst3_n444), .A2(inst3_n321), .ZN(inst3_n2029) );
  AOI22_X1 inst3_U166 ( .A1(inst3_n74), .A2(inst3_n2555), .B1(key3[24]), .B2(
        inst3_n2713), .ZN(inst3_n2033) );
  INV_X1 inst3_U165 ( .A(inst3_n2668), .ZN(inst3_n2555) );
  OAI211_X1 inst3_U164 ( .C1(inst3_n2858), .C2(inst3_n2799), .A(inst3_n2006),
        .B(inst3_n2005), .ZN(inst3_KeyArray_S30reg_gff_1_SFF_5_n6) );
  OAI21_X1 inst3_U163 ( .B1(inst3_n228), .B2(inst3_n2004), .A(inst3_n2003),
        .ZN(inst3_n2005) );
  AOI21_X1 inst3_U162 ( .B1(inst3_n228), .B2(inst3_n2004), .A(inst3_n2648),
        .ZN(inst3_n2003) );
  INV_X2 inst3_U161 ( .A(inst3_n2119), .ZN(inst3_n2662) );
  XNOR2_X1 inst3_U160 ( .A(inst3_n2001), .B(inst3_n2141), .ZN(inst3_n2004) );
  XOR2_X1 inst3_U159 ( .A(inst3_n2000), .B(inst3_n2020), .Z(inst3_n2141) );
  NAND2_X1 inst3_U158 ( .A1(inst3_n1999), .A2(inst3_n1998), .ZN(inst3_n2020)
         );
  XNOR2_X1 inst3_U157 ( .A(inst3_n1997), .B(inst3_n1996), .ZN(inst3_n2000) );
  NAND2_X1 inst3_U156 ( .A1(inst3_n1995), .A2(inst3_n1994), .ZN(inst3_n1996)
         );
  XNOR2_X1 inst3_U155 ( .A(inst3_n2052), .B(inst3_n2078), .ZN(inst3_n1997) );
  XNOR2_X1 inst3_U154 ( .A(inst3_n1993), .B(inst3_n2011), .ZN(inst3_n2078) );
  XNOR2_X1 inst3_U153 ( .A(inst3_n1992), .B(inst3_n2089), .ZN(inst3_n2011) );
  NAND2_X1 inst3_U152 ( .A1(inst3_n1991), .A2(inst3_n2007), .ZN(inst3_n2089)
         );
  XOR2_X1 inst3_U151 ( .A(inst3_n1990), .B(inst3_n1989), .Z(inst3_n2007) );
  XOR2_X1 inst3_U150 ( .A(inst3_n1988), .B(inst3_n2022), .Z(inst3_n1990) );
  XOR2_X1 inst3_U149 ( .A(inst3_n2040), .B(inst3_n1987), .Z(inst3_n2022) );
  XNOR2_X1 inst3_U148 ( .A(inst3_n2063), .B(inst3_n2107), .ZN(inst3_n1992) );
  NOR2_X1 inst3_U147 ( .A1(inst3_n2071), .A2(inst3_n2072), .ZN(inst3_n2107) );
  XOR2_X1 inst3_U146 ( .A(inst3_n2012), .B(inst3_n1986), .Z(inst3_n2072) );
  AND2_X1 inst3_U145 ( .A1(inst3_n1985), .A2(inst3_n2038), .ZN(inst3_n2063) );
  AOI22_X1 inst3_U144 ( .A1(inst3_n1984), .A2(inst3_n1983), .B1(inst3_n2040),
        .B2(inst3_n1982), .ZN(inst3_n2038) );
  INV_X1 inst3_U143 ( .A(inst3_n1981), .ZN(inst3_n1982) );
  XNOR2_X1 inst3_U142 ( .A(inst3_n1980), .B(inst3_n2088), .ZN(inst3_n1993) );
  NAND2_X1 inst3_U141 ( .A1(inst3_n1979), .A2(inst3_n1994), .ZN(inst3_n2088)
         );
  XNOR2_X1 inst3_U140 ( .A(inst3_n1978), .B(inst3_n2013), .ZN(inst3_n1994) );
  XNOR2_X1 inst3_U139 ( .A(inst3_n1977), .B(inst3_n1987), .ZN(inst3_n2013) );
  NAND3_X1 inst3_U138 ( .A1(inst3_n1976), .A2(inst3_n1975), .A3(inst3_n1974),
        .ZN(inst3_n1987) );
  INV_X1 inst3_U137 ( .A(inst3_n1973), .ZN(inst3_n1976) );
  XNOR2_X1 inst3_U136 ( .A(inst3_n2041), .B(inst3_n1972), .ZN(inst3_n1977) );
  XNOR2_X1 inst3_U135 ( .A(inst3_n1971), .B(inst3_n2023), .ZN(inst3_n2041) );
  NOR2_X1 inst3_U134 ( .A1(inst3_n1983), .A2(inst3_n1984), .ZN(inst3_n1971) );
  NAND2_X1 inst3_U133 ( .A1(inst3_n1981), .A2(inst3_n1970), .ZN(inst3_n1984)
         );
  XNOR2_X1 inst3_U132 ( .A(inst3_n2069), .B(inst3_n1969), .ZN(inst3_n1978) );
  NOR2_X1 inst3_U131 ( .A1(inst3_n2009), .A2(inst3_n1968), .ZN(inst3_n1980) );
  XNOR2_X1 inst3_U130 ( .A(inst3_n2014), .B(inst3_n1967), .ZN(inst3_n2009) );
  NAND2_X1 inst3_U129 ( .A1(inst3_n1966), .A2(inst3_n1998), .ZN(inst3_n2052)
         );
  XNOR2_X1 inst3_U128 ( .A(inst3_n1965), .B(inst3_n1964), .ZN(inst3_n1998) );
  XOR2_X1 inst3_U127 ( .A(inst3_n1989), .B(inst3_n2012), .Z(inst3_n1964) );
  XOR2_X1 inst3_U126 ( .A(inst3_n1963), .B(inst3_n1962), .Z(inst3_n2012) );
  OAI211_X1 inst3_U125 ( .C1(inst3_n2040), .C2(inst3_n1970), .A(inst3_n1981),
        .B(inst3_n1961), .ZN(inst3_n1962) );
  NAND2_X1 inst3_U124 ( .A1(inst3_n2040), .A2(inst3_n1970), .ZN(inst3_n1961)
         );
  XNOR2_X1 inst3_U123 ( .A(inst3_n2039), .B(inst3_n2023), .ZN(inst3_n1981) );
  NAND2_X1 inst3_U122 ( .A1(inst3_n2025), .A2(inst3_n2024), .ZN(inst3_n2023)
         );
  XOR2_X1 inst3_U121 ( .A(inst3_n1960), .B(inst3_n1959), .Z(inst3_n2039) );
  XNOR2_X1 inst3_U120 ( .A(inst3_n1958), .B(inst3_n1957), .ZN(inst3_n1960) );
  XNOR2_X1 inst3_U119 ( .A(inst3_n1956), .B(inst3_n1967), .ZN(inst3_n1970) );
  XNOR2_X1 inst3_U118 ( .A(inst3_n1955), .B(inst3_n1954), .ZN(inst3_n1967) );
  XNOR2_X1 inst3_U117 ( .A(inst3_n2015), .B(inst3_n2069), .ZN(inst3_n1955) );
  XNOR2_X1 inst3_U116 ( .A(inst3_n1953), .B(inst3_n2014), .ZN(inst3_n1989) );
  XNOR2_X1 inst3_U115 ( .A(inst3_n1956), .B(inst3_n1952), .ZN(inst3_n2014) );
  AOI211_X1 inst3_U114 ( .C1(inst3_n1975), .C2(inst3_n2040), .A(inst3_n2021),
        .B(inst3_n1951), .ZN(inst3_n1952) );
  NOR2_X1 inst3_U113 ( .A1(inst3_n1975), .A2(inst3_n2040), .ZN(inst3_n1951) );
  INV_X1 inst3_U112 ( .A(inst3_n1974), .ZN(inst3_n2021) );
  XNOR2_X1 inst3_U111 ( .A(inst3_n2069), .B(inst3_n1950), .ZN(inst3_n1974) );
  XNOR2_X1 inst3_U110 ( .A(inst3_n1949), .B(inst3_n1948), .ZN(inst3_n1950) );
  NAND2_X1 inst3_U109 ( .A1(inst3_n1958), .A2(inst3_n1947), .ZN(inst3_n1948)
         );
  XOR2_X1 inst3_U108 ( .A(inst3_n1972), .B(inst3_n1957), .Z(inst3_n1949) );
  NOR2_X1 inst3_U107 ( .A1(inst3_n1983), .A2(inst3_n1973), .ZN(inst3_n2040) );
  XNOR2_X1 inst3_U106 ( .A(inst3_n1946), .B(inst3_n1956), .ZN(inst3_n1973) );
  XNOR2_X1 inst3_U105 ( .A(inst3_n1953), .B(inst3_n1988), .ZN(inst3_n1946) );
  XNOR2_X1 inst3_U104 ( .A(inst3_n1945), .B(inst3_n1944), .ZN(inst3_n1988) );
  INV_X1 inst3_U103 ( .A(inst3_n1943), .ZN(inst3_n1944) );
  XOR2_X1 inst3_U102 ( .A(inst3_n1972), .B(inst3_n1958), .Z(inst3_n1945) );
  NAND2_X1 inst3_U101 ( .A1(inst3_n2018), .A2(inst3_n1947), .ZN(inst3_n1958)
         );
  XOR2_X1 inst3_U100 ( .A(inst3_n1942), .B(inst3_n2048), .Z(inst3_n2018) );
  NAND2_X1 inst3_U99 ( .A1(inst3_n2043), .A2(inst3_n2059), .ZN(inst3_n1972) );
  XNOR2_X1 inst3_U98 ( .A(inst3_n2071), .B(inst3_n1985), .ZN(inst3_n2059) );
  XNOR2_X1 inst3_U97 ( .A(inst3_n1941), .B(inst3_n1940), .ZN(inst3_n2043) );
  XNOR2_X1 inst3_U96 ( .A(inst3_n2025), .B(inst3_n2051), .ZN(inst3_n1941) );
  INV_X1 inst3_U95 ( .A(inst3_n2049), .ZN(inst3_n2051) );
  XNOR2_X1 inst3_U94 ( .A(inst3_n1942), .B(inst3_n1947), .ZN(inst3_n2049) );
  XNOR2_X1 inst3_U93 ( .A(inst3_n1939), .B(inst3_n1938), .ZN(inst3_n1983) );
  XNOR2_X1 inst3_U92 ( .A(inst3_n1937), .B(inst3_n1936), .ZN(inst3_n1939) );
  NAND2_X1 inst3_U91 ( .A1(inst3_n2035), .A2(inst3_n2025), .ZN(inst3_n1936) );
  INV_X1 inst3_U90 ( .A(inst3_n2024), .ZN(inst3_n2035) );
  XOR2_X1 inst3_U89 ( .A(inst3_n2015), .B(inst3_n1935), .Z(inst3_n2024) );
  XNOR2_X1 inst3_U88 ( .A(inst3_n1963), .B(inst3_n1934), .ZN(inst3_n1937) );
  XOR2_X1 inst3_U87 ( .A(inst3_n1933), .B(inst3_n1932), .Z(inst3_n1934) );
  AOI21_X1 inst3_U86 ( .B1(inst3_n2048), .B2(inst3_n1947), .A(inst3_n1931),
        .ZN(inst3_n1932) );
  NOR2_X1 inst3_U85 ( .A1(inst3_n1942), .A2(inst3_n1947), .ZN(inst3_n1931) );
  XOR2_X1 inst3_U84 ( .A(inst3_n1963), .B(inst3_n1986), .Z(inst3_n1975) );
  XNOR2_X1 inst3_U83 ( .A(inst3_n1969), .B(inst3_n1954), .ZN(inst3_n1986) );
  XNOR2_X1 inst3_U82 ( .A(inst3_n1943), .B(inst3_n1957), .ZN(inst3_n1954) );
  NAND2_X1 inst3_U81 ( .A1(inst3_n1979), .A2(inst3_n1995), .ZN(inst3_n1957) );
  XOR2_X1 inst3_U80 ( .A(inst3_n1942), .B(inst3_n1953), .Z(inst3_n1995) );
  XNOR2_X1 inst3_U79 ( .A(inst3_n1930), .B(inst3_n1929), .ZN(inst3_n1979) );
  XOR2_X1 inst3_U78 ( .A(inst3_n1928), .B(inst3_n1947), .Z(inst3_n1930) );
  XNOR2_X1 inst3_U77 ( .A(inst3_n1927), .B(inst3_n1938), .ZN(inst3_n1943) );
  NAND2_X1 inst3_U76 ( .A1(inst3_n1999), .A2(inst3_n1966), .ZN(inst3_n1938) );
  AOI21_X1 inst3_U75 ( .B1(inst3_n1927), .B2(inst3_n1926), .A(inst3_n1925),
        .ZN(inst3_n1969) );
  NOR2_X1 inst3_U74 ( .A1(inst3_n1947), .A2(inst3_n1940), .ZN(inst3_n1925) );
  NAND2_X1 inst3_U73 ( .A1(inst3_n1947), .A2(inst3_n1940), .ZN(inst3_n1926) );
  NAND2_X1 inst3_U72 ( .A1(inst3_n2008), .A2(inst3_n1991), .ZN(inst3_n1963) );
  XOR2_X1 inst3_U71 ( .A(inst3_n2025), .B(inst3_n1953), .Z(inst3_n1991) );
  XOR2_X1 inst3_U70 ( .A(inst3_n2015), .B(inst3_n1927), .Z(inst3_n2008) );
  XNOR2_X1 inst3_U69 ( .A(inst3_n1924), .B(inst3_n1923), .ZN(inst3_n1956) );
  INV_X1 inst3_U68 ( .A(inst3_n1929), .ZN(inst3_n1923) );
  NAND2_X1 inst3_U67 ( .A1(inst3_n2037), .A2(inst3_n1985), .ZN(inst3_n1924) );
  XNOR2_X1 inst3_U66 ( .A(inst3_n1928), .B(inst3_n1922), .ZN(inst3_n1985) );
  INV_X1 inst3_U65 ( .A(inst3_n1999), .ZN(inst3_n1922) );
  XNOR2_X1 inst3_U64 ( .A(inst3_n1942), .B(inst3_n1921), .ZN(inst3_n2037) );
  XNOR2_X1 inst3_U63 ( .A(inst3_n2025), .B(inst3_n1999), .ZN(inst3_n1921) );
  XOR2_X1 inst3_U62 ( .A(inst3_n1953), .B(inst3_n2048), .Z(inst3_n1999) );
  NOR2_X1 inst3_U61 ( .A1(inst3_n2069), .A2(inst3_n1959), .ZN(inst3_n1965) );
  NOR2_X1 inst3_U60 ( .A1(inst3_n2010), .A2(inst3_n1968), .ZN(inst3_n1959) );
  XNOR2_X1 inst3_U59 ( .A(inst3_n1947), .B(inst3_n1940), .ZN(inst3_n1968) );
  XNOR2_X1 inst3_U58 ( .A(inst3_n2015), .B(inst3_n1953), .ZN(inst3_n1947) );
  AOI22_X1 inst3_U57 ( .A1(inst3_n2002), .A2(inst3_n9), .B1(inst3_n2124), .B2(
        inst3_n2800), .ZN(inst3_n1953) );
  AOI22_X1 inst3_U56 ( .A1(inst3_n221), .A2(inst3_n218), .B1(ciphertext3[127]),
        .B2(inst3_n2804), .ZN(inst3_n2124) );
  XNOR2_X1 inst3_U55 ( .A(inst3_n1927), .B(inst3_n1940), .ZN(inst3_n2010) );
  INV_X1 inst3_U54 ( .A(inst3_n1935), .ZN(inst3_n1940) );
  XOR2_X1 inst3_U53 ( .A(inst3_n2071), .B(inst3_n1920), .Z(inst3_n1935) );
  NOR2_X1 inst3_U52 ( .A1(inst3_n2071), .A2(inst3_n2070), .ZN(inst3_n2069) );
  XNOR2_X1 inst3_U51 ( .A(inst3_n2015), .B(inst3_n1929), .ZN(inst3_n2070) );
  XOR2_X1 inst3_U50 ( .A(inst3_n1920), .B(inst3_n2048), .Z(inst3_n1929) );
  AOI22_X1 inst3_U49 ( .A1(inst3_n2002), .A2(inst3_n11), .B1(inst3_n2151),
        .B2(inst3_n2800), .ZN(inst3_n2048) );
  AOI22_X1 inst3_U48 ( .A1(inst3_n223), .A2(inst3_n2802), .B1(ciphertext3[124]), .B2(inst3_n2818), .ZN(inst3_n2151) );
  AOI22_X1 inst3_U47 ( .A1(inst3_n2002), .A2(inst3_n10), .B1(inst3_n2142),
        .B2(inst3_n2800), .ZN(inst3_n2015) );
  AOI22_X1 inst3_U46 ( .A1(inst3_n228), .A2(inst3_n214), .B1(ciphertext3[125]),
        .B2(inst3_n2817), .ZN(inst3_n2142) );
  AOI22_X1 inst3_U45 ( .A1(inst3_n2002), .A2(inst3_n22), .B1(inst3_n2192),
        .B2(inst3_n2800), .ZN(inst3_n2071) );
  AOI22_X1 inst3_U44 ( .A1(inst3_n227), .A2(inst3_n210), .B1(ciphertext3[120]),
        .B2(inst3_n2820), .ZN(inst3_n2192) );
  XOR2_X1 inst3_U43 ( .A(inst3_n1927), .B(inst3_n1920), .Z(inst3_n1966) );
  AOI22_X1 inst3_U42 ( .A1(inst3_n2002), .A2(inst3_n24), .B1(inst3_n2134),
        .B2(inst3_n2800), .ZN(inst3_n1920) );
  AOI22_X1 inst3_U41 ( .A1(inst3_n222), .A2(inst3_n216), .B1(ciphertext3[126]),
        .B2(inst3_n2816), .ZN(inst3_n2134) );
  XOR2_X1 inst3_U40 ( .A(inst3_n1942), .B(inst3_n1928), .Z(inst3_n1927) );
  XOR2_X1 inst3_U39 ( .A(inst3_n2025), .B(inst3_n1933), .Z(inst3_n1928) );
  AOI22_X1 inst3_U38 ( .A1(inst3_n2002), .A2(inst3_n12), .B1(inst3_n2161),
        .B2(inst3_n2800), .ZN(inst3_n1933) );
  AOI22_X1 inst3_U37 ( .A1(inst3_n224), .A2(inst3_n202), .B1(ciphertext3[123]),
        .B2(inst3_n2819), .ZN(inst3_n2161) );
  AOI22_X1 inst3_U36 ( .A1(inst3_n2002), .A2(inst3_n17), .B1(inst3_n2180),
        .B2(inst3_n2800), .ZN(inst3_n2025) );
  AOI22_X1 inst3_U35 ( .A1(inst3_n198), .A2(inst3_n226), .B1(inst3_n2814),
        .B2(ciphertext3[121]), .ZN(inst3_n2180) );
  AOI22_X1 inst3_U34 ( .A1(inst3_n2002), .A2(inst3_n14), .B1(inst3_n2169),
        .B2(inst3_n2800), .ZN(inst3_n1942) );
  AOI22_X1 inst3_U33 ( .A1(ciphertext3[122]), .A2(inst3_n2815), .B1(inst3_n225), .B2(inst3_n2805), .ZN(inst3_n2169) );
  NOR2_X1 inst3_U32 ( .A1(inst3_n1080), .A2(inst3_n321), .ZN(inst3_n2001) );
  AOI22_X1 inst3_U31 ( .A1(inst3_n69), .A2(inst3_n2610), .B1(key3[29]), .B2(
        inst3_n2727), .ZN(inst3_n2006) );
  INV_X1 inst3_U30 ( .A(inst3_n2668), .ZN(inst3_n2610) );
  NAND2_X1 inst3_U29 ( .A1(inst3_n6), .A2(inst3_ctrl_n6), .ZN(inst3_n2800) );
  NAND2_X1 inst3_U28 ( .A1(inst3_n2753), .A2(inst3_n25), .ZN(
        inst3_ctrl_seq4_SFF_0_n5) );
  AOI21_X1 inst3_U27 ( .B1(inst3_n230), .B2(inst3_n1918), .A(inst3_n2774),
        .ZN(inst3_n1919) );
  INV_X1 inst3_U26 ( .A(inst3_n1917), .ZN(inst3_n1918) );
  OAI221_X1 inst3_U25 ( .B1(inst3_n232), .B2(inst3_n1290), .C1(inst3_n1916),
        .C2(inst3_n2756), .A(inst3_n6), .ZN(inst3_ctrl_seq6_SFF_0_n5) );
  INV_X1 inst3_U24 ( .A(inst3_n2720), .ZN(inst3_n2756) );
  NAND2_X1 inst3_U23 ( .A1(inst3_n232), .A2(inst3_n1290), .ZN(inst3_n1916) );
  NAND2_X1 inst3_U22 ( .A1(inst3_n6), .A2(inst3_n231), .ZN(
        inst3_ctrl_seq6_SFF_4_n5) );
  INV_X1 inst3_U21 ( .A(done3), .ZN(inst3_n2720) );
  INV_X1 inst3_U20 ( .A(inst3_n2708), .ZN(done3) );
  INV_X1 inst3_U19 ( .A(inst3_n1914), .ZN(inst3_n2708) );
  OR2_X4 inst3_U18 ( .A1(inst3_ctrl_seq6_SFF_2_n5), .A2(inst3_n1917), .ZN(
        inst3_n2799) );
  NAND4_X1 inst3_U17 ( .A1(inst3_n233), .A2(inst3_n232), .A3(inst3_n1290),
        .A4(inst3_n231), .ZN(inst3_n1917) );
  INV_X1 inst3_U16 ( .A(inst3_n2116), .ZN(inst3_n2123) );
  INV_X1 inst3_U15 ( .A(reset3), .ZN(inst3_n1096) );
  NAND2_X1 inst3_U14 ( .A1(inst3_n6), .A2(inst3_n230), .ZN(
        inst3_ctrl_seq6_SFF_2_n5) );
  INV_X1 inst3_U13 ( .A(inst3_n2775), .ZN(inst3_n2753) );
  NAND2_X1 inst3_U12 ( .A1(inst3_n1919), .A2(inst3_n2800), .ZN(inst3_n2668) );
  NOR4_X1 inst3_U11 ( .A1(inst3_n25), .A2(inst3_n2123), .A3(inst3_n2799), .A4(
        inst3_n2812), .ZN(inst3_n1914) );
  INV_X1 inst3_U10 ( .A(inst3_n6), .ZN(inst3_n2710) );
  NOR4_X1 inst3_U9 ( .A1(inst3_n1081), .A2(inst3_n499), .A3(inst3_n581), .A4(
        inst3_n1080), .ZN(inst3_n2116) );
  NAND2_X1 inst3_U8 ( .A1(inst3_n2002), .A2(inst3_n2799), .ZN(inst3_n2119) );
  INV_X1 inst3_U7 ( .A(inst3_n2800), .ZN(inst3_n2002) );
  INV_X1 inst3_U6 ( .A(inst3_n6), .ZN(inst3_n2727) );
  INV_X2 inst3_U5 ( .A(inst3_n6), .ZN(inst3_n2774) );
  INV_X4 inst3_U4 ( .A(inst3_n1919), .ZN(inst3_n2775) );
  INV_X2 inst3_U3 ( .A(inst3_n2117), .ZN(inst3_n2792) );
  DFF_X2 inst3_nReset_reg_FF_FF ( .D(inst3_n1096), .CK(clk), .Q(inst3_n6),
        .QN(inst3_n2806) );
  DFF_X1 inst3_calcRCon_s_current_state_reg_7__FF_FF ( .D(inst3_calcRCon_n44),
        .CK(clk), .Q(inst3_n2803), .QN(inst3_n1071) );
  DFF_X1 inst3_calcRCon_s_current_state_reg_6__FF_FF ( .D(inst3_calcRCon_n45),
        .CK(clk), .QN(inst3_n718) );
  DFF_X1 inst3_calcRCon_s_current_state_reg_5__FF_FF ( .D(inst3_calcRCon_n46),
        .CK(clk), .QN(inst3_n1080) );
  DFF_X1 inst3_calcRCon_s_current_state_reg_4__FF_FF ( .D(inst3_calcRCon_n47),
        .CK(clk), .QN(inst3_n1081) );
  DFF_X1 inst3_calcRCon_s_current_state_reg_3__FF_FF ( .D(inst3_calcRCon_n48),
        .CK(clk), .Q(inst3_n2813), .QN(inst3_n706) );
  DFF_X1 inst3_calcRCon_s_current_state_reg_2__FF_FF ( .D(inst3_calcRCon_n49),
        .CK(clk), .Q(inst3_n2838), .QN(inst3_n581) );
  DFF_X1 inst3_calcRCon_s_current_state_reg_1__FF_FF ( .D(inst3_calcRCon_n50),
        .CK(clk), .QN(inst3_n499) );
  DFF_X1 inst3_calcRCon_s_current_state_reg_0__FF_FF ( .D(inst3_calcRCon_n51),
        .CK(clk), .Q(inst3_n2839), .QN(inst3_n444) );
  DFF_X1 inst3_KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S33reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst3_n1082) );
  DFF_X1 inst3_KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S33reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst3_n1083) );
  DFF_X1 inst3_KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S33reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst3_n1084) );
  DFF_X1 inst3_KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S33reg_gff_1_SFF_4_n5), .CK(clk), .QN(inst3_n1085) );
  DFF_X1 inst3_KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S33reg_gff_1_SFF_3_n5), .CK(clk), .QN(inst3_n1086) );
  DFF_X1 inst3_KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S33reg_gff_1_SFF_2_n5), .CK(clk), .QN(inst3_n1087) );
  DFF_X1 inst3_KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S33reg_gff_1_SFF_1_n5), .CK(clk), .Q(inst3_n57) );
  DFF_X1 inst3_KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S33reg_gff_1_SFF_0_n5), .CK(clk), .QN(inst3_n1089) );
  DFF_X1 inst3_KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S32reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst3_n1090) );
  DFF_X1 inst3_KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S32reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst3_n1091) );
  DFF_X1 inst3_KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S32reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst3_n1092) );
  DFF_X1 inst3_KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S32reg_gff_1_SFF_4_n6), .CK(clk), .QN(inst3_n1093) );
  DFF_X1 inst3_KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S32reg_gff_1_SFF_3_n6), .CK(clk), .QN(inst3_n1094) );
  DFF_X1 inst3_KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S32reg_gff_1_SFF_2_n6), .CK(clk), .QN(inst3_n1095) );
  DFF_X1 inst3_KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S32reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst3_n65) );
  DFF_X1 inst3_KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S32reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst3_n1097) );
  DFF_X1 inst3_KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S31reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst3_n67) );
  DFF_X1 inst3_KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S31reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst3_n68) );
  DFF_X1 inst3_KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S31reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst3_n69) );
  DFF_X1 inst3_KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S31reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst3_n70), .QN(
        inst3_n2837) );
  DFF_X1 inst3_KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S31reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst3_n71) );
  DFF_X1 inst3_KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S31reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst3_n72) );
  DFF_X1 inst3_KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S31reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst3_n73) );
  DFF_X1 inst3_KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S31reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst3_n74) );
  DFF_X1 inst3_KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S30reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst3_n75), .QN(
        inst3_n2860) );
  DFF_X1 inst3_KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S30reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst3_n76), .QN(
        inst3_n2863) );
  DFF_X1 inst3_KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S30reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst3_n77), .QN(
        inst3_n2858) );
  DFF_X1 inst3_KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S30reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst3_n78) );
  DFF_X1 inst3_KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S30reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst3_n79), .QN(
        inst3_n2864) );
  DFF_X1 inst3_KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S30reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst3_n80), .QN(
        inst3_n2861) );
  DFF_X1 inst3_KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S30reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst3_n81), .QN(
        inst3_n2862) );
  DFF_X1 inst3_KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S30reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst3_n82), .QN(
        inst3_n2859) );
  DFF_X1 inst3_KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S23reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst3_n83) );
  DFF_X1 inst3_KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S23reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst3_n84) );
  DFF_X1 inst3_KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S23reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst3_n85) );
  DFF_X1 inst3_KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S23reg_gff_1_SFF_4_n5), .CK(clk), .Q(inst3_n86) );
  DFF_X1 inst3_KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S23reg_gff_1_SFF_3_n5), .CK(clk), .Q(inst3_n87) );
  DFF_X1 inst3_KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S23reg_gff_1_SFF_2_n5), .CK(clk), .Q(inst3_n88) );
  DFF_X1 inst3_KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S23reg_gff_1_SFF_1_n5), .CK(clk), .Q(inst3_n89) );
  DFF_X1 inst3_KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S23reg_gff_1_SFF_0_n5), .CK(clk), .Q(inst3_n90) );
  DFF_X1 inst3_KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S22reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst3_n91) );
  DFF_X1 inst3_KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S22reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst3_n92) );
  DFF_X1 inst3_KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S22reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst3_n93) );
  DFF_X1 inst3_KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S22reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst3_n94) );
  DFF_X1 inst3_KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S22reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst3_n95) );
  DFF_X1 inst3_KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S22reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst3_n96) );
  DFF_X1 inst3_KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S22reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst3_n97) );
  DFF_X1 inst3_KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S22reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst3_n98) );
  DFF_X1 inst3_KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S21reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst3_n107) );
  DFF_X1 inst3_KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S21reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst3_n108) );
  DFF_X1 inst3_KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S21reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst3_n109) );
  DFF_X1 inst3_KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S21reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst3_n110) );
  DFF_X1 inst3_KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S21reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst3_n111) );
  DFF_X1 inst3_KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S21reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst3_n112) );
  DFF_X1 inst3_KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S21reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst3_n113) );
  DFF_X1 inst3_KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S21reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst3_n114) );
  DFF_X1 inst3_KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S20reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst3_n115) );
  DFF_X1 inst3_KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S20reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst3_n116) );
  DFF_X1 inst3_KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S20reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst3_n117) );
  DFF_X1 inst3_KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S20reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst3_n118) );
  DFF_X1 inst3_KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S20reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst3_n119) );
  DFF_X1 inst3_KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S20reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst3_n120) );
  DFF_X1 inst3_KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S20reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst3_n121) );
  DFF_X1 inst3_KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S20reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst3_n122), .QN(
        inst3_n2865) );
  DFF_X1 inst3_KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S13reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst3_n9), .QN(
        inst3_n2850) );
  DFF_X1 inst3_KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S13reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst3_n24), .QN(
        inst3_n2851) );
  DFF_X1 inst3_KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S13reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst3_n10), .QN(
        inst3_n2852) );
  DFF_X1 inst3_KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S13reg_gff_1_SFF_4_n5), .CK(clk), .Q(inst3_n11), .QN(
        inst3_n2853) );
  DFF_X1 inst3_KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S13reg_gff_1_SFF_3_n5), .CK(clk), .Q(inst3_n12), .QN(
        inst3_n2854) );
  DFF_X1 inst3_KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S13reg_gff_1_SFF_2_n5), .CK(clk), .Q(inst3_n14), .QN(
        inst3_n2855) );
  DFF_X1 inst3_KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S13reg_gff_1_SFF_1_n5), .CK(clk), .Q(inst3_n17), .QN(
        inst3_n2856) );
  DFF_X1 inst3_KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S13reg_gff_1_SFF_0_n5), .CK(clk), .Q(inst3_n22), .QN(
        inst3_n2857) );
  DFF_X1 inst3_KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S12reg_gff_1_SFF_7_n5), .CK(clk), .Q(inst3_n123), .QN(
        inst3_n2866) );
  DFF_X1 inst3_KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S12reg_gff_1_SFF_6_n5), .CK(clk), .Q(inst3_n124), .QN(
        inst3_n2867) );
  DFF_X1 inst3_KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S12reg_gff_1_SFF_5_n5), .CK(clk), .Q(inst3_n125), .QN(
        inst3_n2868) );
  DFF_X1 inst3_KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S12reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst3_n126), .QN(
        inst3_n2869) );
  DFF_X1 inst3_KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S12reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst3_n127), .QN(
        inst3_n2870) );
  DFF_X1 inst3_KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S12reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst3_n128), .QN(
        inst3_n2871) );
  DFF_X1 inst3_KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S12reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst3_n129), .QN(
        inst3_n2872) );
  DFF_X1 inst3_KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S12reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst3_n130), .QN(
        inst3_n2873) );
  DFF_X1 inst3_KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S11reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst3_n131) );
  DFF_X1 inst3_KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S11reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst3_n132) );
  DFF_X1 inst3_KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S11reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst3_n133) );
  DFF_X1 inst3_KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S11reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst3_n134) );
  DFF_X1 inst3_KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S11reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst3_n135) );
  DFF_X1 inst3_KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S11reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst3_n136) );
  DFF_X1 inst3_KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S11reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst3_n137) );
  DFF_X1 inst3_KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S11reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst3_n1161) );
  DFF_X1 inst3_KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S10reg_gff_1_SFF_7_n6), .CK(clk), .QN(inst3_n1162) );
  DFF_X1 inst3_KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S10reg_gff_1_SFF_6_n6), .CK(clk), .QN(inst3_n1163) );
  DFF_X1 inst3_KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S10reg_gff_1_SFF_5_n6), .CK(clk), .QN(inst3_n1164) );
  DFF_X1 inst3_KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S10reg_gff_1_SFF_4_n6), .CK(clk), .QN(inst3_n1165) );
  DFF_X1 inst3_KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S10reg_gff_1_SFF_3_n6), .CK(clk), .QN(inst3_n1166) );
  DFF_X1 inst3_KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S10reg_gff_1_SFF_2_n6), .CK(clk), .QN(inst3_n1167) );
  DFF_X1 inst3_KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S10reg_gff_1_SFF_1_n6), .CK(clk), .QN(inst3_n1168) );
  DFF_X1 inst3_KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S10reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst3_n1169) );
  DFF_X1 inst3_KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S03reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst3_n1170) );
  DFF_X1 inst3_KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S03reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst3_n1171) );
  DFF_X1 inst3_KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S03reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst3_n1172) );
  DFF_X1 inst3_KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S03reg_gff_1_SFF_4_n5), .CK(clk), .QN(inst3_n1173) );
  DFF_X1 inst3_KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S03reg_gff_1_SFF_3_n5), .CK(clk), .QN(inst3_n1174) );
  DFF_X1 inst3_KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S03reg_gff_1_SFF_2_n5), .CK(clk), .QN(inst3_n1175) );
  DFF_X1 inst3_KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S03reg_gff_1_SFF_1_n5), .CK(clk), .QN(inst3_n1176) );
  DFF_X1 inst3_KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S03reg_gff_1_SFF_0_n5), .CK(clk), .QN(inst3_n1177) );
  DFF_X1 inst3_KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S02reg_gff_1_SFF_7_n5), .CK(clk), .QN(inst3_n1178) );
  DFF_X1 inst3_KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S02reg_gff_1_SFF_6_n5), .CK(clk), .QN(inst3_n1179) );
  DFF_X1 inst3_KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S02reg_gff_1_SFF_5_n5), .CK(clk), .QN(inst3_n1180) );
  DFF_X1 inst3_KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S02reg_gff_1_SFF_4_n6), .CK(clk), .QN(inst3_n1181) );
  DFF_X1 inst3_KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S02reg_gff_1_SFF_3_n6), .CK(clk), .QN(inst3_n1182) );
  DFF_X1 inst3_KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S02reg_gff_1_SFF_2_n6), .CK(clk), .QN(inst3_n1183) );
  DFF_X1 inst3_KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S02reg_gff_1_SFF_1_n6), .CK(clk), .QN(inst3_n1184) );
  DFF_X1 inst3_KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S02reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst3_n1185) );
  DFF_X1 inst3_KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S01reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst3_n2824), .QN(
        inst3_n1186) );
  DFF_X1 inst3_KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S01reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst3_n2825), .QN(
        inst3_n1187) );
  DFF_X1 inst3_KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S01reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst3_n2826), .QN(
        inst3_n1188) );
  DFF_X1 inst3_KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S01reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst3_n2840), .QN(
        inst3_n1189) );
  DFF_X1 inst3_KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S01reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst3_n2827), .QN(
        inst3_n1190) );
  DFF_X1 inst3_KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S01reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst3_n2828), .QN(
        inst3_n1191) );
  DFF_X1 inst3_KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S01reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst3_n2841), .QN(
        inst3_n1192) );
  DFF_X1 inst3_KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S01reg_gff_1_SFF_0_n6), .CK(clk), .QN(inst3_n1193) );
  DFF_X1 inst3_KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S00reg_gff_1_SFF_7_n6), .CK(clk), .Q(inst3_n2804), .QN(
        inst3_n221) );
  DFF_X1 inst3_KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S00reg_gff_1_SFF_6_n6), .CK(clk), .Q(inst3_n2816), .QN(
        inst3_n222) );
  DFF_X1 inst3_KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S00reg_gff_1_SFF_5_n6), .CK(clk), .Q(inst3_n2817), .QN(
        inst3_n228) );
  DFF_X1 inst3_KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S00reg_gff_1_SFF_4_n6), .CK(clk), .Q(inst3_n2818), .QN(
        inst3_n223) );
  DFF_X1 inst3_KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S00reg_gff_1_SFF_3_n6), .CK(clk), .Q(inst3_n2819), .QN(
        inst3_n224) );
  DFF_X1 inst3_KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S00reg_gff_1_SFF_2_n6), .CK(clk), .Q(inst3_n2815), .QN(
        inst3_n225) );
  DFF_X1 inst3_KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S00reg_gff_1_SFF_1_n6), .CK(clk), .Q(inst3_n2814), .QN(
        inst3_n226) );
  DFF_X1 inst3_KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_KeyArray_S00reg_gff_1_SFF_0_n6), .CK(clk), .Q(inst3_n2820), .QN(
        inst3_n227) );
  DFF_X1 inst3_stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S33reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext3[7]),
        .QN(inst3_n1194) );
  DFF_X1 inst3_stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S33reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext3[6]),
        .QN(inst3_n1195) );
  DFF_X1 inst3_stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S33reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext3[5]),
        .QN(inst3_n1196) );
  DFF_X1 inst3_stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S33reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext3[4]),
        .QN(inst3_n1197) );
  DFF_X1 inst3_stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S33reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext3[3]),
        .QN(inst3_n1198) );
  DFF_X1 inst3_stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S33reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext3[2]),
        .QN(inst3_n1199) );
  DFF_X1 inst3_stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S33reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext3[1]),
        .QN(inst3_n1200) );
  DFF_X1 inst3_stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S33reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext3[0]),
        .QN(inst3_n1201) );
  DFF_X1 inst3_stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S32reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext3[15]),
        .QN(inst3_n1202) );
  DFF_X1 inst3_stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S32reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext3[14]),
        .QN(inst3_n1203) );
  DFF_X1 inst3_stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S32reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext3[13]),
        .QN(inst3_n1204) );
  DFF_X1 inst3_stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S32reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[12]),
        .QN(inst3_n1205) );
  DFF_X1 inst3_stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S32reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[11]),
        .QN(inst3_n1206) );
  DFF_X1 inst3_stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S32reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[10]),
        .QN(inst3_n1207) );
  DFF_X1 inst3_stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S32reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[9]),
        .QN(inst3_n1208) );
  DFF_X1 inst3_stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S32reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[8]),
        .QN(inst3_n1209) );
  DFF_X1 inst3_stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S31reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext3[23]),
        .QN(inst3_n2830) );
  DFF_X1 inst3_stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S31reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext3[22]),
        .QN(inst3_n2829) );
  DFF_X1 inst3_stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S31reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext3[21]),
        .QN(inst3_n2831) );
  DFF_X1 inst3_stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S31reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[20]),
        .QN(inst3_n2832) );
  DFF_X1 inst3_stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S31reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[19]),
        .QN(inst3_n2833) );
  DFF_X1 inst3_stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S31reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[18]),
        .QN(inst3_n2834) );
  DFF_X1 inst3_stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S31reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[17]),
        .QN(inst3_n2835) );
  DFF_X1 inst3_stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S31reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[16]),
        .QN(inst3_n2836) );
  DFF_X1 inst3_stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S30reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext3[31]),
        .QN(inst3_n2808) );
  DFF_X1 inst3_stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S30reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext3[30]),
        .QN(inst3_n215) );
  DFF_X1 inst3_stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S30reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext3[29]),
        .QN(inst3_n2807) );
  DFF_X1 inst3_stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S30reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext3[28]),
        .QN(inst3_n207) );
  DFF_X1 inst3_stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S30reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext3[27]),
        .QN(inst3_n2821) );
  DFF_X1 inst3_stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S30reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext3[26]),
        .QN(inst3_n203) );
  DFF_X1 inst3_stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S30reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext3[25]),
        .QN(inst3_n191) );
  DFF_X1 inst3_stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S30reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext3[24]),
        .QN(inst3_n199) );
  DFF_X1 inst3_stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S23reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext3[39]),
        .QN(inst3_n1218) );
  DFF_X1 inst3_stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S23reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext3[38]),
        .QN(inst3_n1219) );
  DFF_X1 inst3_stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S23reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext3[37]),
        .QN(inst3_n1220) );
  DFF_X1 inst3_stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S23reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[36]),
        .QN(inst3_n1221) );
  DFF_X1 inst3_stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S23reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[35]),
        .QN(inst3_n1222) );
  DFF_X1 inst3_stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S23reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[34]),
        .QN(inst3_n1223) );
  DFF_X1 inst3_stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S23reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[33]),
        .QN(inst3_n1224) );
  DFF_X1 inst3_stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S23reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[32]),
        .QN(inst3_n1225) );
  DFF_X1 inst3_stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S22reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext3[47]),
        .QN(inst3_n1226) );
  DFF_X1 inst3_stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S22reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext3[46]),
        .QN(inst3_n1227) );
  DFF_X1 inst3_stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S22reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext3[45]),
        .QN(inst3_n1228) );
  DFF_X1 inst3_stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S22reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[44]),
        .QN(inst3_n1229) );
  DFF_X1 inst3_stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S22reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[43]),
        .QN(inst3_n1230) );
  DFF_X1 inst3_stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S22reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[42]),
        .QN(inst3_n1231) );
  DFF_X1 inst3_stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S22reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[41]),
        .QN(inst3_n1232) );
  DFF_X1 inst3_stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S22reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[40]),
        .QN(inst3_n1233) );
  DFF_X1 inst3_stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S21reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext3[55])
         );
  DFF_X1 inst3_stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S21reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext3[54])
         );
  DFF_X1 inst3_stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S21reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext3[53])
         );
  DFF_X1 inst3_stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S21reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[52])
         );
  DFF_X1 inst3_stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S21reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[51])
         );
  DFF_X1 inst3_stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S21reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[50])
         );
  DFF_X1 inst3_stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S21reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[49])
         );
  DFF_X1 inst3_stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S21reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[48])
         );
  DFF_X1 inst3_stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S20reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext3[63]),
        .QN(inst3_n219) );
  DFF_X1 inst3_stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S20reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext3[62]),
        .QN(inst3_n2809) );
  DFF_X1 inst3_stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S20reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext3[61]),
        .QN(inst3_n2823) );
  DFF_X1 inst3_stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S20reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext3[60]),
        .QN(inst3_n2822) );
  DFF_X1 inst3_stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S20reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext3[59]),
        .QN(inst3_n196) );
  DFF_X1 inst3_stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S20reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext3[58]),
        .QN(inst3_n193) );
  DFF_X1 inst3_stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S20reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext3[57]),
        .QN(inst3_n2811) );
  DFF_X1 inst3_stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S20reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext3[56]),
        .QN(inst3_n2810) );
  DFF_X1 inst3_stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S13reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext3[71])
         );
  DFF_X1 inst3_stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S13reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext3[70])
         );
  DFF_X1 inst3_stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S13reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext3[69])
         );
  DFF_X1 inst3_stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S13reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[68])
         );
  DFF_X1 inst3_stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S13reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[67])
         );
  DFF_X1 inst3_stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S13reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[66])
         );
  DFF_X1 inst3_stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S13reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[65])
         );
  DFF_X1 inst3_stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S13reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[64])
         );
  DFF_X1 inst3_stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S12reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext3[79]),
        .QN(inst3_n1250) );
  DFF_X1 inst3_stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S12reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext3[78]),
        .QN(inst3_n1251) );
  DFF_X1 inst3_stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S12reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext3[77]),
        .QN(inst3_n1252) );
  DFF_X1 inst3_stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S12reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[76]),
        .QN(inst3_n1253) );
  DFF_X1 inst3_stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S12reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[75]),
        .QN(inst3_n1254) );
  DFF_X1 inst3_stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S12reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[74]),
        .QN(inst3_n1255) );
  DFF_X1 inst3_stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S12reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[73]),
        .QN(inst3_n1256) );
  DFF_X1 inst3_stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S12reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[72]),
        .QN(inst3_n1257) );
  DFF_X1 inst3_stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S11reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext3[87]),
        .QN(inst3_n1258) );
  DFF_X1 inst3_stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S11reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext3[86]),
        .QN(inst3_n1259) );
  DFF_X1 inst3_stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S11reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext3[85]),
        .QN(inst3_n1260) );
  DFF_X1 inst3_stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S11reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[84]),
        .QN(inst3_n1261) );
  DFF_X1 inst3_stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S11reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[83]),
        .QN(inst3_n1262) );
  DFF_X1 inst3_stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S11reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[82]),
        .QN(inst3_n1263) );
  DFF_X1 inst3_stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S11reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[81]),
        .QN(inst3_n1264) );
  DFF_X1 inst3_stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S11reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[80]),
        .QN(inst3_n1265) );
  DFF_X1 inst3_stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S10reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext3[95]),
        .QN(inst3_n220) );
  DFF_X1 inst3_stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S10reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext3[94]),
        .QN(inst3_n206) );
  DFF_X1 inst3_stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S10reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext3[93]),
        .QN(inst3_n190) );
  DFF_X1 inst3_stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S10reg_gff_1_SFF_4_n5), .CK(clk), .Q(ciphertext3[92]),
        .QN(inst3_n212) );
  DFF_X1 inst3_stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S10reg_gff_1_SFF_3_n5), .CK(clk), .Q(ciphertext3[91]),
        .QN(inst3_n201) );
  DFF_X1 inst3_stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S10reg_gff_1_SFF_2_n5), .CK(clk), .Q(ciphertext3[90]),
        .QN(inst3_n194) );
  DFF_X1 inst3_stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S10reg_gff_1_SFF_1_n5), .CK(clk), .Q(ciphertext3[89]),
        .QN(inst3_n197) );
  DFF_X1 inst3_stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S10reg_gff_1_SFF_0_n5), .CK(clk), .Q(ciphertext3[88]),
        .QN(inst3_n209) );
  DFF_X1 inst3_stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S03reg_gff_1_SFF_7_n5), .CK(clk), .Q(ciphertext3[103]), .QN(inst3_n1266) );
  DFF_X1 inst3_stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S03reg_gff_1_SFF_6_n5), .CK(clk), .Q(ciphertext3[102]), .QN(inst3_n1267) );
  DFF_X1 inst3_stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S03reg_gff_1_SFF_5_n5), .CK(clk), .Q(ciphertext3[101]), .QN(inst3_n1268) );
  DFF_X1 inst3_stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S03reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[100]), .QN(inst3_n1269) );
  DFF_X1 inst3_stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S03reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[99]),
        .QN(inst3_n1270) );
  DFF_X1 inst3_stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S03reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[98]),
        .QN(inst3_n1271) );
  DFF_X1 inst3_stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S03reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[97]),
        .QN(inst3_n1272) );
  DFF_X1 inst3_stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S03reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[96]),
        .QN(inst3_n1273) );
  DFF_X1 inst3_stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S02reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext3[111]) );
  DFF_X1 inst3_stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S02reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext3[110]) );
  DFF_X1 inst3_stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S02reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext3[109]) );
  DFF_X1 inst3_stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S02reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[108]) );
  DFF_X1 inst3_stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S02reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[107]) );
  DFF_X1 inst3_stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S02reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[106]) );
  DFF_X1 inst3_stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S02reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[105]) );
  DFF_X1 inst3_stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S02reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[104]) );
  DFF_X1 inst3_stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S01reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext3[119]), .QN(inst3_n2842) );
  DFF_X1 inst3_stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S01reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext3[118]), .QN(inst3_n2843) );
  DFF_X1 inst3_stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S01reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext3[117]), .QN(inst3_n2844) );
  DFF_X1 inst3_stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S01reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[116]), .QN(inst3_n2845) );
  DFF_X1 inst3_stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S01reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[115]), .QN(inst3_n2846) );
  DFF_X1 inst3_stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S01reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[114]), .QN(inst3_n2847) );
  DFF_X1 inst3_stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S01reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[113]), .QN(inst3_n2848) );
  DFF_X1 inst3_stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S01reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[112]), .QN(inst3_n2849) );
  DFF_X1 inst3_stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        inst3_stateArray_S00reg_gff_1_SFF_7_n6), .CK(clk), .Q(ciphertext3[127]), .QN(inst3_n218) );
  DFF_X1 inst3_stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        inst3_stateArray_S00reg_gff_1_SFF_6_n6), .CK(clk), .Q(ciphertext3[126]), .QN(inst3_n216) );
  DFF_X1 inst3_stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        inst3_stateArray_S00reg_gff_1_SFF_5_n6), .CK(clk), .Q(ciphertext3[125]), .QN(inst3_n214) );
  DFF_X1 inst3_stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        inst3_stateArray_S00reg_gff_1_SFF_4_n6), .CK(clk), .Q(ciphertext3[124]), .QN(inst3_n2802) );
  DFF_X1 inst3_stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        inst3_stateArray_S00reg_gff_1_SFF_3_n6), .CK(clk), .Q(ciphertext3[123]), .QN(inst3_n202) );
  DFF_X1 inst3_stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        inst3_stateArray_S00reg_gff_1_SFF_2_n6), .CK(clk), .Q(ciphertext3[122]), .QN(inst3_n2805) );
  DFF_X1 inst3_stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        inst3_stateArray_S00reg_gff_1_SFF_1_n6), .CK(clk), .Q(ciphertext3[121]), .QN(inst3_n198) );
  DFF_X1 inst3_stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        inst3_stateArray_S00reg_gff_1_SFF_0_n6), .CK(clk), .Q(ciphertext3[120]), .QN(inst3_n210) );
  DFF_X1 inst3_ctrl_CSenRC_reg_FF_FF ( .D(inst3_n2543), .CK(clk), .QN(
        inst3_n321) );
  DFF_X1 inst3_ctrl_CSselMC_reg_FF_FF ( .D(inst3_n1088), .CK(clk), .Q(
        inst3_ctrl_n6) );
  DFF_X1 inst3_ctrl_seq4_SFF_1_Q_reg_FF_FF ( .D(inst3_ctrl_seq4_SFF_1_n5),
        .CK(clk), .Q(inst3_n25) );
  DFF_X1 inst3_ctrl_seq4_SFF_0_Q_reg_FF_FF ( .D(inst3_ctrl_seq4_SFF_0_n5),
        .CK(clk), .Q(inst3_n143), .QN(inst3_n2812) );
  DFF_X1 inst3_ctrl_seq6_SFF_4_Q_reg_FF_FF ( .D(inst3_ctrl_seq6_SFF_4_n5),
        .CK(clk), .QN(inst3_n1290) );
  DFF_X1 inst3_ctrl_seq6_SFF_3_Q_reg_FF_FF ( .D(inst3_ctrl_seq6_SFF_3_n5),
        .CK(clk), .QN(inst3_n231) );
  DFF_X1 inst3_ctrl_seq6_SFF_2_Q_reg_FF_FF ( .D(inst3_ctrl_seq6_SFF_2_n5),
        .CK(clk), .QN(inst3_n233) );
  DFF_X1 inst3_ctrl_seq6_SFF_1_Q_reg_FF_FF ( .D(inst3_ctrl_seq6_SFF_1_n5),
        .CK(clk), .QN(inst3_n230) );
  DFF_X1 inst3_ctrl_seq6_SFF_0_Q_reg_FF_FF ( .D(inst3_ctrl_seq6_SFF_0_n5),
        .CK(clk), .QN(inst3_n232) );
  NAND2_X1 mv_0_U384 ( .A1(mv_0_n256), .A2(mv_0_n255), .ZN(ciphertext[127]) );
  NAND2_X1 mv_0_U383 ( .A1(ciphertext3[127]), .A2(ciphertext1[127]), .ZN(
        mv_0_n255) );
  OAI21_X1 mv_0_U382 ( .B1(ciphertext3[127]), .B2(ciphertext1[127]), .A(
        ciphertext2[127]), .ZN(mv_0_n256) );
  NAND2_X1 mv_0_U381 ( .A1(mv_0_n254), .A2(mv_0_n253), .ZN(ciphertext[126]) );
  NAND2_X1 mv_0_U380 ( .A1(ciphertext3[126]), .A2(ciphertext1[126]), .ZN(
        mv_0_n253) );
  OAI21_X1 mv_0_U379 ( .B1(ciphertext3[126]), .B2(ciphertext1[126]), .A(
        ciphertext2[126]), .ZN(mv_0_n254) );
  NAND2_X1 mv_0_U378 ( .A1(mv_0_n252), .A2(mv_0_n251), .ZN(ciphertext[125]) );
  NAND2_X1 mv_0_U377 ( .A1(ciphertext3[125]), .A2(ciphertext1[125]), .ZN(
        mv_0_n251) );
  OAI21_X1 mv_0_U376 ( .B1(ciphertext3[125]), .B2(ciphertext1[125]), .A(
        ciphertext2[125]), .ZN(mv_0_n252) );
  NAND2_X1 mv_0_U375 ( .A1(mv_0_n250), .A2(mv_0_n249), .ZN(ciphertext[124]) );
  NAND2_X1 mv_0_U374 ( .A1(ciphertext3[124]), .A2(ciphertext1[124]), .ZN(
        mv_0_n249) );
  OAI21_X1 mv_0_U373 ( .B1(ciphertext3[124]), .B2(ciphertext1[124]), .A(
        ciphertext2[124]), .ZN(mv_0_n250) );
  NAND2_X1 mv_0_U372 ( .A1(mv_0_n248), .A2(mv_0_n247), .ZN(ciphertext[123]) );
  NAND2_X1 mv_0_U371 ( .A1(ciphertext3[123]), .A2(ciphertext1[123]), .ZN(
        mv_0_n247) );
  OAI21_X1 mv_0_U370 ( .B1(ciphertext3[123]), .B2(ciphertext1[123]), .A(
        ciphertext2[123]), .ZN(mv_0_n248) );
  NAND2_X1 mv_0_U369 ( .A1(mv_0_n246), .A2(mv_0_n245), .ZN(ciphertext[122]) );
  NAND2_X1 mv_0_U368 ( .A1(ciphertext3[122]), .A2(ciphertext1[122]), .ZN(
        mv_0_n245) );
  OAI21_X1 mv_0_U367 ( .B1(ciphertext3[122]), .B2(ciphertext1[122]), .A(
        ciphertext2[122]), .ZN(mv_0_n246) );
  NAND2_X1 mv_0_U366 ( .A1(mv_0_n244), .A2(mv_0_n243), .ZN(ciphertext[121]) );
  NAND2_X1 mv_0_U365 ( .A1(ciphertext3[121]), .A2(ciphertext1[121]), .ZN(
        mv_0_n243) );
  OAI21_X1 mv_0_U364 ( .B1(ciphertext3[121]), .B2(ciphertext1[121]), .A(
        ciphertext2[121]), .ZN(mv_0_n244) );
  NAND2_X1 mv_0_U363 ( .A1(mv_0_n242), .A2(mv_0_n241), .ZN(ciphertext[120]) );
  NAND2_X1 mv_0_U362 ( .A1(ciphertext3[120]), .A2(ciphertext1[120]), .ZN(
        mv_0_n241) );
  OAI21_X1 mv_0_U361 ( .B1(ciphertext3[120]), .B2(ciphertext1[120]), .A(
        ciphertext2[120]), .ZN(mv_0_n242) );
  NAND2_X1 mv_0_U360 ( .A1(mv_0_n240), .A2(mv_0_n239), .ZN(ciphertext[119]) );
  NAND2_X1 mv_0_U359 ( .A1(ciphertext3[119]), .A2(ciphertext1[119]), .ZN(
        mv_0_n239) );
  OAI21_X1 mv_0_U358 ( .B1(ciphertext3[119]), .B2(ciphertext1[119]), .A(
        ciphertext2[119]), .ZN(mv_0_n240) );
  NAND2_X1 mv_0_U357 ( .A1(mv_0_n238), .A2(mv_0_n237), .ZN(ciphertext[118]) );
  NAND2_X1 mv_0_U356 ( .A1(ciphertext3[118]), .A2(ciphertext1[118]), .ZN(
        mv_0_n237) );
  OAI21_X1 mv_0_U355 ( .B1(ciphertext3[118]), .B2(ciphertext1[118]), .A(
        ciphertext2[118]), .ZN(mv_0_n238) );
  NAND2_X1 mv_0_U354 ( .A1(mv_0_n236), .A2(mv_0_n235), .ZN(ciphertext[117]) );
  NAND2_X1 mv_0_U353 ( .A1(ciphertext3[117]), .A2(ciphertext1[117]), .ZN(
        mv_0_n235) );
  OAI21_X1 mv_0_U352 ( .B1(ciphertext3[117]), .B2(ciphertext1[117]), .A(
        ciphertext2[117]), .ZN(mv_0_n236) );
  NAND2_X1 mv_0_U351 ( .A1(mv_0_n234), .A2(mv_0_n233), .ZN(ciphertext[116]) );
  NAND2_X1 mv_0_U350 ( .A1(ciphertext3[116]), .A2(ciphertext1[116]), .ZN(
        mv_0_n233) );
  OAI21_X1 mv_0_U349 ( .B1(ciphertext3[116]), .B2(ciphertext1[116]), .A(
        ciphertext2[116]), .ZN(mv_0_n234) );
  NAND2_X1 mv_0_U348 ( .A1(mv_0_n232), .A2(mv_0_n231), .ZN(ciphertext[115]) );
  NAND2_X1 mv_0_U347 ( .A1(ciphertext3[115]), .A2(ciphertext1[115]), .ZN(
        mv_0_n231) );
  OAI21_X1 mv_0_U346 ( .B1(ciphertext3[115]), .B2(ciphertext1[115]), .A(
        ciphertext2[115]), .ZN(mv_0_n232) );
  NAND2_X1 mv_0_U345 ( .A1(mv_0_n230), .A2(mv_0_n229), .ZN(ciphertext[114]) );
  NAND2_X1 mv_0_U344 ( .A1(ciphertext3[114]), .A2(ciphertext1[114]), .ZN(
        mv_0_n229) );
  OAI21_X1 mv_0_U343 ( .B1(ciphertext3[114]), .B2(ciphertext1[114]), .A(
        ciphertext2[114]), .ZN(mv_0_n230) );
  NAND2_X1 mv_0_U342 ( .A1(mv_0_n228), .A2(mv_0_n227), .ZN(ciphertext[113]) );
  NAND2_X1 mv_0_U341 ( .A1(ciphertext3[113]), .A2(ciphertext1[113]), .ZN(
        mv_0_n227) );
  OAI21_X1 mv_0_U340 ( .B1(ciphertext3[113]), .B2(ciphertext1[113]), .A(
        ciphertext2[113]), .ZN(mv_0_n228) );
  NAND2_X1 mv_0_U339 ( .A1(mv_0_n226), .A2(mv_0_n225), .ZN(ciphertext[112]) );
  NAND2_X1 mv_0_U338 ( .A1(ciphertext3[112]), .A2(ciphertext1[112]), .ZN(
        mv_0_n225) );
  OAI21_X1 mv_0_U337 ( .B1(ciphertext3[112]), .B2(ciphertext1[112]), .A(
        ciphertext2[112]), .ZN(mv_0_n226) );
  NAND2_X1 mv_0_U336 ( .A1(mv_0_n224), .A2(mv_0_n223), .ZN(ciphertext[111]) );
  NAND2_X1 mv_0_U335 ( .A1(ciphertext3[111]), .A2(ciphertext1[111]), .ZN(
        mv_0_n223) );
  OAI21_X1 mv_0_U334 ( .B1(ciphertext3[111]), .B2(ciphertext1[111]), .A(
        ciphertext2[111]), .ZN(mv_0_n224) );
  NAND2_X1 mv_0_U333 ( .A1(mv_0_n222), .A2(mv_0_n221), .ZN(ciphertext[110]) );
  NAND2_X1 mv_0_U332 ( .A1(ciphertext3[110]), .A2(ciphertext1[110]), .ZN(
        mv_0_n221) );
  OAI21_X1 mv_0_U331 ( .B1(ciphertext3[110]), .B2(ciphertext1[110]), .A(
        ciphertext2[110]), .ZN(mv_0_n222) );
  NAND2_X1 mv_0_U330 ( .A1(mv_0_n220), .A2(mv_0_n219), .ZN(ciphertext[109]) );
  NAND2_X1 mv_0_U329 ( .A1(ciphertext3[109]), .A2(ciphertext1[109]), .ZN(
        mv_0_n219) );
  OAI21_X1 mv_0_U328 ( .B1(ciphertext3[109]), .B2(ciphertext1[109]), .A(
        ciphertext2[109]), .ZN(mv_0_n220) );
  NAND2_X1 mv_0_U327 ( .A1(mv_0_n218), .A2(mv_0_n217), .ZN(ciphertext[108]) );
  NAND2_X1 mv_0_U326 ( .A1(ciphertext3[108]), .A2(ciphertext1[108]), .ZN(
        mv_0_n217) );
  OAI21_X1 mv_0_U325 ( .B1(ciphertext3[108]), .B2(ciphertext1[108]), .A(
        ciphertext2[108]), .ZN(mv_0_n218) );
  NAND2_X1 mv_0_U324 ( .A1(mv_0_n216), .A2(mv_0_n215), .ZN(ciphertext[107]) );
  NAND2_X1 mv_0_U323 ( .A1(ciphertext3[107]), .A2(ciphertext1[107]), .ZN(
        mv_0_n215) );
  OAI21_X1 mv_0_U322 ( .B1(ciphertext3[107]), .B2(ciphertext1[107]), .A(
        ciphertext2[107]), .ZN(mv_0_n216) );
  NAND2_X1 mv_0_U321 ( .A1(mv_0_n214), .A2(mv_0_n213), .ZN(ciphertext[106]) );
  NAND2_X1 mv_0_U320 ( .A1(ciphertext3[106]), .A2(ciphertext1[106]), .ZN(
        mv_0_n213) );
  OAI21_X1 mv_0_U319 ( .B1(ciphertext3[106]), .B2(ciphertext1[106]), .A(
        ciphertext2[106]), .ZN(mv_0_n214) );
  NAND2_X1 mv_0_U318 ( .A1(mv_0_n212), .A2(mv_0_n211), .ZN(ciphertext[105]) );
  NAND2_X1 mv_0_U317 ( .A1(ciphertext3[105]), .A2(ciphertext1[105]), .ZN(
        mv_0_n211) );
  OAI21_X1 mv_0_U316 ( .B1(ciphertext3[105]), .B2(ciphertext1[105]), .A(
        ciphertext2[105]), .ZN(mv_0_n212) );
  NAND2_X1 mv_0_U315 ( .A1(mv_0_n210), .A2(mv_0_n209), .ZN(ciphertext[104]) );
  NAND2_X1 mv_0_U314 ( .A1(ciphertext3[104]), .A2(ciphertext1[104]), .ZN(
        mv_0_n209) );
  OAI21_X1 mv_0_U313 ( .B1(ciphertext3[104]), .B2(ciphertext1[104]), .A(
        ciphertext2[104]), .ZN(mv_0_n210) );
  NAND2_X1 mv_0_U312 ( .A1(mv_0_n208), .A2(mv_0_n207), .ZN(ciphertext[103]) );
  NAND2_X1 mv_0_U311 ( .A1(ciphertext3[103]), .A2(ciphertext1[103]), .ZN(
        mv_0_n207) );
  OAI21_X1 mv_0_U310 ( .B1(ciphertext3[103]), .B2(ciphertext1[103]), .A(
        ciphertext2[103]), .ZN(mv_0_n208) );
  NAND2_X1 mv_0_U309 ( .A1(mv_0_n206), .A2(mv_0_n205), .ZN(ciphertext[102]) );
  NAND2_X1 mv_0_U308 ( .A1(ciphertext3[102]), .A2(ciphertext1[102]), .ZN(
        mv_0_n205) );
  OAI21_X1 mv_0_U307 ( .B1(ciphertext3[102]), .B2(ciphertext1[102]), .A(
        ciphertext2[102]), .ZN(mv_0_n206) );
  NAND2_X1 mv_0_U306 ( .A1(mv_0_n204), .A2(mv_0_n203), .ZN(ciphertext[101]) );
  NAND2_X1 mv_0_U305 ( .A1(ciphertext3[101]), .A2(ciphertext1[101]), .ZN(
        mv_0_n203) );
  OAI21_X1 mv_0_U304 ( .B1(ciphertext3[101]), .B2(ciphertext1[101]), .A(
        ciphertext2[101]), .ZN(mv_0_n204) );
  NAND2_X1 mv_0_U303 ( .A1(mv_0_n202), .A2(mv_0_n201), .ZN(ciphertext[100]) );
  NAND2_X1 mv_0_U302 ( .A1(ciphertext3[100]), .A2(ciphertext1[100]), .ZN(
        mv_0_n201) );
  OAI21_X1 mv_0_U301 ( .B1(ciphertext3[100]), .B2(ciphertext1[100]), .A(
        ciphertext2[100]), .ZN(mv_0_n202) );
  NAND2_X1 mv_0_U300 ( .A1(mv_0_n200), .A2(mv_0_n199), .ZN(ciphertext[99]) );
  NAND2_X1 mv_0_U299 ( .A1(ciphertext3[99]), .A2(ciphertext1[99]), .ZN(
        mv_0_n199) );
  OAI21_X1 mv_0_U298 ( .B1(ciphertext3[99]), .B2(ciphertext1[99]), .A(
        ciphertext2[99]), .ZN(mv_0_n200) );
  NAND2_X1 mv_0_U297 ( .A1(mv_0_n198), .A2(mv_0_n197), .ZN(ciphertext[98]) );
  NAND2_X1 mv_0_U296 ( .A1(ciphertext3[98]), .A2(ciphertext1[98]), .ZN(
        mv_0_n197) );
  OAI21_X1 mv_0_U295 ( .B1(ciphertext3[98]), .B2(ciphertext1[98]), .A(
        ciphertext2[98]), .ZN(mv_0_n198) );
  NAND2_X1 mv_0_U294 ( .A1(mv_0_n196), .A2(mv_0_n195), .ZN(ciphertext[97]) );
  NAND2_X1 mv_0_U293 ( .A1(ciphertext3[97]), .A2(ciphertext1[97]), .ZN(
        mv_0_n195) );
  OAI21_X1 mv_0_U292 ( .B1(ciphertext3[97]), .B2(ciphertext1[97]), .A(
        ciphertext2[97]), .ZN(mv_0_n196) );
  NAND2_X1 mv_0_U291 ( .A1(mv_0_n194), .A2(mv_0_n193), .ZN(ciphertext[96]) );
  NAND2_X1 mv_0_U290 ( .A1(ciphertext3[96]), .A2(ciphertext1[96]), .ZN(
        mv_0_n193) );
  OAI21_X1 mv_0_U289 ( .B1(ciphertext3[96]), .B2(ciphertext1[96]), .A(
        ciphertext2[96]), .ZN(mv_0_n194) );
  NAND2_X1 mv_0_U288 ( .A1(mv_0_n192), .A2(mv_0_n191), .ZN(ciphertext[95]) );
  NAND2_X1 mv_0_U287 ( .A1(ciphertext3[95]), .A2(ciphertext1[95]), .ZN(
        mv_0_n191) );
  OAI21_X1 mv_0_U286 ( .B1(ciphertext3[95]), .B2(ciphertext1[95]), .A(
        ciphertext2[95]), .ZN(mv_0_n192) );
  NAND2_X1 mv_0_U285 ( .A1(mv_0_n190), .A2(mv_0_n189), .ZN(ciphertext[94]) );
  NAND2_X1 mv_0_U284 ( .A1(ciphertext3[94]), .A2(ciphertext1[94]), .ZN(
        mv_0_n189) );
  OAI21_X1 mv_0_U283 ( .B1(ciphertext3[94]), .B2(ciphertext1[94]), .A(
        ciphertext2[94]), .ZN(mv_0_n190) );
  NAND2_X1 mv_0_U282 ( .A1(mv_0_n188), .A2(mv_0_n187), .ZN(ciphertext[93]) );
  NAND2_X1 mv_0_U281 ( .A1(ciphertext3[93]), .A2(ciphertext1[93]), .ZN(
        mv_0_n187) );
  OAI21_X1 mv_0_U280 ( .B1(ciphertext3[93]), .B2(ciphertext1[93]), .A(
        ciphertext2[93]), .ZN(mv_0_n188) );
  NAND2_X1 mv_0_U279 ( .A1(mv_0_n186), .A2(mv_0_n185), .ZN(ciphertext[92]) );
  NAND2_X1 mv_0_U278 ( .A1(ciphertext3[92]), .A2(ciphertext1[92]), .ZN(
        mv_0_n185) );
  OAI21_X1 mv_0_U277 ( .B1(ciphertext3[92]), .B2(ciphertext1[92]), .A(
        ciphertext2[92]), .ZN(mv_0_n186) );
  NAND2_X1 mv_0_U276 ( .A1(mv_0_n184), .A2(mv_0_n183), .ZN(ciphertext[91]) );
  NAND2_X1 mv_0_U275 ( .A1(ciphertext3[91]), .A2(ciphertext1[91]), .ZN(
        mv_0_n183) );
  OAI21_X1 mv_0_U274 ( .B1(ciphertext3[91]), .B2(ciphertext1[91]), .A(
        ciphertext2[91]), .ZN(mv_0_n184) );
  NAND2_X1 mv_0_U273 ( .A1(mv_0_n182), .A2(mv_0_n181), .ZN(ciphertext[90]) );
  NAND2_X1 mv_0_U272 ( .A1(ciphertext3[90]), .A2(ciphertext1[90]), .ZN(
        mv_0_n181) );
  OAI21_X1 mv_0_U271 ( .B1(ciphertext3[90]), .B2(ciphertext1[90]), .A(
        ciphertext2[90]), .ZN(mv_0_n182) );
  NAND2_X1 mv_0_U270 ( .A1(mv_0_n180), .A2(mv_0_n179), .ZN(ciphertext[89]) );
  NAND2_X1 mv_0_U269 ( .A1(ciphertext3[89]), .A2(ciphertext1[89]), .ZN(
        mv_0_n179) );
  OAI21_X1 mv_0_U268 ( .B1(ciphertext3[89]), .B2(ciphertext1[89]), .A(
        ciphertext2[89]), .ZN(mv_0_n180) );
  NAND2_X1 mv_0_U267 ( .A1(mv_0_n178), .A2(mv_0_n177), .ZN(ciphertext[88]) );
  NAND2_X1 mv_0_U266 ( .A1(ciphertext3[88]), .A2(ciphertext1[88]), .ZN(
        mv_0_n177) );
  OAI21_X1 mv_0_U265 ( .B1(ciphertext3[88]), .B2(ciphertext1[88]), .A(
        ciphertext2[88]), .ZN(mv_0_n178) );
  NAND2_X1 mv_0_U264 ( .A1(mv_0_n176), .A2(mv_0_n175), .ZN(ciphertext[87]) );
  NAND2_X1 mv_0_U263 ( .A1(ciphertext3[87]), .A2(ciphertext1[87]), .ZN(
        mv_0_n175) );
  OAI21_X1 mv_0_U262 ( .B1(ciphertext3[87]), .B2(ciphertext1[87]), .A(
        ciphertext2[87]), .ZN(mv_0_n176) );
  NAND2_X1 mv_0_U261 ( .A1(mv_0_n174), .A2(mv_0_n173), .ZN(ciphertext[86]) );
  NAND2_X1 mv_0_U260 ( .A1(ciphertext3[86]), .A2(ciphertext1[86]), .ZN(
        mv_0_n173) );
  OAI21_X1 mv_0_U259 ( .B1(ciphertext3[86]), .B2(ciphertext1[86]), .A(
        ciphertext2[86]), .ZN(mv_0_n174) );
  NAND2_X1 mv_0_U258 ( .A1(mv_0_n172), .A2(mv_0_n171), .ZN(ciphertext[85]) );
  NAND2_X1 mv_0_U257 ( .A1(ciphertext3[85]), .A2(ciphertext1[85]), .ZN(
        mv_0_n171) );
  OAI21_X1 mv_0_U256 ( .B1(ciphertext3[85]), .B2(ciphertext1[85]), .A(
        ciphertext2[85]), .ZN(mv_0_n172) );
  NAND2_X1 mv_0_U255 ( .A1(mv_0_n170), .A2(mv_0_n169), .ZN(ciphertext[84]) );
  NAND2_X1 mv_0_U254 ( .A1(ciphertext3[84]), .A2(ciphertext1[84]), .ZN(
        mv_0_n169) );
  OAI21_X1 mv_0_U253 ( .B1(ciphertext3[84]), .B2(ciphertext1[84]), .A(
        ciphertext2[84]), .ZN(mv_0_n170) );
  NAND2_X1 mv_0_U252 ( .A1(mv_0_n168), .A2(mv_0_n167), .ZN(ciphertext[83]) );
  NAND2_X1 mv_0_U251 ( .A1(ciphertext3[83]), .A2(ciphertext1[83]), .ZN(
        mv_0_n167) );
  OAI21_X1 mv_0_U250 ( .B1(ciphertext3[83]), .B2(ciphertext1[83]), .A(
        ciphertext2[83]), .ZN(mv_0_n168) );
  NAND2_X1 mv_0_U249 ( .A1(mv_0_n166), .A2(mv_0_n165), .ZN(ciphertext[82]) );
  NAND2_X1 mv_0_U248 ( .A1(ciphertext3[82]), .A2(ciphertext1[82]), .ZN(
        mv_0_n165) );
  OAI21_X1 mv_0_U247 ( .B1(ciphertext3[82]), .B2(ciphertext1[82]), .A(
        ciphertext2[82]), .ZN(mv_0_n166) );
  NAND2_X1 mv_0_U246 ( .A1(mv_0_n164), .A2(mv_0_n163), .ZN(ciphertext[81]) );
  NAND2_X1 mv_0_U245 ( .A1(ciphertext3[81]), .A2(ciphertext1[81]), .ZN(
        mv_0_n163) );
  OAI21_X1 mv_0_U244 ( .B1(ciphertext3[81]), .B2(ciphertext1[81]), .A(
        ciphertext2[81]), .ZN(mv_0_n164) );
  NAND2_X1 mv_0_U243 ( .A1(mv_0_n162), .A2(mv_0_n161), .ZN(ciphertext[80]) );
  NAND2_X1 mv_0_U242 ( .A1(ciphertext3[80]), .A2(ciphertext1[80]), .ZN(
        mv_0_n161) );
  OAI21_X1 mv_0_U241 ( .B1(ciphertext3[80]), .B2(ciphertext1[80]), .A(
        ciphertext2[80]), .ZN(mv_0_n162) );
  NAND2_X1 mv_0_U240 ( .A1(mv_0_n160), .A2(mv_0_n159), .ZN(ciphertext[79]) );
  NAND2_X1 mv_0_U239 ( .A1(ciphertext3[79]), .A2(ciphertext1[79]), .ZN(
        mv_0_n159) );
  OAI21_X1 mv_0_U238 ( .B1(ciphertext3[79]), .B2(ciphertext1[79]), .A(
        ciphertext2[79]), .ZN(mv_0_n160) );
  NAND2_X1 mv_0_U237 ( .A1(mv_0_n158), .A2(mv_0_n157), .ZN(ciphertext[78]) );
  NAND2_X1 mv_0_U236 ( .A1(ciphertext3[78]), .A2(ciphertext1[78]), .ZN(
        mv_0_n157) );
  OAI21_X1 mv_0_U235 ( .B1(ciphertext3[78]), .B2(ciphertext1[78]), .A(
        ciphertext2[78]), .ZN(mv_0_n158) );
  NAND2_X1 mv_0_U234 ( .A1(mv_0_n156), .A2(mv_0_n155), .ZN(ciphertext[77]) );
  NAND2_X1 mv_0_U233 ( .A1(ciphertext3[77]), .A2(ciphertext1[77]), .ZN(
        mv_0_n155) );
  OAI21_X1 mv_0_U232 ( .B1(ciphertext3[77]), .B2(ciphertext1[77]), .A(
        ciphertext2[77]), .ZN(mv_0_n156) );
  NAND2_X1 mv_0_U231 ( .A1(mv_0_n154), .A2(mv_0_n153), .ZN(ciphertext[76]) );
  NAND2_X1 mv_0_U230 ( .A1(ciphertext3[76]), .A2(ciphertext1[76]), .ZN(
        mv_0_n153) );
  OAI21_X1 mv_0_U229 ( .B1(ciphertext3[76]), .B2(ciphertext1[76]), .A(
        ciphertext2[76]), .ZN(mv_0_n154) );
  NAND2_X1 mv_0_U228 ( .A1(mv_0_n152), .A2(mv_0_n151), .ZN(ciphertext[75]) );
  NAND2_X1 mv_0_U227 ( .A1(ciphertext3[75]), .A2(ciphertext1[75]), .ZN(
        mv_0_n151) );
  OAI21_X1 mv_0_U226 ( .B1(ciphertext3[75]), .B2(ciphertext1[75]), .A(
        ciphertext2[75]), .ZN(mv_0_n152) );
  NAND2_X1 mv_0_U225 ( .A1(mv_0_n150), .A2(mv_0_n149), .ZN(ciphertext[74]) );
  NAND2_X1 mv_0_U224 ( .A1(ciphertext3[74]), .A2(ciphertext1[74]), .ZN(
        mv_0_n149) );
  OAI21_X1 mv_0_U223 ( .B1(ciphertext3[74]), .B2(ciphertext1[74]), .A(
        ciphertext2[74]), .ZN(mv_0_n150) );
  NAND2_X1 mv_0_U222 ( .A1(mv_0_n148), .A2(mv_0_n147), .ZN(ciphertext[73]) );
  NAND2_X1 mv_0_U221 ( .A1(ciphertext3[73]), .A2(ciphertext1[73]), .ZN(
        mv_0_n147) );
  OAI21_X1 mv_0_U220 ( .B1(ciphertext3[73]), .B2(ciphertext1[73]), .A(
        ciphertext2[73]), .ZN(mv_0_n148) );
  NAND2_X1 mv_0_U219 ( .A1(mv_0_n146), .A2(mv_0_n145), .ZN(ciphertext[72]) );
  NAND2_X1 mv_0_U218 ( .A1(ciphertext3[72]), .A2(ciphertext1[72]), .ZN(
        mv_0_n145) );
  OAI21_X1 mv_0_U217 ( .B1(ciphertext3[72]), .B2(ciphertext1[72]), .A(
        ciphertext2[72]), .ZN(mv_0_n146) );
  NAND2_X1 mv_0_U216 ( .A1(mv_0_n144), .A2(mv_0_n143), .ZN(ciphertext[71]) );
  NAND2_X1 mv_0_U215 ( .A1(ciphertext3[71]), .A2(ciphertext1[71]), .ZN(
        mv_0_n143) );
  OAI21_X1 mv_0_U214 ( .B1(ciphertext3[71]), .B2(ciphertext1[71]), .A(
        ciphertext2[71]), .ZN(mv_0_n144) );
  NAND2_X1 mv_0_U213 ( .A1(mv_0_n142), .A2(mv_0_n141), .ZN(ciphertext[70]) );
  NAND2_X1 mv_0_U212 ( .A1(ciphertext3[70]), .A2(ciphertext1[70]), .ZN(
        mv_0_n141) );
  OAI21_X1 mv_0_U211 ( .B1(ciphertext3[70]), .B2(ciphertext1[70]), .A(
        ciphertext2[70]), .ZN(mv_0_n142) );
  NAND2_X1 mv_0_U210 ( .A1(mv_0_n140), .A2(mv_0_n139), .ZN(ciphertext[69]) );
  NAND2_X1 mv_0_U209 ( .A1(ciphertext3[69]), .A2(ciphertext1[69]), .ZN(
        mv_0_n139) );
  OAI21_X1 mv_0_U208 ( .B1(ciphertext3[69]), .B2(ciphertext1[69]), .A(
        ciphertext2[69]), .ZN(mv_0_n140) );
  NAND2_X1 mv_0_U207 ( .A1(mv_0_n138), .A2(mv_0_n137), .ZN(ciphertext[68]) );
  NAND2_X1 mv_0_U206 ( .A1(ciphertext3[68]), .A2(ciphertext1[68]), .ZN(
        mv_0_n137) );
  OAI21_X1 mv_0_U205 ( .B1(ciphertext3[68]), .B2(ciphertext1[68]), .A(
        ciphertext2[68]), .ZN(mv_0_n138) );
  NAND2_X1 mv_0_U204 ( .A1(mv_0_n136), .A2(mv_0_n135), .ZN(ciphertext[67]) );
  NAND2_X1 mv_0_U203 ( .A1(ciphertext3[67]), .A2(ciphertext1[67]), .ZN(
        mv_0_n135) );
  OAI21_X1 mv_0_U202 ( .B1(ciphertext3[67]), .B2(ciphertext1[67]), .A(
        ciphertext2[67]), .ZN(mv_0_n136) );
  NAND2_X1 mv_0_U201 ( .A1(mv_0_n134), .A2(mv_0_n133), .ZN(ciphertext[66]) );
  NAND2_X1 mv_0_U200 ( .A1(ciphertext3[66]), .A2(ciphertext1[66]), .ZN(
        mv_0_n133) );
  OAI21_X1 mv_0_U199 ( .B1(ciphertext3[66]), .B2(ciphertext1[66]), .A(
        ciphertext2[66]), .ZN(mv_0_n134) );
  NAND2_X1 mv_0_U198 ( .A1(mv_0_n132), .A2(mv_0_n131), .ZN(ciphertext[65]) );
  NAND2_X1 mv_0_U197 ( .A1(ciphertext3[65]), .A2(ciphertext1[65]), .ZN(
        mv_0_n131) );
  OAI21_X1 mv_0_U196 ( .B1(ciphertext3[65]), .B2(ciphertext1[65]), .A(
        ciphertext2[65]), .ZN(mv_0_n132) );
  NAND2_X1 mv_0_U195 ( .A1(mv_0_n130), .A2(mv_0_n129), .ZN(ciphertext[64]) );
  NAND2_X1 mv_0_U194 ( .A1(ciphertext3[64]), .A2(ciphertext1[64]), .ZN(
        mv_0_n129) );
  OAI21_X1 mv_0_U193 ( .B1(ciphertext3[64]), .B2(ciphertext1[64]), .A(
        ciphertext2[64]), .ZN(mv_0_n130) );
  NAND2_X1 mv_0_U192 ( .A1(mv_0_n128), .A2(mv_0_n127), .ZN(ciphertext[63]) );
  NAND2_X1 mv_0_U191 ( .A1(ciphertext3[63]), .A2(ciphertext1[63]), .ZN(
        mv_0_n127) );
  OAI21_X1 mv_0_U190 ( .B1(ciphertext3[63]), .B2(ciphertext1[63]), .A(
        ciphertext2[63]), .ZN(mv_0_n128) );
  NAND2_X1 mv_0_U189 ( .A1(mv_0_n126), .A2(mv_0_n125), .ZN(ciphertext[62]) );
  NAND2_X1 mv_0_U188 ( .A1(ciphertext3[62]), .A2(ciphertext1[62]), .ZN(
        mv_0_n125) );
  OAI21_X1 mv_0_U187 ( .B1(ciphertext3[62]), .B2(ciphertext1[62]), .A(
        ciphertext2[62]), .ZN(mv_0_n126) );
  NAND2_X1 mv_0_U186 ( .A1(mv_0_n124), .A2(mv_0_n123), .ZN(ciphertext[61]) );
  NAND2_X1 mv_0_U185 ( .A1(ciphertext3[61]), .A2(ciphertext1[61]), .ZN(
        mv_0_n123) );
  OAI21_X1 mv_0_U184 ( .B1(ciphertext3[61]), .B2(ciphertext1[61]), .A(
        ciphertext2[61]), .ZN(mv_0_n124) );
  NAND2_X1 mv_0_U183 ( .A1(mv_0_n122), .A2(mv_0_n121), .ZN(ciphertext[60]) );
  NAND2_X1 mv_0_U182 ( .A1(ciphertext3[60]), .A2(ciphertext1[60]), .ZN(
        mv_0_n121) );
  OAI21_X1 mv_0_U181 ( .B1(ciphertext3[60]), .B2(ciphertext1[60]), .A(
        ciphertext2[60]), .ZN(mv_0_n122) );
  NAND2_X1 mv_0_U180 ( .A1(mv_0_n120), .A2(mv_0_n119), .ZN(ciphertext[59]) );
  NAND2_X1 mv_0_U179 ( .A1(ciphertext3[59]), .A2(ciphertext1[59]), .ZN(
        mv_0_n119) );
  OAI21_X1 mv_0_U178 ( .B1(ciphertext3[59]), .B2(ciphertext1[59]), .A(
        ciphertext2[59]), .ZN(mv_0_n120) );
  NAND2_X1 mv_0_U177 ( .A1(mv_0_n118), .A2(mv_0_n117), .ZN(ciphertext[58]) );
  NAND2_X1 mv_0_U176 ( .A1(ciphertext3[58]), .A2(ciphertext1[58]), .ZN(
        mv_0_n117) );
  OAI21_X1 mv_0_U175 ( .B1(ciphertext3[58]), .B2(ciphertext1[58]), .A(
        ciphertext2[58]), .ZN(mv_0_n118) );
  NAND2_X1 mv_0_U174 ( .A1(mv_0_n116), .A2(mv_0_n115), .ZN(ciphertext[57]) );
  NAND2_X1 mv_0_U173 ( .A1(ciphertext3[57]), .A2(ciphertext1[57]), .ZN(
        mv_0_n115) );
  OAI21_X1 mv_0_U172 ( .B1(ciphertext3[57]), .B2(ciphertext1[57]), .A(
        ciphertext2[57]), .ZN(mv_0_n116) );
  NAND2_X1 mv_0_U171 ( .A1(mv_0_n114), .A2(mv_0_n113), .ZN(ciphertext[56]) );
  NAND2_X1 mv_0_U170 ( .A1(ciphertext3[56]), .A2(ciphertext1[56]), .ZN(
        mv_0_n113) );
  OAI21_X1 mv_0_U169 ( .B1(ciphertext3[56]), .B2(ciphertext1[56]), .A(
        ciphertext2[56]), .ZN(mv_0_n114) );
  NAND2_X1 mv_0_U168 ( .A1(mv_0_n112), .A2(mv_0_n111), .ZN(ciphertext[55]) );
  NAND2_X1 mv_0_U167 ( .A1(ciphertext3[55]), .A2(ciphertext1[55]), .ZN(
        mv_0_n111) );
  OAI21_X1 mv_0_U166 ( .B1(ciphertext3[55]), .B2(ciphertext1[55]), .A(
        ciphertext2[55]), .ZN(mv_0_n112) );
  NAND2_X1 mv_0_U165 ( .A1(mv_0_n110), .A2(mv_0_n109), .ZN(ciphertext[54]) );
  NAND2_X1 mv_0_U164 ( .A1(ciphertext3[54]), .A2(ciphertext1[54]), .ZN(
        mv_0_n109) );
  OAI21_X1 mv_0_U163 ( .B1(ciphertext3[54]), .B2(ciphertext1[54]), .A(
        ciphertext2[54]), .ZN(mv_0_n110) );
  NAND2_X1 mv_0_U162 ( .A1(mv_0_n108), .A2(mv_0_n107), .ZN(ciphertext[53]) );
  NAND2_X1 mv_0_U161 ( .A1(ciphertext3[53]), .A2(ciphertext1[53]), .ZN(
        mv_0_n107) );
  OAI21_X1 mv_0_U160 ( .B1(ciphertext3[53]), .B2(ciphertext1[53]), .A(
        ciphertext2[53]), .ZN(mv_0_n108) );
  NAND2_X1 mv_0_U159 ( .A1(mv_0_n106), .A2(mv_0_n105), .ZN(ciphertext[52]) );
  NAND2_X1 mv_0_U158 ( .A1(ciphertext3[52]), .A2(ciphertext1[52]), .ZN(
        mv_0_n105) );
  OAI21_X1 mv_0_U157 ( .B1(ciphertext3[52]), .B2(ciphertext1[52]), .A(
        ciphertext2[52]), .ZN(mv_0_n106) );
  NAND2_X1 mv_0_U156 ( .A1(mv_0_n104), .A2(mv_0_n103), .ZN(ciphertext[51]) );
  NAND2_X1 mv_0_U155 ( .A1(ciphertext3[51]), .A2(ciphertext1[51]), .ZN(
        mv_0_n103) );
  OAI21_X1 mv_0_U154 ( .B1(ciphertext3[51]), .B2(ciphertext1[51]), .A(
        ciphertext2[51]), .ZN(mv_0_n104) );
  NAND2_X1 mv_0_U153 ( .A1(mv_0_n102), .A2(mv_0_n101), .ZN(ciphertext[50]) );
  NAND2_X1 mv_0_U152 ( .A1(ciphertext3[50]), .A2(ciphertext1[50]), .ZN(
        mv_0_n101) );
  OAI21_X1 mv_0_U151 ( .B1(ciphertext3[50]), .B2(ciphertext1[50]), .A(
        ciphertext2[50]), .ZN(mv_0_n102) );
  NAND2_X1 mv_0_U150 ( .A1(mv_0_n100), .A2(mv_0_n99), .ZN(ciphertext[49]) );
  NAND2_X1 mv_0_U149 ( .A1(ciphertext3[49]), .A2(ciphertext1[49]), .ZN(
        mv_0_n99) );
  OAI21_X1 mv_0_U148 ( .B1(ciphertext3[49]), .B2(ciphertext1[49]), .A(
        ciphertext2[49]), .ZN(mv_0_n100) );
  NAND2_X1 mv_0_U147 ( .A1(mv_0_n98), .A2(mv_0_n97), .ZN(ciphertext[48]) );
  NAND2_X1 mv_0_U146 ( .A1(ciphertext3[48]), .A2(ciphertext1[48]), .ZN(
        mv_0_n97) );
  OAI21_X1 mv_0_U145 ( .B1(ciphertext3[48]), .B2(ciphertext1[48]), .A(
        ciphertext2[48]), .ZN(mv_0_n98) );
  NAND2_X1 mv_0_U144 ( .A1(mv_0_n96), .A2(mv_0_n95), .ZN(ciphertext[47]) );
  NAND2_X1 mv_0_U143 ( .A1(ciphertext3[47]), .A2(ciphertext1[47]), .ZN(
        mv_0_n95) );
  OAI21_X1 mv_0_U142 ( .B1(ciphertext3[47]), .B2(ciphertext1[47]), .A(
        ciphertext2[47]), .ZN(mv_0_n96) );
  NAND2_X1 mv_0_U141 ( .A1(mv_0_n94), .A2(mv_0_n93), .ZN(ciphertext[46]) );
  NAND2_X1 mv_0_U140 ( .A1(ciphertext3[46]), .A2(ciphertext1[46]), .ZN(
        mv_0_n93) );
  OAI21_X1 mv_0_U139 ( .B1(ciphertext3[46]), .B2(ciphertext1[46]), .A(
        ciphertext2[46]), .ZN(mv_0_n94) );
  NAND2_X1 mv_0_U138 ( .A1(mv_0_n92), .A2(mv_0_n91), .ZN(ciphertext[45]) );
  NAND2_X1 mv_0_U137 ( .A1(ciphertext3[45]), .A2(ciphertext1[45]), .ZN(
        mv_0_n91) );
  OAI21_X1 mv_0_U136 ( .B1(ciphertext3[45]), .B2(ciphertext1[45]), .A(
        ciphertext2[45]), .ZN(mv_0_n92) );
  NAND2_X1 mv_0_U135 ( .A1(mv_0_n90), .A2(mv_0_n89), .ZN(ciphertext[44]) );
  NAND2_X1 mv_0_U134 ( .A1(ciphertext3[44]), .A2(ciphertext1[44]), .ZN(
        mv_0_n89) );
  OAI21_X1 mv_0_U133 ( .B1(ciphertext3[44]), .B2(ciphertext1[44]), .A(
        ciphertext2[44]), .ZN(mv_0_n90) );
  NAND2_X1 mv_0_U132 ( .A1(mv_0_n88), .A2(mv_0_n87), .ZN(ciphertext[43]) );
  NAND2_X1 mv_0_U131 ( .A1(ciphertext3[43]), .A2(ciphertext1[43]), .ZN(
        mv_0_n87) );
  OAI21_X1 mv_0_U130 ( .B1(ciphertext3[43]), .B2(ciphertext1[43]), .A(
        ciphertext2[43]), .ZN(mv_0_n88) );
  NAND2_X1 mv_0_U129 ( .A1(mv_0_n86), .A2(mv_0_n85), .ZN(ciphertext[42]) );
  NAND2_X1 mv_0_U128 ( .A1(ciphertext3[42]), .A2(ciphertext1[42]), .ZN(
        mv_0_n85) );
  OAI21_X1 mv_0_U127 ( .B1(ciphertext3[42]), .B2(ciphertext1[42]), .A(
        ciphertext2[42]), .ZN(mv_0_n86) );
  NAND2_X1 mv_0_U126 ( .A1(mv_0_n84), .A2(mv_0_n83), .ZN(ciphertext[41]) );
  NAND2_X1 mv_0_U125 ( .A1(ciphertext3[41]), .A2(ciphertext1[41]), .ZN(
        mv_0_n83) );
  OAI21_X1 mv_0_U124 ( .B1(ciphertext3[41]), .B2(ciphertext1[41]), .A(
        ciphertext2[41]), .ZN(mv_0_n84) );
  NAND2_X1 mv_0_U123 ( .A1(mv_0_n82), .A2(mv_0_n81), .ZN(ciphertext[40]) );
  NAND2_X1 mv_0_U122 ( .A1(ciphertext3[40]), .A2(ciphertext1[40]), .ZN(
        mv_0_n81) );
  OAI21_X1 mv_0_U121 ( .B1(ciphertext3[40]), .B2(ciphertext1[40]), .A(
        ciphertext2[40]), .ZN(mv_0_n82) );
  NAND2_X1 mv_0_U120 ( .A1(mv_0_n80), .A2(mv_0_n79), .ZN(ciphertext[39]) );
  NAND2_X1 mv_0_U119 ( .A1(ciphertext3[39]), .A2(ciphertext1[39]), .ZN(
        mv_0_n79) );
  OAI21_X1 mv_0_U118 ( .B1(ciphertext3[39]), .B2(ciphertext1[39]), .A(
        ciphertext2[39]), .ZN(mv_0_n80) );
  NAND2_X1 mv_0_U117 ( .A1(mv_0_n78), .A2(mv_0_n77), .ZN(ciphertext[38]) );
  NAND2_X1 mv_0_U116 ( .A1(ciphertext3[38]), .A2(ciphertext1[38]), .ZN(
        mv_0_n77) );
  OAI21_X1 mv_0_U115 ( .B1(ciphertext3[38]), .B2(ciphertext1[38]), .A(
        ciphertext2[38]), .ZN(mv_0_n78) );
  NAND2_X1 mv_0_U114 ( .A1(mv_0_n76), .A2(mv_0_n75), .ZN(ciphertext[37]) );
  NAND2_X1 mv_0_U113 ( .A1(ciphertext3[37]), .A2(ciphertext1[37]), .ZN(
        mv_0_n75) );
  OAI21_X1 mv_0_U112 ( .B1(ciphertext3[37]), .B2(ciphertext1[37]), .A(
        ciphertext2[37]), .ZN(mv_0_n76) );
  NAND2_X1 mv_0_U111 ( .A1(mv_0_n74), .A2(mv_0_n73), .ZN(ciphertext[36]) );
  NAND2_X1 mv_0_U110 ( .A1(ciphertext3[36]), .A2(ciphertext1[36]), .ZN(
        mv_0_n73) );
  OAI21_X1 mv_0_U109 ( .B1(ciphertext3[36]), .B2(ciphertext1[36]), .A(
        ciphertext2[36]), .ZN(mv_0_n74) );
  NAND2_X1 mv_0_U108 ( .A1(mv_0_n72), .A2(mv_0_n71), .ZN(ciphertext[35]) );
  NAND2_X1 mv_0_U107 ( .A1(ciphertext3[35]), .A2(ciphertext1[35]), .ZN(
        mv_0_n71) );
  OAI21_X1 mv_0_U106 ( .B1(ciphertext3[35]), .B2(ciphertext1[35]), .A(
        ciphertext2[35]), .ZN(mv_0_n72) );
  NAND2_X1 mv_0_U105 ( .A1(mv_0_n70), .A2(mv_0_n69), .ZN(ciphertext[34]) );
  NAND2_X1 mv_0_U104 ( .A1(ciphertext3[34]), .A2(ciphertext1[34]), .ZN(
        mv_0_n69) );
  OAI21_X1 mv_0_U103 ( .B1(ciphertext3[34]), .B2(ciphertext1[34]), .A(
        ciphertext2[34]), .ZN(mv_0_n70) );
  NAND2_X1 mv_0_U102 ( .A1(mv_0_n68), .A2(mv_0_n67), .ZN(ciphertext[33]) );
  NAND2_X1 mv_0_U101 ( .A1(ciphertext3[33]), .A2(ciphertext1[33]), .ZN(
        mv_0_n67) );
  OAI21_X1 mv_0_U100 ( .B1(ciphertext3[33]), .B2(ciphertext1[33]), .A(
        ciphertext2[33]), .ZN(mv_0_n68) );
  NAND2_X1 mv_0_U99 ( .A1(mv_0_n66), .A2(mv_0_n65), .ZN(ciphertext[32]) );
  NAND2_X1 mv_0_U98 ( .A1(ciphertext3[32]), .A2(ciphertext1[32]), .ZN(mv_0_n65) );
  OAI21_X1 mv_0_U97 ( .B1(ciphertext3[32]), .B2(ciphertext1[32]), .A(
        ciphertext2[32]), .ZN(mv_0_n66) );
  NAND2_X1 mv_0_U96 ( .A1(mv_0_n64), .A2(mv_0_n63), .ZN(ciphertext[31]) );
  NAND2_X1 mv_0_U95 ( .A1(ciphertext3[31]), .A2(ciphertext1[31]), .ZN(mv_0_n63) );
  OAI21_X1 mv_0_U94 ( .B1(ciphertext3[31]), .B2(ciphertext1[31]), .A(
        ciphertext2[31]), .ZN(mv_0_n64) );
  NAND2_X1 mv_0_U93 ( .A1(mv_0_n62), .A2(mv_0_n61), .ZN(ciphertext[30]) );
  NAND2_X1 mv_0_U92 ( .A1(ciphertext3[30]), .A2(ciphertext1[30]), .ZN(mv_0_n61) );
  OAI21_X1 mv_0_U91 ( .B1(ciphertext3[30]), .B2(ciphertext1[30]), .A(
        ciphertext2[30]), .ZN(mv_0_n62) );
  NAND2_X1 mv_0_U90 ( .A1(mv_0_n60), .A2(mv_0_n59), .ZN(ciphertext[29]) );
  NAND2_X1 mv_0_U89 ( .A1(ciphertext3[29]), .A2(ciphertext1[29]), .ZN(mv_0_n59) );
  OAI21_X1 mv_0_U88 ( .B1(ciphertext3[29]), .B2(ciphertext1[29]), .A(
        ciphertext2[29]), .ZN(mv_0_n60) );
  NAND2_X1 mv_0_U87 ( .A1(mv_0_n58), .A2(mv_0_n57), .ZN(ciphertext[28]) );
  NAND2_X1 mv_0_U86 ( .A1(ciphertext3[28]), .A2(ciphertext1[28]), .ZN(mv_0_n57) );
  OAI21_X1 mv_0_U85 ( .B1(ciphertext3[28]), .B2(ciphertext1[28]), .A(
        ciphertext2[28]), .ZN(mv_0_n58) );
  NAND2_X1 mv_0_U84 ( .A1(mv_0_n56), .A2(mv_0_n55), .ZN(ciphertext[27]) );
  NAND2_X1 mv_0_U83 ( .A1(ciphertext3[27]), .A2(ciphertext1[27]), .ZN(mv_0_n55) );
  OAI21_X1 mv_0_U82 ( .B1(ciphertext3[27]), .B2(ciphertext1[27]), .A(
        ciphertext2[27]), .ZN(mv_0_n56) );
  NAND2_X1 mv_0_U81 ( .A1(mv_0_n54), .A2(mv_0_n53), .ZN(ciphertext[26]) );
  NAND2_X1 mv_0_U80 ( .A1(ciphertext3[26]), .A2(ciphertext1[26]), .ZN(mv_0_n53) );
  OAI21_X1 mv_0_U79 ( .B1(ciphertext3[26]), .B2(ciphertext1[26]), .A(
        ciphertext2[26]), .ZN(mv_0_n54) );
  NAND2_X1 mv_0_U78 ( .A1(mv_0_n52), .A2(mv_0_n51), .ZN(ciphertext[25]) );
  NAND2_X1 mv_0_U77 ( .A1(ciphertext3[25]), .A2(ciphertext1[25]), .ZN(mv_0_n51) );
  OAI21_X1 mv_0_U76 ( .B1(ciphertext3[25]), .B2(ciphertext1[25]), .A(
        ciphertext2[25]), .ZN(mv_0_n52) );
  NAND2_X1 mv_0_U75 ( .A1(mv_0_n50), .A2(mv_0_n49), .ZN(ciphertext[24]) );
  NAND2_X1 mv_0_U74 ( .A1(ciphertext3[24]), .A2(ciphertext1[24]), .ZN(mv_0_n49) );
  OAI21_X1 mv_0_U73 ( .B1(ciphertext3[24]), .B2(ciphertext1[24]), .A(
        ciphertext2[24]), .ZN(mv_0_n50) );
  NAND2_X1 mv_0_U72 ( .A1(mv_0_n48), .A2(mv_0_n47), .ZN(ciphertext[23]) );
  NAND2_X1 mv_0_U71 ( .A1(ciphertext3[23]), .A2(ciphertext1[23]), .ZN(mv_0_n47) );
  OAI21_X1 mv_0_U70 ( .B1(ciphertext3[23]), .B2(ciphertext1[23]), .A(
        ciphertext2[23]), .ZN(mv_0_n48) );
  NAND2_X1 mv_0_U69 ( .A1(mv_0_n46), .A2(mv_0_n45), .ZN(ciphertext[22]) );
  NAND2_X1 mv_0_U68 ( .A1(ciphertext3[22]), .A2(ciphertext1[22]), .ZN(mv_0_n45) );
  OAI21_X1 mv_0_U67 ( .B1(ciphertext3[22]), .B2(ciphertext1[22]), .A(
        ciphertext2[22]), .ZN(mv_0_n46) );
  NAND2_X1 mv_0_U66 ( .A1(mv_0_n44), .A2(mv_0_n43), .ZN(ciphertext[21]) );
  NAND2_X1 mv_0_U65 ( .A1(ciphertext3[21]), .A2(ciphertext1[21]), .ZN(mv_0_n43) );
  OAI21_X1 mv_0_U64 ( .B1(ciphertext3[21]), .B2(ciphertext1[21]), .A(
        ciphertext2[21]), .ZN(mv_0_n44) );
  NAND2_X1 mv_0_U63 ( .A1(mv_0_n42), .A2(mv_0_n41), .ZN(ciphertext[20]) );
  NAND2_X1 mv_0_U62 ( .A1(ciphertext3[20]), .A2(ciphertext1[20]), .ZN(mv_0_n41) );
  OAI21_X1 mv_0_U61 ( .B1(ciphertext3[20]), .B2(ciphertext1[20]), .A(
        ciphertext2[20]), .ZN(mv_0_n42) );
  NAND2_X1 mv_0_U60 ( .A1(mv_0_n40), .A2(mv_0_n39), .ZN(ciphertext[19]) );
  NAND2_X1 mv_0_U59 ( .A1(ciphertext3[19]), .A2(ciphertext1[19]), .ZN(mv_0_n39) );
  OAI21_X1 mv_0_U58 ( .B1(ciphertext3[19]), .B2(ciphertext1[19]), .A(
        ciphertext2[19]), .ZN(mv_0_n40) );
  NAND2_X1 mv_0_U57 ( .A1(mv_0_n38), .A2(mv_0_n37), .ZN(ciphertext[18]) );
  NAND2_X1 mv_0_U56 ( .A1(ciphertext3[18]), .A2(ciphertext1[18]), .ZN(mv_0_n37) );
  OAI21_X1 mv_0_U55 ( .B1(ciphertext3[18]), .B2(ciphertext1[18]), .A(
        ciphertext2[18]), .ZN(mv_0_n38) );
  NAND2_X1 mv_0_U54 ( .A1(mv_0_n36), .A2(mv_0_n35), .ZN(ciphertext[17]) );
  NAND2_X1 mv_0_U53 ( .A1(ciphertext3[17]), .A2(ciphertext1[17]), .ZN(mv_0_n35) );
  OAI21_X1 mv_0_U52 ( .B1(ciphertext3[17]), .B2(ciphertext1[17]), .A(
        ciphertext2[17]), .ZN(mv_0_n36) );
  NAND2_X1 mv_0_U51 ( .A1(mv_0_n34), .A2(mv_0_n33), .ZN(ciphertext[16]) );
  NAND2_X1 mv_0_U50 ( .A1(ciphertext3[16]), .A2(ciphertext1[16]), .ZN(mv_0_n33) );
  OAI21_X1 mv_0_U49 ( .B1(ciphertext3[16]), .B2(ciphertext1[16]), .A(
        ciphertext2[16]), .ZN(mv_0_n34) );
  NAND2_X1 mv_0_U48 ( .A1(mv_0_n32), .A2(mv_0_n31), .ZN(ciphertext[15]) );
  NAND2_X1 mv_0_U47 ( .A1(ciphertext3[15]), .A2(ciphertext1[15]), .ZN(mv_0_n31) );
  OAI21_X1 mv_0_U46 ( .B1(ciphertext3[15]), .B2(ciphertext1[15]), .A(
        ciphertext2[15]), .ZN(mv_0_n32) );
  NAND2_X1 mv_0_U45 ( .A1(mv_0_n30), .A2(mv_0_n29), .ZN(ciphertext[14]) );
  NAND2_X1 mv_0_U44 ( .A1(ciphertext3[14]), .A2(ciphertext1[14]), .ZN(mv_0_n29) );
  OAI21_X1 mv_0_U43 ( .B1(ciphertext3[14]), .B2(ciphertext1[14]), .A(
        ciphertext2[14]), .ZN(mv_0_n30) );
  NAND2_X1 mv_0_U42 ( .A1(mv_0_n28), .A2(mv_0_n27), .ZN(ciphertext[13]) );
  NAND2_X1 mv_0_U41 ( .A1(ciphertext3[13]), .A2(ciphertext1[13]), .ZN(mv_0_n27) );
  OAI21_X1 mv_0_U40 ( .B1(ciphertext3[13]), .B2(ciphertext1[13]), .A(
        ciphertext2[13]), .ZN(mv_0_n28) );
  NAND2_X1 mv_0_U39 ( .A1(mv_0_n26), .A2(mv_0_n25), .ZN(ciphertext[12]) );
  NAND2_X1 mv_0_U38 ( .A1(ciphertext3[12]), .A2(ciphertext1[12]), .ZN(mv_0_n25) );
  OAI21_X1 mv_0_U37 ( .B1(ciphertext3[12]), .B2(ciphertext1[12]), .A(
        ciphertext2[12]), .ZN(mv_0_n26) );
  NAND2_X1 mv_0_U36 ( .A1(mv_0_n24), .A2(mv_0_n23), .ZN(ciphertext[11]) );
  NAND2_X1 mv_0_U35 ( .A1(ciphertext3[11]), .A2(ciphertext1[11]), .ZN(mv_0_n23) );
  OAI21_X1 mv_0_U34 ( .B1(ciphertext3[11]), .B2(ciphertext1[11]), .A(
        ciphertext2[11]), .ZN(mv_0_n24) );
  NAND2_X1 mv_0_U33 ( .A1(mv_0_n22), .A2(mv_0_n21), .ZN(ciphertext[10]) );
  NAND2_X1 mv_0_U32 ( .A1(ciphertext3[10]), .A2(ciphertext1[10]), .ZN(mv_0_n21) );
  OAI21_X1 mv_0_U31 ( .B1(ciphertext3[10]), .B2(ciphertext1[10]), .A(
        ciphertext2[10]), .ZN(mv_0_n22) );
  NAND2_X1 mv_0_U30 ( .A1(mv_0_n20), .A2(mv_0_n19), .ZN(ciphertext[9]) );
  NAND2_X1 mv_0_U29 ( .A1(ciphertext3[9]), .A2(ciphertext1[9]), .ZN(mv_0_n19)
         );
  OAI21_X1 mv_0_U28 ( .B1(ciphertext3[9]), .B2(ciphertext1[9]), .A(
        ciphertext2[9]), .ZN(mv_0_n20) );
  NAND2_X1 mv_0_U27 ( .A1(mv_0_n18), .A2(mv_0_n17), .ZN(ciphertext[8]) );
  NAND2_X1 mv_0_U26 ( .A1(ciphertext3[8]), .A2(ciphertext1[8]), .ZN(mv_0_n17)
         );
  OAI21_X1 mv_0_U25 ( .B1(ciphertext3[8]), .B2(ciphertext1[8]), .A(
        ciphertext2[8]), .ZN(mv_0_n18) );
  NAND2_X1 mv_0_U24 ( .A1(mv_0_n16), .A2(mv_0_n15), .ZN(ciphertext[7]) );
  NAND2_X1 mv_0_U23 ( .A1(ciphertext3[7]), .A2(ciphertext1[7]), .ZN(mv_0_n15)
         );
  OAI21_X1 mv_0_U22 ( .B1(ciphertext3[7]), .B2(ciphertext1[7]), .A(
        ciphertext2[7]), .ZN(mv_0_n16) );
  NAND2_X1 mv_0_U21 ( .A1(mv_0_n14), .A2(mv_0_n13), .ZN(ciphertext[6]) );
  NAND2_X1 mv_0_U20 ( .A1(ciphertext3[6]), .A2(ciphertext1[6]), .ZN(mv_0_n13)
         );
  OAI21_X1 mv_0_U19 ( .B1(ciphertext3[6]), .B2(ciphertext1[6]), .A(
        ciphertext2[6]), .ZN(mv_0_n14) );
  NAND2_X1 mv_0_U18 ( .A1(mv_0_n12), .A2(mv_0_n11), .ZN(ciphertext[5]) );
  NAND2_X1 mv_0_U17 ( .A1(ciphertext3[5]), .A2(ciphertext1[5]), .ZN(mv_0_n11)
         );
  OAI21_X1 mv_0_U16 ( .B1(ciphertext3[5]), .B2(ciphertext1[5]), .A(
        ciphertext2[5]), .ZN(mv_0_n12) );
  NAND2_X1 mv_0_U15 ( .A1(mv_0_n10), .A2(mv_0_n9), .ZN(ciphertext[4]) );
  NAND2_X1 mv_0_U14 ( .A1(ciphertext3[4]), .A2(ciphertext1[4]), .ZN(mv_0_n9)
         );
  OAI21_X1 mv_0_U13 ( .B1(ciphertext3[4]), .B2(ciphertext1[4]), .A(
        ciphertext2[4]), .ZN(mv_0_n10) );
  NAND2_X1 mv_0_U12 ( .A1(mv_0_n8), .A2(mv_0_n7), .ZN(ciphertext[3]) );
  NAND2_X1 mv_0_U11 ( .A1(ciphertext3[3]), .A2(ciphertext1[3]), .ZN(mv_0_n7)
         );
  OAI21_X1 mv_0_U10 ( .B1(ciphertext3[3]), .B2(ciphertext1[3]), .A(
        ciphertext2[3]), .ZN(mv_0_n8) );
  NAND2_X1 mv_0_U9 ( .A1(mv_0_n6), .A2(mv_0_n5), .ZN(ciphertext[2]) );
  NAND2_X1 mv_0_U8 ( .A1(ciphertext3[2]), .A2(ciphertext1[2]), .ZN(mv_0_n5) );
  OAI21_X1 mv_0_U7 ( .B1(ciphertext3[2]), .B2(ciphertext1[2]), .A(
        ciphertext2[2]), .ZN(mv_0_n6) );
  NAND2_X1 mv_0_U6 ( .A1(mv_0_n4), .A2(mv_0_n3), .ZN(ciphertext[1]) );
  NAND2_X1 mv_0_U5 ( .A1(ciphertext3[1]), .A2(ciphertext1[1]), .ZN(mv_0_n3) );
  OAI21_X1 mv_0_U4 ( .B1(ciphertext3[1]), .B2(ciphertext1[1]), .A(
        ciphertext2[1]), .ZN(mv_0_n4) );
  NAND2_X1 mv_0_U3 ( .A1(mv_0_n2), .A2(mv_0_n1), .ZN(ciphertext[0]) );
  NAND2_X1 mv_0_U2 ( .A1(ciphertext3[0]), .A2(ciphertext1[0]), .ZN(mv_0_n1) );
  OAI21_X1 mv_0_U1 ( .B1(ciphertext3[0]), .B2(ciphertext1[0]), .A(
        ciphertext2[0]), .ZN(mv_0_n2) );
  NAND2_X1 mv_1_U3 ( .A1(mv_1_n2), .A2(mv_1_n1), .ZN(done) );
  NAND2_X1 mv_1_U2 ( .A1(done3), .A2(done1), .ZN(mv_1_n1) );
  OAI21_X1 mv_1_U1 ( .B1(done3), .B2(done1), .A(done2), .ZN(mv_1_n2) );
endmodule

