
module circuit ( CLK, RESET, FRESH, DONE, KEY1, KEY2, KEY3, PLAINTEXT1, 
        PLAINTEXT2, PLAINTEXT3, CIPHERTEXT1, CIPHERTEXT2, CIPHERTEXT3 );
  input [127:0] FRESH;
  input [63:0] KEY1;
  input [63:0] KEY2;
  input [63:0] KEY3;
  input [63:0] PLAINTEXT1;
  input [63:0] PLAINTEXT2;
  input [63:0] PLAINTEXT3;
  output [63:0] CIPHERTEXT1;
  output [63:0] CIPHERTEXT2;
  output [63:0] CIPHERTEXT3;
  input CLK, RESET;
  output DONE;
  wire   KEY_EN, RF1_KA_n18, RF1_KA_n17, RF1_KA_n16, RF1_KA_n15, RF1_KA_n14,
         RF1_KA_n13, RF2_KA_n18, RF2_KA_n17, RF2_KA_n16, RF2_KA_n15,
         RF2_KA_n14, RF2_KA_n13, RF3_KA_n18, RF3_KA_n17, RF3_KA_n16,
         RF3_KA_n15, RF3_KA_n14, RF3_KA_n13, S_0_F_n4, S_0_F_n3, S_0_F_n2,
         S_0_F_n1, S_0_F_N5, S_0_F_N4, S_0_F_N3, S_0_F_N2, S_0_F_N1, S_0_F_N0,
         S_0_F_Inst_0__CF_Inst_n3, S_0_F_Inst_1__CF_Inst_n3,
         S_0_F_Inst_3__CF_Inst_n3, S_0_F_Inst_4__CF_Inst_n3,
         S_0_F_Inst_6__CF_Inst_n7, S_0_F_Inst_9__CF_Inst_n3,
         S_0_F_Inst_11__CF_Inst_n3, S_0_F_Inst_12__CF_Inst_n3,
         S_0_F_Inst_13__CF_Inst_n3, S_0_F_Inst_15__CF_Inst_n7,
         S_0_F_Inst_16__CF_Inst_n3, S_0_F_Inst_17__CF_Inst_n3,
         S_0_F_InstXOR_0__Compression1_n3, S_0_F_InstXOR_0__Compression2_n3,
         S_0_F_InstXOR_0__Compression3_n3, S_0_F_InstXOR_1__Compression1_n3,
         S_0_F_InstXOR_1__Compression2_n3, S_0_F_InstXOR_1__Compression3_n3,
         S_0_G_Inst_1__CF_Inst_n3, S_0_G_Inst_2__CF_Inst_n3,
         S_0_G_Inst_3__CF_Inst_n6, S_0_G_Inst_3__CF_Inst_n5,
         S_0_G_Inst_7__CF_Inst_n3, S_0_G_Inst_9__CF_Inst_n3,
         S_0_G_Inst_10__CF_Inst_n3, S_0_G_Inst_11__CF_Inst_n6,
         S_0_G_Inst_11__CF_Inst_n5, S_0_G_Inst_12__CF_Inst_n3,
         S_0_G_Inst_14__CF_Inst_n6, S_0_G_Inst_14__CF_Inst_n5,
         S_0_G_Inst_15__CF_Inst_n3, S_0_G_Inst_17__CF_Inst_n3,
         S_0_G_InstXOR_0__Compression1_n3, S_0_G_InstXOR_0__Compression2_n3,
         S_0_G_InstXOR_0__Compression3_n3, S_0_G_InstXOR_1__Compression1_n3,
         S_0_G_InstXOR_1__Compression2_n3, S_0_G_InstXOR_1__Compression3_n3,
         S_1_F_n12, S_1_F_n11, S_1_F_n10, S_1_F_n9, S_1_F_N5, S_1_F_N4,
         S_1_F_N3, S_1_F_N2, S_1_F_N1, S_1_F_N0, S_1_F_Inst_0__CF_Inst_n3,
         S_1_F_Inst_1__CF_Inst_n3, S_1_F_Inst_3__CF_Inst_n3,
         S_1_F_Inst_4__CF_Inst_n3, S_1_F_Inst_6__CF_Inst_n7,
         S_1_F_Inst_9__CF_Inst_n3, S_1_F_Inst_11__CF_Inst_n3,
         S_1_F_Inst_12__CF_Inst_n3, S_1_F_Inst_13__CF_Inst_n3,
         S_1_F_Inst_15__CF_Inst_n7, S_1_F_Inst_16__CF_Inst_n3,
         S_1_F_Inst_17__CF_Inst_n3, S_1_F_InstXOR_0__Compression1_n3,
         S_1_F_InstXOR_0__Compression2_n3, S_1_F_InstXOR_0__Compression3_n3,
         S_1_F_InstXOR_1__Compression1_n3, S_1_F_InstXOR_1__Compression2_n3,
         S_1_F_InstXOR_1__Compression3_n3, S_1_G_Inst_1__CF_Inst_n3,
         S_1_G_Inst_2__CF_Inst_n3, S_1_G_Inst_3__CF_Inst_n6,
         S_1_G_Inst_3__CF_Inst_n5, S_1_G_Inst_7__CF_Inst_n3,
         S_1_G_Inst_9__CF_Inst_n3, S_1_G_Inst_10__CF_Inst_n3,
         S_1_G_Inst_11__CF_Inst_n6, S_1_G_Inst_11__CF_Inst_n5,
         S_1_G_Inst_12__CF_Inst_n3, S_1_G_Inst_14__CF_Inst_n6,
         S_1_G_Inst_14__CF_Inst_n5, S_1_G_Inst_15__CF_Inst_n3,
         S_1_G_Inst_17__CF_Inst_n3, S_1_G_InstXOR_0__Compression1_n3,
         S_1_G_InstXOR_0__Compression2_n3, S_1_G_InstXOR_0__Compression3_n3,
         S_1_G_InstXOR_1__Compression1_n3, S_1_G_InstXOR_1__Compression2_n3,
         S_1_G_InstXOR_1__Compression3_n3, S_2_F_n12, S_2_F_n11, S_2_F_n10,
         S_2_F_n9, S_2_F_N5, S_2_F_N4, S_2_F_N3, S_2_F_N2, S_2_F_N1, S_2_F_N0,
         S_2_F_Inst_0__CF_Inst_n3, S_2_F_Inst_1__CF_Inst_n3,
         S_2_F_Inst_3__CF_Inst_n3, S_2_F_Inst_4__CF_Inst_n3,
         S_2_F_Inst_6__CF_Inst_n7, S_2_F_Inst_9__CF_Inst_n3,
         S_2_F_Inst_11__CF_Inst_n3, S_2_F_Inst_12__CF_Inst_n3,
         S_2_F_Inst_13__CF_Inst_n3, S_2_F_Inst_15__CF_Inst_n7,
         S_2_F_Inst_16__CF_Inst_n3, S_2_F_Inst_17__CF_Inst_n3,
         S_2_F_InstXOR_0__Compression1_n3, S_2_F_InstXOR_0__Compression2_n3,
         S_2_F_InstXOR_0__Compression3_n3, S_2_F_InstXOR_1__Compression1_n3,
         S_2_F_InstXOR_1__Compression2_n3, S_2_F_InstXOR_1__Compression3_n3,
         S_2_G_Inst_1__CF_Inst_n3, S_2_G_Inst_2__CF_Inst_n3,
         S_2_G_Inst_3__CF_Inst_n6, S_2_G_Inst_3__CF_Inst_n5,
         S_2_G_Inst_7__CF_Inst_n3, S_2_G_Inst_9__CF_Inst_n3,
         S_2_G_Inst_10__CF_Inst_n3, S_2_G_Inst_11__CF_Inst_n6,
         S_2_G_Inst_11__CF_Inst_n5, S_2_G_Inst_12__CF_Inst_n3,
         S_2_G_Inst_14__CF_Inst_n6, S_2_G_Inst_14__CF_Inst_n5,
         S_2_G_Inst_15__CF_Inst_n3, S_2_G_Inst_17__CF_Inst_n3,
         S_2_G_InstXOR_0__Compression1_n3, S_2_G_InstXOR_0__Compression2_n3,
         S_2_G_InstXOR_0__Compression3_n3, S_2_G_InstXOR_1__Compression1_n3,
         S_2_G_InstXOR_1__Compression2_n3, S_2_G_InstXOR_1__Compression3_n3,
         S_3_F_n12, S_3_F_n11, S_3_F_n10, S_3_F_n9, S_3_F_N5, S_3_F_N4,
         S_3_F_N3, S_3_F_N2, S_3_F_N1, S_3_F_N0, S_3_F_Inst_0__CF_Inst_n3,
         S_3_F_Inst_1__CF_Inst_n3, S_3_F_Inst_3__CF_Inst_n3,
         S_3_F_Inst_4__CF_Inst_n3, S_3_F_Inst_6__CF_Inst_n7,
         S_3_F_Inst_9__CF_Inst_n3, S_3_F_Inst_11__CF_Inst_n3,
         S_3_F_Inst_12__CF_Inst_n3, S_3_F_Inst_13__CF_Inst_n3,
         S_3_F_Inst_15__CF_Inst_n7, S_3_F_Inst_16__CF_Inst_n3,
         S_3_F_Inst_17__CF_Inst_n3, S_3_F_InstXOR_0__Compression1_n3,
         S_3_F_InstXOR_0__Compression2_n3, S_3_F_InstXOR_0__Compression3_n3,
         S_3_F_InstXOR_1__Compression1_n3, S_3_F_InstXOR_1__Compression2_n3,
         S_3_F_InstXOR_1__Compression3_n3, S_3_G_Inst_1__CF_Inst_n3,
         S_3_G_Inst_2__CF_Inst_n3, S_3_G_Inst_3__CF_Inst_n6,
         S_3_G_Inst_3__CF_Inst_n5, S_3_G_Inst_7__CF_Inst_n3,
         S_3_G_Inst_9__CF_Inst_n3, S_3_G_Inst_10__CF_Inst_n3,
         S_3_G_Inst_11__CF_Inst_n6, S_3_G_Inst_11__CF_Inst_n5,
         S_3_G_Inst_12__CF_Inst_n3, S_3_G_Inst_14__CF_Inst_n6,
         S_3_G_Inst_14__CF_Inst_n5, S_3_G_Inst_15__CF_Inst_n3,
         S_3_G_Inst_17__CF_Inst_n3, S_3_G_InstXOR_0__Compression1_n3,
         S_3_G_InstXOR_0__Compression2_n3, S_3_G_InstXOR_0__Compression3_n3,
         S_3_G_InstXOR_1__Compression1_n3, S_3_G_InstXOR_1__Compression2_n3,
         S_3_G_InstXOR_1__Compression3_n3, S_4_F_n12, S_4_F_n11, S_4_F_n10,
         S_4_F_n9, S_4_F_N5, S_4_F_N4, S_4_F_N3, S_4_F_N2, S_4_F_N1, S_4_F_N0,
         S_4_F_Inst_0__CF_Inst_n3, S_4_F_Inst_1__CF_Inst_n3,
         S_4_F_Inst_3__CF_Inst_n3, S_4_F_Inst_4__CF_Inst_n3,
         S_4_F_Inst_6__CF_Inst_n7, S_4_F_Inst_9__CF_Inst_n3,
         S_4_F_Inst_11__CF_Inst_n3, S_4_F_Inst_12__CF_Inst_n3,
         S_4_F_Inst_13__CF_Inst_n3, S_4_F_Inst_15__CF_Inst_n7,
         S_4_F_Inst_16__CF_Inst_n3, S_4_F_Inst_17__CF_Inst_n3,
         S_4_F_InstXOR_0__Compression1_n3, S_4_F_InstXOR_0__Compression2_n3,
         S_4_F_InstXOR_0__Compression3_n3, S_4_F_InstXOR_1__Compression1_n3,
         S_4_F_InstXOR_1__Compression2_n3, S_4_F_InstXOR_1__Compression3_n3,
         S_4_G_Inst_1__CF_Inst_n3, S_4_G_Inst_2__CF_Inst_n3,
         S_4_G_Inst_3__CF_Inst_n6, S_4_G_Inst_3__CF_Inst_n5,
         S_4_G_Inst_7__CF_Inst_n3, S_4_G_Inst_9__CF_Inst_n3,
         S_4_G_Inst_10__CF_Inst_n3, S_4_G_Inst_11__CF_Inst_n6,
         S_4_G_Inst_11__CF_Inst_n5, S_4_G_Inst_12__CF_Inst_n3,
         S_4_G_Inst_14__CF_Inst_n6, S_4_G_Inst_14__CF_Inst_n5,
         S_4_G_Inst_15__CF_Inst_n3, S_4_G_Inst_17__CF_Inst_n3,
         S_4_G_InstXOR_0__Compression1_n3, S_4_G_InstXOR_0__Compression2_n3,
         S_4_G_InstXOR_0__Compression3_n3, S_4_G_InstXOR_1__Compression1_n3,
         S_4_G_InstXOR_1__Compression2_n3, S_4_G_InstXOR_1__Compression3_n3,
         S_5_F_n12, S_5_F_n11, S_5_F_n10, S_5_F_n9, S_5_F_N5, S_5_F_N4,
         S_5_F_N3, S_5_F_N2, S_5_F_N1, S_5_F_N0, S_5_F_Inst_0__CF_Inst_n3,
         S_5_F_Inst_1__CF_Inst_n3, S_5_F_Inst_3__CF_Inst_n3,
         S_5_F_Inst_4__CF_Inst_n3, S_5_F_Inst_6__CF_Inst_n7,
         S_5_F_Inst_9__CF_Inst_n3, S_5_F_Inst_11__CF_Inst_n3,
         S_5_F_Inst_12__CF_Inst_n3, S_5_F_Inst_13__CF_Inst_n3,
         S_5_F_Inst_15__CF_Inst_n7, S_5_F_Inst_16__CF_Inst_n3,
         S_5_F_Inst_17__CF_Inst_n3, S_5_F_InstXOR_0__Compression1_n3,
         S_5_F_InstXOR_0__Compression2_n3, S_5_F_InstXOR_0__Compression3_n3,
         S_5_F_InstXOR_1__Compression1_n3, S_5_F_InstXOR_1__Compression2_n3,
         S_5_F_InstXOR_1__Compression3_n3, S_5_G_Inst_1__CF_Inst_n3,
         S_5_G_Inst_2__CF_Inst_n3, S_5_G_Inst_3__CF_Inst_n6,
         S_5_G_Inst_3__CF_Inst_n5, S_5_G_Inst_7__CF_Inst_n3,
         S_5_G_Inst_9__CF_Inst_n3, S_5_G_Inst_10__CF_Inst_n3,
         S_5_G_Inst_11__CF_Inst_n6, S_5_G_Inst_11__CF_Inst_n5,
         S_5_G_Inst_12__CF_Inst_n3, S_5_G_Inst_14__CF_Inst_n6,
         S_5_G_Inst_14__CF_Inst_n5, S_5_G_Inst_15__CF_Inst_n3,
         S_5_G_Inst_17__CF_Inst_n3, S_5_G_InstXOR_0__Compression1_n3,
         S_5_G_InstXOR_0__Compression2_n3, S_5_G_InstXOR_0__Compression3_n3,
         S_5_G_InstXOR_1__Compression1_n3, S_5_G_InstXOR_1__Compression2_n3,
         S_5_G_InstXOR_1__Compression3_n3, S_6_F_n12, S_6_F_n11, S_6_F_n10,
         S_6_F_n9, S_6_F_N5, S_6_F_N4, S_6_F_N3, S_6_F_N2, S_6_F_N1, S_6_F_N0,
         S_6_F_Inst_0__CF_Inst_n3, S_6_F_Inst_1__CF_Inst_n3,
         S_6_F_Inst_3__CF_Inst_n3, S_6_F_Inst_4__CF_Inst_n3,
         S_6_F_Inst_6__CF_Inst_n7, S_6_F_Inst_9__CF_Inst_n3,
         S_6_F_Inst_11__CF_Inst_n3, S_6_F_Inst_12__CF_Inst_n3,
         S_6_F_Inst_13__CF_Inst_n3, S_6_F_Inst_15__CF_Inst_n7,
         S_6_F_Inst_16__CF_Inst_n3, S_6_F_Inst_17__CF_Inst_n3,
         S_6_F_InstXOR_0__Compression1_n3, S_6_F_InstXOR_0__Compression2_n3,
         S_6_F_InstXOR_0__Compression3_n3, S_6_F_InstXOR_1__Compression1_n3,
         S_6_F_InstXOR_1__Compression2_n3, S_6_F_InstXOR_1__Compression3_n3,
         S_6_G_Inst_1__CF_Inst_n3, S_6_G_Inst_2__CF_Inst_n3,
         S_6_G_Inst_3__CF_Inst_n6, S_6_G_Inst_3__CF_Inst_n5,
         S_6_G_Inst_7__CF_Inst_n3, S_6_G_Inst_9__CF_Inst_n3,
         S_6_G_Inst_10__CF_Inst_n3, S_6_G_Inst_11__CF_Inst_n6,
         S_6_G_Inst_11__CF_Inst_n5, S_6_G_Inst_12__CF_Inst_n3,
         S_6_G_Inst_14__CF_Inst_n6, S_6_G_Inst_14__CF_Inst_n5,
         S_6_G_Inst_15__CF_Inst_n3, S_6_G_Inst_17__CF_Inst_n3,
         S_6_G_InstXOR_0__Compression1_n3, S_6_G_InstXOR_0__Compression2_n3,
         S_6_G_InstXOR_0__Compression3_n3, S_6_G_InstXOR_1__Compression1_n3,
         S_6_G_InstXOR_1__Compression2_n3, S_6_G_InstXOR_1__Compression3_n3,
         S_7_F_n12, S_7_F_n11, S_7_F_n10, S_7_F_n9, S_7_F_N5, S_7_F_N4,
         S_7_F_N3, S_7_F_N2, S_7_F_N1, S_7_F_N0, S_7_F_Inst_0__CF_Inst_n3,
         S_7_F_Inst_1__CF_Inst_n3, S_7_F_Inst_3__CF_Inst_n3,
         S_7_F_Inst_4__CF_Inst_n3, S_7_F_Inst_6__CF_Inst_n7,
         S_7_F_Inst_9__CF_Inst_n3, S_7_F_Inst_11__CF_Inst_n3,
         S_7_F_Inst_12__CF_Inst_n3, S_7_F_Inst_13__CF_Inst_n3,
         S_7_F_Inst_15__CF_Inst_n7, S_7_F_Inst_16__CF_Inst_n3,
         S_7_F_Inst_17__CF_Inst_n3, S_7_F_InstXOR_0__Compression1_n3,
         S_7_F_InstXOR_0__Compression2_n3, S_7_F_InstXOR_0__Compression3_n3,
         S_7_F_InstXOR_1__Compression1_n3, S_7_F_InstXOR_1__Compression2_n3,
         S_7_F_InstXOR_1__Compression3_n3, S_7_G_Inst_1__CF_Inst_n3,
         S_7_G_Inst_2__CF_Inst_n3, S_7_G_Inst_3__CF_Inst_n6,
         S_7_G_Inst_3__CF_Inst_n5, S_7_G_Inst_7__CF_Inst_n3,
         S_7_G_Inst_9__CF_Inst_n3, S_7_G_Inst_10__CF_Inst_n3,
         S_7_G_Inst_11__CF_Inst_n6, S_7_G_Inst_11__CF_Inst_n5,
         S_7_G_Inst_12__CF_Inst_n3, S_7_G_Inst_14__CF_Inst_n6,
         S_7_G_Inst_14__CF_Inst_n5, S_7_G_Inst_15__CF_Inst_n3,
         S_7_G_Inst_17__CF_Inst_n3, S_7_G_InstXOR_0__Compression1_n3,
         S_7_G_InstXOR_0__Compression2_n3, S_7_G_InstXOR_0__Compression3_n3,
         S_7_G_InstXOR_1__Compression1_n3, S_7_G_InstXOR_1__Compression2_n3,
         S_7_G_InstXOR_1__Compression3_n3, S_8_F_n12, S_8_F_n11, S_8_F_n10,
         S_8_F_n9, S_8_F_N5, S_8_F_N4, S_8_F_N3, S_8_F_N2, S_8_F_N1, S_8_F_N0,
         S_8_F_Inst_0__CF_Inst_n3, S_8_F_Inst_1__CF_Inst_n3,
         S_8_F_Inst_3__CF_Inst_n3, S_8_F_Inst_4__CF_Inst_n3,
         S_8_F_Inst_6__CF_Inst_n7, S_8_F_Inst_9__CF_Inst_n3,
         S_8_F_Inst_11__CF_Inst_n3, S_8_F_Inst_12__CF_Inst_n3,
         S_8_F_Inst_13__CF_Inst_n3, S_8_F_Inst_15__CF_Inst_n7,
         S_8_F_Inst_16__CF_Inst_n3, S_8_F_Inst_17__CF_Inst_n3,
         S_8_F_InstXOR_0__Compression1_n3, S_8_F_InstXOR_0__Compression2_n3,
         S_8_F_InstXOR_0__Compression3_n3, S_8_F_InstXOR_1__Compression1_n3,
         S_8_F_InstXOR_1__Compression2_n3, S_8_F_InstXOR_1__Compression3_n3,
         S_8_G_Inst_1__CF_Inst_n3, S_8_G_Inst_2__CF_Inst_n3,
         S_8_G_Inst_3__CF_Inst_n6, S_8_G_Inst_3__CF_Inst_n5,
         S_8_G_Inst_7__CF_Inst_n3, S_8_G_Inst_9__CF_Inst_n3,
         S_8_G_Inst_10__CF_Inst_n3, S_8_G_Inst_11__CF_Inst_n6,
         S_8_G_Inst_11__CF_Inst_n5, S_8_G_Inst_12__CF_Inst_n3,
         S_8_G_Inst_14__CF_Inst_n6, S_8_G_Inst_14__CF_Inst_n5,
         S_8_G_Inst_15__CF_Inst_n3, S_8_G_Inst_17__CF_Inst_n3,
         S_8_G_InstXOR_0__Compression1_n3, S_8_G_InstXOR_0__Compression2_n3,
         S_8_G_InstXOR_0__Compression3_n3, S_8_G_InstXOR_1__Compression1_n3,
         S_8_G_InstXOR_1__Compression2_n3, S_8_G_InstXOR_1__Compression3_n3,
         S_9_F_n12, S_9_F_n11, S_9_F_n10, S_9_F_n9, S_9_F_N5, S_9_F_N4,
         S_9_F_N3, S_9_F_N2, S_9_F_N1, S_9_F_N0, S_9_F_Inst_0__CF_Inst_n3,
         S_9_F_Inst_1__CF_Inst_n3, S_9_F_Inst_3__CF_Inst_n3,
         S_9_F_Inst_4__CF_Inst_n3, S_9_F_Inst_6__CF_Inst_n7,
         S_9_F_Inst_9__CF_Inst_n3, S_9_F_Inst_11__CF_Inst_n3,
         S_9_F_Inst_12__CF_Inst_n3, S_9_F_Inst_13__CF_Inst_n3,
         S_9_F_Inst_15__CF_Inst_n7, S_9_F_Inst_16__CF_Inst_n3,
         S_9_F_Inst_17__CF_Inst_n3, S_9_F_InstXOR_0__Compression1_n3,
         S_9_F_InstXOR_0__Compression2_n3, S_9_F_InstXOR_0__Compression3_n3,
         S_9_F_InstXOR_1__Compression1_n3, S_9_F_InstXOR_1__Compression2_n3,
         S_9_F_InstXOR_1__Compression3_n3, S_9_G_Inst_1__CF_Inst_n3,
         S_9_G_Inst_2__CF_Inst_n3, S_9_G_Inst_3__CF_Inst_n6,
         S_9_G_Inst_3__CF_Inst_n5, S_9_G_Inst_7__CF_Inst_n3,
         S_9_G_Inst_9__CF_Inst_n3, S_9_G_Inst_10__CF_Inst_n3,
         S_9_G_Inst_11__CF_Inst_n6, S_9_G_Inst_11__CF_Inst_n5,
         S_9_G_Inst_12__CF_Inst_n3, S_9_G_Inst_14__CF_Inst_n6,
         S_9_G_Inst_14__CF_Inst_n5, S_9_G_Inst_15__CF_Inst_n3,
         S_9_G_Inst_17__CF_Inst_n3, S_9_G_InstXOR_0__Compression1_n3,
         S_9_G_InstXOR_0__Compression2_n3, S_9_G_InstXOR_0__Compression3_n3,
         S_9_G_InstXOR_1__Compression1_n3, S_9_G_InstXOR_1__Compression2_n3,
         S_9_G_InstXOR_1__Compression3_n3, S_10_F_n12, S_10_F_n11, S_10_F_n10,
         S_10_F_n9, S_10_F_N5, S_10_F_N4, S_10_F_N3, S_10_F_N2, S_10_F_N1,
         S_10_F_N0, S_10_F_Inst_0__CF_Inst_n3, S_10_F_Inst_1__CF_Inst_n3,
         S_10_F_Inst_3__CF_Inst_n3, S_10_F_Inst_4__CF_Inst_n3,
         S_10_F_Inst_6__CF_Inst_n7, S_10_F_Inst_9__CF_Inst_n3,
         S_10_F_Inst_11__CF_Inst_n3, S_10_F_Inst_12__CF_Inst_n3,
         S_10_F_Inst_13__CF_Inst_n3, S_10_F_Inst_15__CF_Inst_n7,
         S_10_F_Inst_16__CF_Inst_n3, S_10_F_Inst_17__CF_Inst_n3,
         S_10_F_InstXOR_0__Compression1_n3, S_10_F_InstXOR_0__Compression2_n3,
         S_10_F_InstXOR_0__Compression3_n3, S_10_F_InstXOR_1__Compression1_n3,
         S_10_F_InstXOR_1__Compression2_n3, S_10_F_InstXOR_1__Compression3_n3,
         S_10_G_Inst_1__CF_Inst_n3, S_10_G_Inst_2__CF_Inst_n3,
         S_10_G_Inst_3__CF_Inst_n6, S_10_G_Inst_3__CF_Inst_n5,
         S_10_G_Inst_7__CF_Inst_n3, S_10_G_Inst_9__CF_Inst_n3,
         S_10_G_Inst_10__CF_Inst_n3, S_10_G_Inst_11__CF_Inst_n6,
         S_10_G_Inst_11__CF_Inst_n5, S_10_G_Inst_12__CF_Inst_n3,
         S_10_G_Inst_14__CF_Inst_n6, S_10_G_Inst_14__CF_Inst_n5,
         S_10_G_Inst_15__CF_Inst_n3, S_10_G_Inst_17__CF_Inst_n3,
         S_10_G_InstXOR_0__Compression1_n3, S_10_G_InstXOR_0__Compression2_n3,
         S_10_G_InstXOR_0__Compression3_n3, S_10_G_InstXOR_1__Compression1_n3,
         S_10_G_InstXOR_1__Compression2_n3, S_10_G_InstXOR_1__Compression3_n3,
         S_11_F_n12, S_11_F_n11, S_11_F_n10, S_11_F_n9, S_11_F_N5, S_11_F_N4,
         S_11_F_N3, S_11_F_N2, S_11_F_N1, S_11_F_N0, S_11_F_Inst_0__CF_Inst_n3,
         S_11_F_Inst_1__CF_Inst_n3, S_11_F_Inst_3__CF_Inst_n3,
         S_11_F_Inst_4__CF_Inst_n3, S_11_F_Inst_6__CF_Inst_n7,
         S_11_F_Inst_9__CF_Inst_n3, S_11_F_Inst_11__CF_Inst_n3,
         S_11_F_Inst_12__CF_Inst_n3, S_11_F_Inst_13__CF_Inst_n3,
         S_11_F_Inst_15__CF_Inst_n7, S_11_F_Inst_16__CF_Inst_n3,
         S_11_F_Inst_17__CF_Inst_n3, S_11_F_InstXOR_0__Compression1_n3,
         S_11_F_InstXOR_0__Compression2_n3, S_11_F_InstXOR_0__Compression3_n3,
         S_11_F_InstXOR_1__Compression1_n3, S_11_F_InstXOR_1__Compression2_n3,
         S_11_F_InstXOR_1__Compression3_n3, S_11_G_Inst_1__CF_Inst_n3,
         S_11_G_Inst_2__CF_Inst_n3, S_11_G_Inst_3__CF_Inst_n6,
         S_11_G_Inst_3__CF_Inst_n5, S_11_G_Inst_7__CF_Inst_n3,
         S_11_G_Inst_9__CF_Inst_n3, S_11_G_Inst_10__CF_Inst_n3,
         S_11_G_Inst_11__CF_Inst_n6, S_11_G_Inst_11__CF_Inst_n5,
         S_11_G_Inst_12__CF_Inst_n3, S_11_G_Inst_14__CF_Inst_n6,
         S_11_G_Inst_14__CF_Inst_n5, S_11_G_Inst_15__CF_Inst_n3,
         S_11_G_Inst_17__CF_Inst_n3, S_11_G_InstXOR_0__Compression1_n3,
         S_11_G_InstXOR_0__Compression2_n3, S_11_G_InstXOR_0__Compression3_n3,
         S_11_G_InstXOR_1__Compression1_n3, S_11_G_InstXOR_1__Compression2_n3,
         S_11_G_InstXOR_1__Compression3_n3, S_12_F_n12, S_12_F_n11, S_12_F_n10,
         S_12_F_n9, S_12_F_N5, S_12_F_N4, S_12_F_N3, S_12_F_N2, S_12_F_N1,
         S_12_F_N0, S_12_F_Inst_0__CF_Inst_n3, S_12_F_Inst_1__CF_Inst_n3,
         S_12_F_Inst_3__CF_Inst_n3, S_12_F_Inst_4__CF_Inst_n3,
         S_12_F_Inst_6__CF_Inst_n7, S_12_F_Inst_9__CF_Inst_n3,
         S_12_F_Inst_11__CF_Inst_n3, S_12_F_Inst_12__CF_Inst_n3,
         S_12_F_Inst_13__CF_Inst_n3, S_12_F_Inst_15__CF_Inst_n7,
         S_12_F_Inst_16__CF_Inst_n3, S_12_F_Inst_17__CF_Inst_n3,
         S_12_F_InstXOR_0__Compression1_n3, S_12_F_InstXOR_0__Compression2_n3,
         S_12_F_InstXOR_0__Compression3_n3, S_12_F_InstXOR_1__Compression1_n3,
         S_12_F_InstXOR_1__Compression2_n3, S_12_F_InstXOR_1__Compression3_n3,
         S_12_G_Inst_1__CF_Inst_n3, S_12_G_Inst_2__CF_Inst_n3,
         S_12_G_Inst_3__CF_Inst_n6, S_12_G_Inst_3__CF_Inst_n5,
         S_12_G_Inst_7__CF_Inst_n3, S_12_G_Inst_9__CF_Inst_n3,
         S_12_G_Inst_10__CF_Inst_n3, S_12_G_Inst_11__CF_Inst_n6,
         S_12_G_Inst_11__CF_Inst_n5, S_12_G_Inst_12__CF_Inst_n3,
         S_12_G_Inst_14__CF_Inst_n6, S_12_G_Inst_14__CF_Inst_n5,
         S_12_G_Inst_15__CF_Inst_n3, S_12_G_Inst_17__CF_Inst_n3,
         S_12_G_InstXOR_0__Compression1_n3, S_12_G_InstXOR_0__Compression2_n3,
         S_12_G_InstXOR_0__Compression3_n3, S_12_G_InstXOR_1__Compression1_n3,
         S_12_G_InstXOR_1__Compression2_n3, S_12_G_InstXOR_1__Compression3_n3,
         S_13_F_n12, S_13_F_n11, S_13_F_n10, S_13_F_n9, S_13_F_N5, S_13_F_N4,
         S_13_F_N3, S_13_F_N2, S_13_F_N1, S_13_F_N0, S_13_F_Inst_0__CF_Inst_n3,
         S_13_F_Inst_1__CF_Inst_n3, S_13_F_Inst_3__CF_Inst_n3,
         S_13_F_Inst_4__CF_Inst_n3, S_13_F_Inst_6__CF_Inst_n7,
         S_13_F_Inst_9__CF_Inst_n3, S_13_F_Inst_11__CF_Inst_n3,
         S_13_F_Inst_12__CF_Inst_n3, S_13_F_Inst_13__CF_Inst_n3,
         S_13_F_Inst_15__CF_Inst_n7, S_13_F_Inst_16__CF_Inst_n3,
         S_13_F_Inst_17__CF_Inst_n3, S_13_F_InstXOR_0__Compression1_n3,
         S_13_F_InstXOR_0__Compression2_n3, S_13_F_InstXOR_0__Compression3_n3,
         S_13_F_InstXOR_1__Compression1_n3, S_13_F_InstXOR_1__Compression2_n3,
         S_13_F_InstXOR_1__Compression3_n3, S_13_G_Inst_1__CF_Inst_n3,
         S_13_G_Inst_2__CF_Inst_n3, S_13_G_Inst_3__CF_Inst_n6,
         S_13_G_Inst_3__CF_Inst_n5, S_13_G_Inst_7__CF_Inst_n3,
         S_13_G_Inst_9__CF_Inst_n3, S_13_G_Inst_10__CF_Inst_n3,
         S_13_G_Inst_11__CF_Inst_n6, S_13_G_Inst_11__CF_Inst_n5,
         S_13_G_Inst_12__CF_Inst_n3, S_13_G_Inst_14__CF_Inst_n6,
         S_13_G_Inst_14__CF_Inst_n5, S_13_G_Inst_15__CF_Inst_n3,
         S_13_G_Inst_17__CF_Inst_n3, S_13_G_InstXOR_0__Compression1_n3,
         S_13_G_InstXOR_0__Compression2_n3, S_13_G_InstXOR_0__Compression3_n3,
         S_13_G_InstXOR_1__Compression1_n3, S_13_G_InstXOR_1__Compression2_n3,
         S_13_G_InstXOR_1__Compression3_n3, S_14_F_n12, S_14_F_n11, S_14_F_n10,
         S_14_F_n9, S_14_F_N5, S_14_F_N4, S_14_F_N3, S_14_F_N2, S_14_F_N1,
         S_14_F_N0, S_14_F_Inst_0__CF_Inst_n3, S_14_F_Inst_1__CF_Inst_n3,
         S_14_F_Inst_3__CF_Inst_n3, S_14_F_Inst_4__CF_Inst_n3,
         S_14_F_Inst_6__CF_Inst_n7, S_14_F_Inst_9__CF_Inst_n3,
         S_14_F_Inst_11__CF_Inst_n3, S_14_F_Inst_12__CF_Inst_n3,
         S_14_F_Inst_13__CF_Inst_n3, S_14_F_Inst_15__CF_Inst_n7,
         S_14_F_Inst_16__CF_Inst_n3, S_14_F_Inst_17__CF_Inst_n3,
         S_14_F_InstXOR_0__Compression1_n3, S_14_F_InstXOR_0__Compression2_n3,
         S_14_F_InstXOR_0__Compression3_n3, S_14_F_InstXOR_1__Compression1_n3,
         S_14_F_InstXOR_1__Compression2_n3, S_14_F_InstXOR_1__Compression3_n3,
         S_14_G_Inst_1__CF_Inst_n3, S_14_G_Inst_2__CF_Inst_n3,
         S_14_G_Inst_3__CF_Inst_n6, S_14_G_Inst_3__CF_Inst_n5,
         S_14_G_Inst_7__CF_Inst_n3, S_14_G_Inst_9__CF_Inst_n3,
         S_14_G_Inst_10__CF_Inst_n3, S_14_G_Inst_11__CF_Inst_n6,
         S_14_G_Inst_11__CF_Inst_n5, S_14_G_Inst_12__CF_Inst_n3,
         S_14_G_Inst_14__CF_Inst_n6, S_14_G_Inst_14__CF_Inst_n5,
         S_14_G_Inst_15__CF_Inst_n3, S_14_G_Inst_17__CF_Inst_n3,
         S_14_G_InstXOR_0__Compression1_n3, S_14_G_InstXOR_0__Compression2_n3,
         S_14_G_InstXOR_0__Compression3_n3, S_14_G_InstXOR_1__Compression1_n3,
         S_14_G_InstXOR_1__Compression2_n3, S_14_G_InstXOR_1__Compression3_n3,
         S_15_F_n12, S_15_F_n11, S_15_F_n10, S_15_F_n9, S_15_F_N5, S_15_F_N4,
         S_15_F_N3, S_15_F_N2, S_15_F_N1, S_15_F_N0, S_15_F_Inst_0__CF_Inst_n3,
         S_15_F_Inst_1__CF_Inst_n3, S_15_F_Inst_3__CF_Inst_n3,
         S_15_F_Inst_4__CF_Inst_n3, S_15_F_Inst_6__CF_Inst_n7,
         S_15_F_Inst_9__CF_Inst_n3, S_15_F_Inst_11__CF_Inst_n3,
         S_15_F_Inst_12__CF_Inst_n3, S_15_F_Inst_13__CF_Inst_n3,
         S_15_F_Inst_15__CF_Inst_n7, S_15_F_Inst_16__CF_Inst_n3,
         S_15_F_Inst_17__CF_Inst_n3, S_15_F_InstXOR_0__Compression1_n3,
         S_15_F_InstXOR_0__Compression2_n3, S_15_F_InstXOR_0__Compression3_n3,
         S_15_F_InstXOR_1__Compression1_n3, S_15_F_InstXOR_1__Compression2_n3,
         S_15_F_InstXOR_1__Compression3_n3, S_15_G_Inst_1__CF_Inst_n3,
         S_15_G_Inst_2__CF_Inst_n3, S_15_G_Inst_3__CF_Inst_n6,
         S_15_G_Inst_3__CF_Inst_n5, S_15_G_Inst_7__CF_Inst_n3,
         S_15_G_Inst_9__CF_Inst_n3, S_15_G_Inst_10__CF_Inst_n3,
         S_15_G_Inst_11__CF_Inst_n6, S_15_G_Inst_11__CF_Inst_n5,
         S_15_G_Inst_12__CF_Inst_n3, S_15_G_Inst_14__CF_Inst_n6,
         S_15_G_Inst_14__CF_Inst_n5, S_15_G_Inst_15__CF_Inst_n3,
         S_15_G_Inst_17__CF_Inst_n3, S_15_G_InstXOR_0__Compression1_n3,
         S_15_G_InstXOR_0__Compression2_n3, S_15_G_InstXOR_0__Compression3_n3,
         S_15_G_InstXOR_1__Compression1_n3, S_15_G_InstXOR_1__Compression2_n3,
         S_15_G_InstXOR_1__Compression3_n3, KE1_RS_n12, KE1_RS_n11, KE1_RS_n10,
         KE1_RS_n9, KE1_RS_n8, KE1_RS_n7, KE1_RS_SFF_0_n10, KE1_RS_SFF_0_n9,
         KE1_RS_SFF_0_n7, KE1_RS_SFF_0_n6, KE1_RS_SFF_1_n11, KE1_RS_SFF_1_n10,
         KE1_RS_SFF_1_n8, KE1_RS_SFF_1_n7, KE1_RS_SFF_2_n11, KE1_RS_SFF_2_n10,
         KE1_RS_SFF_2_n8, KE1_RS_SFF_2_n7, KE1_RS_SFF_3_n10, KE1_RS_SFF_3_n9,
         KE1_RS_SFF_3_n7, KE1_RS_SFF_3_n6, KE1_RS_SFF_4_n10, KE1_RS_SFF_4_n9,
         KE1_RS_SFF_4_n7, KE1_RS_SFF_4_n6, KE1_RS_SFF_5_n10, KE1_RS_SFF_5_n9,
         KE1_RS_SFF_5_n7, KE1_RS_SFF_5_n6, KE1_RS_SFF_6_n10, KE1_RS_SFF_6_n9,
         KE1_RS_SFF_6_n7, KE1_RS_SFF_6_n6, KE1_RS_SFF_7_n10, KE1_RS_SFF_7_n9,
         KE1_RS_SFF_7_n7, KE1_RS_SFF_7_n6, KE1_RS_SFF_8_n10, KE1_RS_SFF_8_n9,
         KE1_RS_SFF_8_n7, KE1_RS_SFF_8_n6, KE1_RS_SFF_9_n10, KE1_RS_SFF_9_n9,
         KE1_RS_SFF_9_n7, KE1_RS_SFF_9_n6, KE1_RS_SFF_10_n10, KE1_RS_SFF_10_n9,
         KE1_RS_SFF_10_n7, KE1_RS_SFF_10_n6, KE1_RS_SFF_11_n10,
         KE1_RS_SFF_11_n9, KE1_RS_SFF_11_n7, KE1_RS_SFF_11_n6,
         KE1_RS_SFF_12_n10, KE1_RS_SFF_12_n9, KE1_RS_SFF_12_n7,
         KE1_RS_SFF_12_n6, KE1_RS_SFF_13_n11, KE1_RS_SFF_13_n10,
         KE1_RS_SFF_13_n8, KE1_RS_SFF_13_n7, KE1_RS_SFF_14_n11,
         KE1_RS_SFF_14_n10, KE1_RS_SFF_14_n8, KE1_RS_SFF_14_n7,
         KE1_RS_SFF_15_n10, KE1_RS_SFF_15_n9, KE1_RS_SFF_15_n7,
         KE1_RS_SFF_15_n6, KE1_RS_SFF_16_n10, KE1_RS_SFF_16_n9,
         KE1_RS_SFF_16_n7, KE1_RS_SFF_16_n6, KE1_RS_SFF_17_n10,
         KE1_RS_SFF_17_n9, KE1_RS_SFF_17_n7, KE1_RS_SFF_17_n6,
         KE1_RS_SFF_18_n10, KE1_RS_SFF_18_n9, KE1_RS_SFF_18_n7,
         KE1_RS_SFF_18_n6, KE1_RS_SFF_19_n10, KE1_RS_SFF_19_n9,
         KE1_RS_SFF_19_n7, KE1_RS_SFF_19_n6, KE1_RS_SFF_20_n10,
         KE1_RS_SFF_20_n9, KE1_RS_SFF_20_n7, KE1_RS_SFF_20_n6,
         KE1_RS_SFF_21_n10, KE1_RS_SFF_21_n9, KE1_RS_SFF_21_n7,
         KE1_RS_SFF_21_n6, KE1_RS_SFF_22_n10, KE1_RS_SFF_22_n9,
         KE1_RS_SFF_22_n7, KE1_RS_SFF_22_n6, KE1_RS_SFF_23_n10,
         KE1_RS_SFF_23_n9, KE1_RS_SFF_23_n7, KE1_RS_SFF_23_n6,
         KE1_RS_SFF_24_n10, KE1_RS_SFF_24_n9, KE1_RS_SFF_24_n7,
         KE1_RS_SFF_24_n6, KE1_RS_SFF_25_n11, KE1_RS_SFF_25_n10,
         KE1_RS_SFF_25_n8, KE1_RS_SFF_25_n7, KE1_RS_SFF_26_n11,
         KE1_RS_SFF_26_n10, KE1_RS_SFF_26_n8, KE1_RS_SFF_26_n7,
         KE1_RS_SFF_27_n10, KE1_RS_SFF_27_n9, KE1_RS_SFF_27_n7,
         KE1_RS_SFF_27_n6, KE1_RS_SFF_28_n10, KE1_RS_SFF_28_n9,
         KE1_RS_SFF_28_n7, KE1_RS_SFF_28_n6, KE1_RS_SFF_29_n10,
         KE1_RS_SFF_29_n9, KE1_RS_SFF_29_n7, KE1_RS_SFF_29_n6,
         KE1_RS_SFF_30_n10, KE1_RS_SFF_30_n9, KE1_RS_SFF_30_n7,
         KE1_RS_SFF_30_n6, KE1_RS_SFF_31_n10, KE1_RS_SFF_31_n9,
         KE1_RS_SFF_31_n7, KE1_RS_SFF_31_n6, KE1_RS_SFF_32_n10,
         KE1_RS_SFF_32_n9, KE1_RS_SFF_32_n7, KE1_RS_SFF_32_n6,
         KE1_RS_SFF_33_n10, KE1_RS_SFF_33_n9, KE1_RS_SFF_33_n7,
         KE1_RS_SFF_33_n6, KE1_RS_SFF_34_n10, KE1_RS_SFF_34_n9,
         KE1_RS_SFF_34_n7, KE1_RS_SFF_34_n6, KE1_RS_SFF_35_n10,
         KE1_RS_SFF_35_n9, KE1_RS_SFF_35_n7, KE1_RS_SFF_35_n6,
         KE1_RS_SFF_36_n10, KE1_RS_SFF_36_n9, KE1_RS_SFF_36_n7,
         KE1_RS_SFF_36_n6, KE1_RS_SFF_37_n11, KE1_RS_SFF_37_n10,
         KE1_RS_SFF_37_n8, KE1_RS_SFF_37_n7, KE1_RS_SFF_38_n11,
         KE1_RS_SFF_38_n10, KE1_RS_SFF_38_n8, KE1_RS_SFF_38_n7,
         KE1_RS_SFF_39_n10, KE1_RS_SFF_39_n9, KE1_RS_SFF_39_n7,
         KE1_RS_SFF_39_n6, KE1_RS_SFF_40_n10, KE1_RS_SFF_40_n9,
         KE1_RS_SFF_40_n7, KE1_RS_SFF_40_n6, KE1_RS_SFF_41_n10,
         KE1_RS_SFF_41_n9, KE1_RS_SFF_41_n7, KE1_RS_SFF_41_n6,
         KE1_RS_SFF_42_n10, KE1_RS_SFF_42_n9, KE1_RS_SFF_42_n7,
         KE1_RS_SFF_42_n6, KE1_RS_SFF_43_n10, KE1_RS_SFF_43_n9,
         KE1_RS_SFF_43_n7, KE1_RS_SFF_43_n6, KE1_RS_SFF_44_n10,
         KE1_RS_SFF_44_n9, KE1_RS_SFF_44_n7, KE1_RS_SFF_44_n6,
         KE1_RS_SFF_45_n10, KE1_RS_SFF_45_n9, KE1_RS_SFF_45_n7,
         KE1_RS_SFF_45_n6, KE1_RS_SFF_46_n10, KE1_RS_SFF_46_n9,
         KE1_RS_SFF_46_n7, KE1_RS_SFF_46_n6, KE1_RS_SFF_47_n10,
         KE1_RS_SFF_47_n9, KE1_RS_SFF_47_n7, KE1_RS_SFF_47_n6,
         KE1_RS_SFF_48_n10, KE1_RS_SFF_48_n9, KE1_RS_SFF_48_n7,
         KE1_RS_SFF_48_n6, KE1_RS_SFF_49_n11, KE1_RS_SFF_49_n10,
         KE1_RS_SFF_49_n8, KE1_RS_SFF_49_n7, KE1_RS_SFF_50_n11,
         KE1_RS_SFF_50_n10, KE1_RS_SFF_50_n8, KE1_RS_SFF_50_n7,
         KE1_RS_SFF_51_n10, KE1_RS_SFF_51_n9, KE1_RS_SFF_51_n7,
         KE1_RS_SFF_51_n6, KE1_RS_SFF_52_n10, KE1_RS_SFF_52_n9,
         KE1_RS_SFF_52_n7, KE1_RS_SFF_52_n6, KE1_RS_SFF_53_n10,
         KE1_RS_SFF_53_n9, KE1_RS_SFF_53_n7, KE1_RS_SFF_53_n6,
         KE1_RS_SFF_54_n10, KE1_RS_SFF_54_n9, KE1_RS_SFF_54_n7,
         KE1_RS_SFF_54_n6, KE1_RS_SFF_55_n10, KE1_RS_SFF_55_n9,
         KE1_RS_SFF_55_n7, KE1_RS_SFF_55_n6, KE1_RS_SFF_56_n10,
         KE1_RS_SFF_56_n9, KE1_RS_SFF_56_n7, KE1_RS_SFF_56_n6,
         KE1_RS_SFF_57_n10, KE1_RS_SFF_57_n9, KE1_RS_SFF_57_n7,
         KE1_RS_SFF_57_n6, KE1_RS_SFF_58_n10, KE1_RS_SFF_58_n9,
         KE1_RS_SFF_58_n7, KE1_RS_SFF_58_n6, KE1_RS_SFF_59_n10,
         KE1_RS_SFF_59_n9, KE1_RS_SFF_59_n7, KE1_RS_SFF_59_n6,
         KE1_RS_SFF_60_n10, KE1_RS_SFF_60_n9, KE1_RS_SFF_60_n7,
         KE1_RS_SFF_60_n6, KE1_RS_SFF_61_n10, KE1_RS_SFF_61_n9,
         KE1_RS_SFF_61_n7, KE1_RS_SFF_61_n6, KE1_RS_SFF_62_n10,
         KE1_RS_SFF_62_n9, KE1_RS_SFF_62_n7, KE1_RS_SFF_62_n6,
         KE1_RS_SFF_63_n10, KE1_RS_SFF_63_n9, KE1_RS_SFF_63_n7,
         KE1_RS_SFF_63_n6, KE2_RS_n11, KE2_RS_n10, KE2_RS_n9, KE2_RS_n8,
         KE2_RS_n7, KE2_RS_n6, KE2_RS_SFF_0_n11, KE2_RS_SFF_0_n10,
         KE2_RS_SFF_0_n8, KE2_RS_SFF_0_n7, KE2_RS_SFF_1_n11, KE2_RS_SFF_1_n10,
         KE2_RS_SFF_1_n8, KE2_RS_SFF_1_n7, KE2_RS_SFF_2_n10, KE2_RS_SFF_2_n9,
         KE2_RS_SFF_2_n7, KE2_RS_SFF_2_n6, KE2_RS_SFF_3_n10, KE2_RS_SFF_3_n9,
         KE2_RS_SFF_3_n7, KE2_RS_SFF_3_n6, KE2_RS_SFF_4_n10, KE2_RS_SFF_4_n9,
         KE2_RS_SFF_4_n7, KE2_RS_SFF_4_n6, KE2_RS_SFF_5_n10, KE2_RS_SFF_5_n9,
         KE2_RS_SFF_5_n7, KE2_RS_SFF_5_n6, KE2_RS_SFF_6_n10, KE2_RS_SFF_6_n9,
         KE2_RS_SFF_6_n7, KE2_RS_SFF_6_n6, KE2_RS_SFF_7_n10, KE2_RS_SFF_7_n9,
         KE2_RS_SFF_7_n7, KE2_RS_SFF_7_n6, KE2_RS_SFF_8_n10, KE2_RS_SFF_8_n9,
         KE2_RS_SFF_8_n7, KE2_RS_SFF_8_n6, KE2_RS_SFF_9_n10, KE2_RS_SFF_9_n9,
         KE2_RS_SFF_9_n7, KE2_RS_SFF_9_n6, KE2_RS_SFF_10_n10, KE2_RS_SFF_10_n9,
         KE2_RS_SFF_10_n7, KE2_RS_SFF_10_n6, KE2_RS_SFF_11_n10,
         KE2_RS_SFF_11_n9, KE2_RS_SFF_11_n7, KE2_RS_SFF_11_n6,
         KE2_RS_SFF_12_n11, KE2_RS_SFF_12_n10, KE2_RS_SFF_12_n8,
         KE2_RS_SFF_12_n7, KE2_RS_SFF_13_n11, KE2_RS_SFF_13_n10,
         KE2_RS_SFF_13_n8, KE2_RS_SFF_13_n7, KE2_RS_SFF_14_n10,
         KE2_RS_SFF_14_n9, KE2_RS_SFF_14_n7, KE2_RS_SFF_14_n6,
         KE2_RS_SFF_15_n10, KE2_RS_SFF_15_n9, KE2_RS_SFF_15_n7,
         KE2_RS_SFF_15_n6, KE2_RS_SFF_16_n10, KE2_RS_SFF_16_n9,
         KE2_RS_SFF_16_n7, KE2_RS_SFF_16_n6, KE2_RS_SFF_17_n10,
         KE2_RS_SFF_17_n9, KE2_RS_SFF_17_n7, KE2_RS_SFF_17_n6,
         KE2_RS_SFF_18_n10, KE2_RS_SFF_18_n9, KE2_RS_SFF_18_n7,
         KE2_RS_SFF_18_n6, KE2_RS_SFF_19_n10, KE2_RS_SFF_19_n9,
         KE2_RS_SFF_19_n7, KE2_RS_SFF_19_n6, KE2_RS_SFF_20_n10,
         KE2_RS_SFF_20_n9, KE2_RS_SFF_20_n7, KE2_RS_SFF_20_n6,
         KE2_RS_SFF_21_n10, KE2_RS_SFF_21_n9, KE2_RS_SFF_21_n7,
         KE2_RS_SFF_21_n6, KE2_RS_SFF_22_n10, KE2_RS_SFF_22_n9,
         KE2_RS_SFF_22_n7, KE2_RS_SFF_22_n6, KE2_RS_SFF_23_n10,
         KE2_RS_SFF_23_n9, KE2_RS_SFF_23_n7, KE2_RS_SFF_23_n6,
         KE2_RS_SFF_24_n11, KE2_RS_SFF_24_n10, KE2_RS_SFF_24_n8,
         KE2_RS_SFF_24_n7, KE2_RS_SFF_25_n11, KE2_RS_SFF_25_n10,
         KE2_RS_SFF_25_n8, KE2_RS_SFF_25_n7, KE2_RS_SFF_26_n10,
         KE2_RS_SFF_26_n9, KE2_RS_SFF_26_n7, KE2_RS_SFF_26_n6,
         KE2_RS_SFF_27_n10, KE2_RS_SFF_27_n9, KE2_RS_SFF_27_n7,
         KE2_RS_SFF_27_n6, KE2_RS_SFF_28_n10, KE2_RS_SFF_28_n9,
         KE2_RS_SFF_28_n7, KE2_RS_SFF_28_n6, KE2_RS_SFF_29_n10,
         KE2_RS_SFF_29_n9, KE2_RS_SFF_29_n7, KE2_RS_SFF_29_n6,
         KE2_RS_SFF_30_n10, KE2_RS_SFF_30_n9, KE2_RS_SFF_30_n7,
         KE2_RS_SFF_30_n6, KE2_RS_SFF_31_n10, KE2_RS_SFF_31_n9,
         KE2_RS_SFF_31_n7, KE2_RS_SFF_31_n6, KE2_RS_SFF_32_n10,
         KE2_RS_SFF_32_n9, KE2_RS_SFF_32_n7, KE2_RS_SFF_32_n6,
         KE2_RS_SFF_33_n10, KE2_RS_SFF_33_n9, KE2_RS_SFF_33_n7,
         KE2_RS_SFF_33_n6, KE2_RS_SFF_34_n10, KE2_RS_SFF_34_n9,
         KE2_RS_SFF_34_n7, KE2_RS_SFF_34_n6, KE2_RS_SFF_35_n10,
         KE2_RS_SFF_35_n9, KE2_RS_SFF_35_n7, KE2_RS_SFF_35_n6,
         KE2_RS_SFF_36_n11, KE2_RS_SFF_36_n10, KE2_RS_SFF_36_n8,
         KE2_RS_SFF_36_n7, KE2_RS_SFF_37_n11, KE2_RS_SFF_37_n10,
         KE2_RS_SFF_37_n8, KE2_RS_SFF_37_n7, KE2_RS_SFF_38_n10,
         KE2_RS_SFF_38_n9, KE2_RS_SFF_38_n7, KE2_RS_SFF_38_n6,
         KE2_RS_SFF_39_n10, KE2_RS_SFF_39_n9, KE2_RS_SFF_39_n7,
         KE2_RS_SFF_39_n6, KE2_RS_SFF_40_n10, KE2_RS_SFF_40_n9,
         KE2_RS_SFF_40_n7, KE2_RS_SFF_40_n6, KE2_RS_SFF_41_n10,
         KE2_RS_SFF_41_n9, KE2_RS_SFF_41_n7, KE2_RS_SFF_41_n6,
         KE2_RS_SFF_42_n10, KE2_RS_SFF_42_n9, KE2_RS_SFF_42_n7,
         KE2_RS_SFF_42_n6, KE2_RS_SFF_43_n10, KE2_RS_SFF_43_n9,
         KE2_RS_SFF_43_n7, KE2_RS_SFF_43_n6, KE2_RS_SFF_44_n10,
         KE2_RS_SFF_44_n9, KE2_RS_SFF_44_n7, KE2_RS_SFF_44_n6,
         KE2_RS_SFF_45_n10, KE2_RS_SFF_45_n9, KE2_RS_SFF_45_n7,
         KE2_RS_SFF_45_n6, KE2_RS_SFF_46_n10, KE2_RS_SFF_46_n9,
         KE2_RS_SFF_46_n7, KE2_RS_SFF_46_n6, KE2_RS_SFF_47_n10,
         KE2_RS_SFF_47_n9, KE2_RS_SFF_47_n7, KE2_RS_SFF_47_n6,
         KE2_RS_SFF_48_n11, KE2_RS_SFF_48_n10, KE2_RS_SFF_48_n8,
         KE2_RS_SFF_48_n7, KE2_RS_SFF_49_n11, KE2_RS_SFF_49_n10,
         KE2_RS_SFF_49_n8, KE2_RS_SFF_49_n7, KE2_RS_SFF_50_n10,
         KE2_RS_SFF_50_n9, KE2_RS_SFF_50_n7, KE2_RS_SFF_50_n6,
         KE2_RS_SFF_51_n10, KE2_RS_SFF_51_n9, KE2_RS_SFF_51_n7,
         KE2_RS_SFF_51_n6, KE2_RS_SFF_52_n10, KE2_RS_SFF_52_n9,
         KE2_RS_SFF_52_n7, KE2_RS_SFF_52_n6, KE2_RS_SFF_53_n10,
         KE2_RS_SFF_53_n9, KE2_RS_SFF_53_n7, KE2_RS_SFF_53_n6,
         KE2_RS_SFF_54_n10, KE2_RS_SFF_54_n9, KE2_RS_SFF_54_n7,
         KE2_RS_SFF_54_n6, KE2_RS_SFF_55_n10, KE2_RS_SFF_55_n9,
         KE2_RS_SFF_55_n7, KE2_RS_SFF_55_n6, KE2_RS_SFF_56_n10,
         KE2_RS_SFF_56_n9, KE2_RS_SFF_56_n7, KE2_RS_SFF_56_n6,
         KE2_RS_SFF_57_n10, KE2_RS_SFF_57_n9, KE2_RS_SFF_57_n7,
         KE2_RS_SFF_57_n6, KE2_RS_SFF_58_n10, KE2_RS_SFF_58_n9,
         KE2_RS_SFF_58_n7, KE2_RS_SFF_58_n6, KE2_RS_SFF_59_n10,
         KE2_RS_SFF_59_n9, KE2_RS_SFF_59_n7, KE2_RS_SFF_59_n6,
         KE2_RS_SFF_60_n10, KE2_RS_SFF_60_n9, KE2_RS_SFF_60_n7,
         KE2_RS_SFF_60_n6, KE2_RS_SFF_61_n10, KE2_RS_SFF_61_n9,
         KE2_RS_SFF_61_n7, KE2_RS_SFF_61_n6, KE2_RS_SFF_62_n10,
         KE2_RS_SFF_62_n9, KE2_RS_SFF_62_n7, KE2_RS_SFF_62_n6,
         KE2_RS_SFF_63_n10, KE2_RS_SFF_63_n9, KE2_RS_SFF_63_n7,
         KE2_RS_SFF_63_n6, KE3_RS_n12, KE3_RS_n11, KE3_RS_n10, KE3_RS_n9,
         KE3_RS_n8, KE3_RS_n7, KE3_RS_SFF_0_n11, KE3_RS_SFF_0_n10,
         KE3_RS_SFF_0_n8, KE3_RS_SFF_0_n7, KE3_RS_SFF_1_n11, KE3_RS_SFF_1_n10,
         KE3_RS_SFF_1_n8, KE3_RS_SFF_1_n7, KE3_RS_SFF_2_n10, KE3_RS_SFF_2_n9,
         KE3_RS_SFF_2_n7, KE3_RS_SFF_2_n6, KE3_RS_SFF_3_n10, KE3_RS_SFF_3_n9,
         KE3_RS_SFF_3_n7, KE3_RS_SFF_3_n6, KE3_RS_SFF_4_n10, KE3_RS_SFF_4_n9,
         KE3_RS_SFF_4_n7, KE3_RS_SFF_4_n6, KE3_RS_SFF_5_n10, KE3_RS_SFF_5_n9,
         KE3_RS_SFF_5_n7, KE3_RS_SFF_5_n6, KE3_RS_SFF_6_n10, KE3_RS_SFF_6_n9,
         KE3_RS_SFF_6_n7, KE3_RS_SFF_6_n6, KE3_RS_SFF_7_n10, KE3_RS_SFF_7_n9,
         KE3_RS_SFF_7_n7, KE3_RS_SFF_7_n6, KE3_RS_SFF_8_n10, KE3_RS_SFF_8_n9,
         KE3_RS_SFF_8_n7, KE3_RS_SFF_8_n6, KE3_RS_SFF_9_n10, KE3_RS_SFF_9_n9,
         KE3_RS_SFF_9_n7, KE3_RS_SFF_9_n6, KE3_RS_SFF_10_n10, KE3_RS_SFF_10_n9,
         KE3_RS_SFF_10_n7, KE3_RS_SFF_10_n6, KE3_RS_SFF_11_n10,
         KE3_RS_SFF_11_n9, KE3_RS_SFF_11_n7, KE3_RS_SFF_11_n6,
         KE3_RS_SFF_12_n11, KE3_RS_SFF_12_n10, KE3_RS_SFF_12_n8,
         KE3_RS_SFF_12_n7, KE3_RS_SFF_13_n11, KE3_RS_SFF_13_n10,
         KE3_RS_SFF_13_n8, KE3_RS_SFF_13_n7, KE3_RS_SFF_14_n10,
         KE3_RS_SFF_14_n9, KE3_RS_SFF_14_n7, KE3_RS_SFF_14_n6,
         KE3_RS_SFF_15_n10, KE3_RS_SFF_15_n9, KE3_RS_SFF_15_n7,
         KE3_RS_SFF_15_n6, KE3_RS_SFF_16_n10, KE3_RS_SFF_16_n9,
         KE3_RS_SFF_16_n7, KE3_RS_SFF_16_n6, KE3_RS_SFF_17_n10,
         KE3_RS_SFF_17_n9, KE3_RS_SFF_17_n7, KE3_RS_SFF_17_n6,
         KE3_RS_SFF_18_n10, KE3_RS_SFF_18_n9, KE3_RS_SFF_18_n7,
         KE3_RS_SFF_18_n6, KE3_RS_SFF_19_n10, KE3_RS_SFF_19_n9,
         KE3_RS_SFF_19_n7, KE3_RS_SFF_19_n6, KE3_RS_SFF_20_n10,
         KE3_RS_SFF_20_n9, KE3_RS_SFF_20_n7, KE3_RS_SFF_20_n6,
         KE3_RS_SFF_21_n10, KE3_RS_SFF_21_n9, KE3_RS_SFF_21_n7,
         KE3_RS_SFF_21_n6, KE3_RS_SFF_22_n10, KE3_RS_SFF_22_n9,
         KE3_RS_SFF_22_n7, KE3_RS_SFF_22_n6, KE3_RS_SFF_23_n10,
         KE3_RS_SFF_23_n9, KE3_RS_SFF_23_n7, KE3_RS_SFF_23_n6,
         KE3_RS_SFF_24_n11, KE3_RS_SFF_24_n10, KE3_RS_SFF_24_n8,
         KE3_RS_SFF_24_n7, KE3_RS_SFF_25_n11, KE3_RS_SFF_25_n10,
         KE3_RS_SFF_25_n8, KE3_RS_SFF_25_n7, KE3_RS_SFF_26_n10,
         KE3_RS_SFF_26_n9, KE3_RS_SFF_26_n7, KE3_RS_SFF_26_n6,
         KE3_RS_SFF_27_n10, KE3_RS_SFF_27_n9, KE3_RS_SFF_27_n7,
         KE3_RS_SFF_27_n6, KE3_RS_SFF_28_n10, KE3_RS_SFF_28_n9,
         KE3_RS_SFF_28_n7, KE3_RS_SFF_28_n6, KE3_RS_SFF_29_n10,
         KE3_RS_SFF_29_n9, KE3_RS_SFF_29_n7, KE3_RS_SFF_29_n6,
         KE3_RS_SFF_30_n10, KE3_RS_SFF_30_n9, KE3_RS_SFF_30_n7,
         KE3_RS_SFF_30_n6, KE3_RS_SFF_31_n10, KE3_RS_SFF_31_n9,
         KE3_RS_SFF_31_n7, KE3_RS_SFF_31_n6, KE3_RS_SFF_32_n10,
         KE3_RS_SFF_32_n9, KE3_RS_SFF_32_n7, KE3_RS_SFF_32_n6,
         KE3_RS_SFF_33_n10, KE3_RS_SFF_33_n9, KE3_RS_SFF_33_n7,
         KE3_RS_SFF_33_n6, KE3_RS_SFF_34_n10, KE3_RS_SFF_34_n9,
         KE3_RS_SFF_34_n7, KE3_RS_SFF_34_n6, KE3_RS_SFF_35_n10,
         KE3_RS_SFF_35_n9, KE3_RS_SFF_35_n7, KE3_RS_SFF_35_n6,
         KE3_RS_SFF_36_n11, KE3_RS_SFF_36_n10, KE3_RS_SFF_36_n8,
         KE3_RS_SFF_36_n7, KE3_RS_SFF_37_n11, KE3_RS_SFF_37_n10,
         KE3_RS_SFF_37_n8, KE3_RS_SFF_37_n7, KE3_RS_SFF_38_n10,
         KE3_RS_SFF_38_n9, KE3_RS_SFF_38_n7, KE3_RS_SFF_38_n6,
         KE3_RS_SFF_39_n10, KE3_RS_SFF_39_n9, KE3_RS_SFF_39_n7,
         KE3_RS_SFF_39_n6, KE3_RS_SFF_40_n10, KE3_RS_SFF_40_n9,
         KE3_RS_SFF_40_n7, KE3_RS_SFF_40_n6, KE3_RS_SFF_41_n10,
         KE3_RS_SFF_41_n9, KE3_RS_SFF_41_n7, KE3_RS_SFF_41_n6,
         KE3_RS_SFF_42_n10, KE3_RS_SFF_42_n9, KE3_RS_SFF_42_n7,
         KE3_RS_SFF_42_n6, KE3_RS_SFF_43_n10, KE3_RS_SFF_43_n9,
         KE3_RS_SFF_43_n7, KE3_RS_SFF_43_n6, KE3_RS_SFF_44_n10,
         KE3_RS_SFF_44_n9, KE3_RS_SFF_44_n7, KE3_RS_SFF_44_n6,
         KE3_RS_SFF_45_n10, KE3_RS_SFF_45_n9, KE3_RS_SFF_45_n7,
         KE3_RS_SFF_45_n6, KE3_RS_SFF_46_n10, KE3_RS_SFF_46_n9,
         KE3_RS_SFF_46_n7, KE3_RS_SFF_46_n6, KE3_RS_SFF_47_n10,
         KE3_RS_SFF_47_n9, KE3_RS_SFF_47_n7, KE3_RS_SFF_47_n6,
         KE3_RS_SFF_48_n11, KE3_RS_SFF_48_n10, KE3_RS_SFF_48_n8,
         KE3_RS_SFF_48_n7, KE3_RS_SFF_49_n11, KE3_RS_SFF_49_n10,
         KE3_RS_SFF_49_n8, KE3_RS_SFF_49_n7, KE3_RS_SFF_50_n10,
         KE3_RS_SFF_50_n9, KE3_RS_SFF_50_n7, KE3_RS_SFF_50_n6,
         KE3_RS_SFF_51_n10, KE3_RS_SFF_51_n9, KE3_RS_SFF_51_n7,
         KE3_RS_SFF_51_n6, KE3_RS_SFF_52_n10, KE3_RS_SFF_52_n9,
         KE3_RS_SFF_52_n7, KE3_RS_SFF_52_n6, KE3_RS_SFF_53_n10,
         KE3_RS_SFF_53_n9, KE3_RS_SFF_53_n7, KE3_RS_SFF_53_n6,
         KE3_RS_SFF_54_n10, KE3_RS_SFF_54_n9, KE3_RS_SFF_54_n7,
         KE3_RS_SFF_54_n6, KE3_RS_SFF_55_n10, KE3_RS_SFF_55_n9,
         KE3_RS_SFF_55_n7, KE3_RS_SFF_55_n6, KE3_RS_SFF_56_n10,
         KE3_RS_SFF_56_n9, KE3_RS_SFF_56_n7, KE3_RS_SFF_56_n6,
         KE3_RS_SFF_57_n10, KE3_RS_SFF_57_n9, KE3_RS_SFF_57_n7,
         KE3_RS_SFF_57_n6, KE3_RS_SFF_58_n10, KE3_RS_SFF_58_n9,
         KE3_RS_SFF_58_n7, KE3_RS_SFF_58_n6, KE3_RS_SFF_59_n10,
         KE3_RS_SFF_59_n9, KE3_RS_SFF_59_n7, KE3_RS_SFF_59_n6,
         KE3_RS_SFF_60_n10, KE3_RS_SFF_60_n9, KE3_RS_SFF_60_n7,
         KE3_RS_SFF_60_n6, KE3_RS_SFF_61_n10, KE3_RS_SFF_61_n9,
         KE3_RS_SFF_61_n7, KE3_RS_SFF_61_n6, KE3_RS_SFF_62_n10,
         KE3_RS_SFF_62_n9, KE3_RS_SFF_62_n7, KE3_RS_SFF_62_n6,
         KE3_RS_SFF_63_n10, KE3_RS_SFF_63_n9, KE3_RS_SFF_63_n7,
         KE3_RS_SFF_63_n6, CL_n26, CL_n25, CL_n20, CL_n13, CL_n11, CL_n24,
         CL_n23, CL_n22, CL_n21, CL_n3, CL_n2, CL_n1, CL_n19, CL_n18, CL_n17,
         CL_n16, CL_n15, CL_n14, CL_n9, CL_n8, CL_n7, CL_n6, CL_n5, CL_n4,
         CL_N11;
  wire   [5:0] ROUND_CST;
  wire   [63:0] SUB_IN1;
  wire   [63:29] SUB_OUT1;
  wire   [63:29] SUB_OUT2;
  wire   [63:29] SUB_OUT3;
  wire   [47:0] RF1_SHIFTROWS;
  wire   [47:0] RF2_SHIFTROWS;
  wire   [47:0] RF3_SHIFTROWS;
  wire   [3:0] S_0_G_out1;
  wire   [3:0] S_0_F_in3;
  wire   [3:0] S_0_F_in2;
  wire   [3:0] S_0_F_in1;
  wire   [3:0] S_0_q3;
  wire   [3:0] S_0_Rq3;
  wire   [3:0] S_0_q2;
  wire   [3:0] S_0_Rq2;
  wire   [3:0] S_0_q1;
  wire   [3:0] S_0_Rq1;
  wire   [3:2] S_0_F_q3;
  wire   [3:2] S_0_F_q2;
  wire   [3:2] S_0_F_q1;
  wire   [17:0] S_0_F_CF_Reg;
  wire   [17:0] S_0_F_CF_Out;
  wire   [17:0] S_0_G_CF_Reg;
  wire   [17:0] S_0_G_CF_Out;
  wire   [3:0] S_1_G_out1;
  wire   [3:0] S_1_F_in3;
  wire   [3:0] S_1_F_in2;
  wire   [3:0] S_1_F_in1;
  wire   [3:0] S_1_q3;
  wire   [3:0] S_1_Rq3;
  wire   [3:0] S_1_q2;
  wire   [3:0] S_1_Rq2;
  wire   [3:0] S_1_q1;
  wire   [3:0] S_1_Rq1;
  wire   [3:2] S_1_F_q3;
  wire   [3:2] S_1_F_q2;
  wire   [3:2] S_1_F_q1;
  wire   [17:0] S_1_F_CF_Reg;
  wire   [17:0] S_1_F_CF_Out;
  wire   [17:0] S_1_G_CF_Reg;
  wire   [17:0] S_1_G_CF_Out;
  wire   [3:0] S_2_G_out1;
  wire   [3:0] S_2_F_in3;
  wire   [3:0] S_2_F_in2;
  wire   [3:0] S_2_F_in1;
  wire   [3:0] S_2_q3;
  wire   [3:0] S_2_Rq3;
  wire   [3:0] S_2_q2;
  wire   [3:0] S_2_Rq2;
  wire   [3:0] S_2_q1;
  wire   [3:0] S_2_Rq1;
  wire   [3:2] S_2_F_q3;
  wire   [3:2] S_2_F_q2;
  wire   [3:2] S_2_F_q1;
  wire   [17:0] S_2_F_CF_Reg;
  wire   [17:0] S_2_F_CF_Out;
  wire   [17:0] S_2_G_CF_Reg;
  wire   [17:0] S_2_G_CF_Out;
  wire   [3:0] S_3_G_out1;
  wire   [3:0] S_3_F_in3;
  wire   [3:0] S_3_F_in2;
  wire   [3:0] S_3_F_in1;
  wire   [3:0] S_3_q3;
  wire   [3:0] S_3_Rq3;
  wire   [3:0] S_3_q2;
  wire   [3:0] S_3_Rq2;
  wire   [3:0] S_3_q1;
  wire   [3:0] S_3_Rq1;
  wire   [3:2] S_3_F_q3;
  wire   [3:2] S_3_F_q2;
  wire   [3:2] S_3_F_q1;
  wire   [17:0] S_3_F_CF_Reg;
  wire   [17:0] S_3_F_CF_Out;
  wire   [17:0] S_3_G_CF_Reg;
  wire   [17:0] S_3_G_CF_Out;
  wire   [3:0] S_4_G_out1;
  wire   [3:0] S_4_F_in3;
  wire   [3:0] S_4_F_in2;
  wire   [3:0] S_4_F_in1;
  wire   [3:0] S_4_q3;
  wire   [3:0] S_4_Rq3;
  wire   [3:0] S_4_q2;
  wire   [3:0] S_4_Rq2;
  wire   [3:0] S_4_q1;
  wire   [3:0] S_4_Rq1;
  wire   [3:2] S_4_F_q3;
  wire   [3:2] S_4_F_q2;
  wire   [3:2] S_4_F_q1;
  wire   [17:0] S_4_F_CF_Reg;
  wire   [17:0] S_4_F_CF_Out;
  wire   [17:0] S_4_G_CF_Reg;
  wire   [17:0] S_4_G_CF_Out;
  wire   [3:0] S_5_G_out1;
  wire   [3:0] S_5_F_in3;
  wire   [3:0] S_5_F_in2;
  wire   [3:0] S_5_F_in1;
  wire   [3:0] S_5_q3;
  wire   [3:0] S_5_Rq3;
  wire   [3:0] S_5_q2;
  wire   [3:0] S_5_Rq2;
  wire   [3:0] S_5_q1;
  wire   [3:0] S_5_Rq1;
  wire   [3:2] S_5_F_q3;
  wire   [3:2] S_5_F_q2;
  wire   [3:2] S_5_F_q1;
  wire   [17:0] S_5_F_CF_Reg;
  wire   [17:0] S_5_F_CF_Out;
  wire   [17:0] S_5_G_CF_Reg;
  wire   [17:0] S_5_G_CF_Out;
  wire   [3:0] S_6_G_out1;
  wire   [3:0] S_6_F_in3;
  wire   [3:0] S_6_F_in2;
  wire   [3:0] S_6_F_in1;
  wire   [3:0] S_6_q3;
  wire   [3:0] S_6_Rq3;
  wire   [3:0] S_6_q2;
  wire   [3:0] S_6_Rq2;
  wire   [3:0] S_6_q1;
  wire   [3:0] S_6_Rq1;
  wire   [3:2] S_6_F_q3;
  wire   [3:2] S_6_F_q2;
  wire   [3:2] S_6_F_q1;
  wire   [17:0] S_6_F_CF_Reg;
  wire   [17:0] S_6_F_CF_Out;
  wire   [17:0] S_6_G_CF_Reg;
  wire   [17:0] S_6_G_CF_Out;
  wire   [3:0] S_7_G_out1;
  wire   [3:0] S_7_F_in3;
  wire   [3:0] S_7_F_in2;
  wire   [3:0] S_7_F_in1;
  wire   [3:0] S_7_q3;
  wire   [3:0] S_7_Rq3;
  wire   [3:0] S_7_q2;
  wire   [3:0] S_7_Rq2;
  wire   [3:0] S_7_q1;
  wire   [3:0] S_7_Rq1;
  wire   [3:2] S_7_F_q3;
  wire   [3:2] S_7_F_q2;
  wire   [3:2] S_7_F_q1;
  wire   [17:0] S_7_F_CF_Reg;
  wire   [17:0] S_7_F_CF_Out;
  wire   [17:0] S_7_G_CF_Reg;
  wire   [17:0] S_7_G_CF_Out;
  wire   [3:0] S_8_G_out1;
  wire   [3:0] S_8_F_in3;
  wire   [3:0] S_8_F_in2;
  wire   [3:0] S_8_F_in1;
  wire   [3:0] S_8_q3;
  wire   [3:0] S_8_Rq3;
  wire   [3:0] S_8_q2;
  wire   [3:0] S_8_Rq2;
  wire   [3:0] S_8_q1;
  wire   [3:0] S_8_Rq1;
  wire   [3:2] S_8_F_q3;
  wire   [3:2] S_8_F_q2;
  wire   [3:2] S_8_F_q1;
  wire   [17:0] S_8_F_CF_Reg;
  wire   [17:0] S_8_F_CF_Out;
  wire   [17:0] S_8_G_CF_Reg;
  wire   [17:0] S_8_G_CF_Out;
  wire   [3:0] S_9_G_out1;
  wire   [3:0] S_9_F_in3;
  wire   [3:0] S_9_F_in2;
  wire   [3:0] S_9_F_in1;
  wire   [3:0] S_9_q3;
  wire   [3:0] S_9_Rq3;
  wire   [3:0] S_9_q2;
  wire   [3:0] S_9_Rq2;
  wire   [3:0] S_9_q1;
  wire   [3:0] S_9_Rq1;
  wire   [3:2] S_9_F_q3;
  wire   [3:2] S_9_F_q2;
  wire   [3:2] S_9_F_q1;
  wire   [17:0] S_9_F_CF_Reg;
  wire   [17:0] S_9_F_CF_Out;
  wire   [17:0] S_9_G_CF_Reg;
  wire   [17:0] S_9_G_CF_Out;
  wire   [3:0] S_10_G_out1;
  wire   [3:0] S_10_F_in3;
  wire   [3:0] S_10_F_in2;
  wire   [3:0] S_10_F_in1;
  wire   [3:0] S_10_q3;
  wire   [3:0] S_10_Rq3;
  wire   [3:0] S_10_q2;
  wire   [3:0] S_10_Rq2;
  wire   [3:0] S_10_q1;
  wire   [3:0] S_10_Rq1;
  wire   [3:2] S_10_F_q3;
  wire   [3:2] S_10_F_q2;
  wire   [3:2] S_10_F_q1;
  wire   [17:0] S_10_F_CF_Reg;
  wire   [17:0] S_10_F_CF_Out;
  wire   [17:0] S_10_G_CF_Reg;
  wire   [17:0] S_10_G_CF_Out;
  wire   [3:0] S_11_G_out1;
  wire   [3:0] S_11_F_in3;
  wire   [3:0] S_11_F_in2;
  wire   [3:0] S_11_F_in1;
  wire   [3:0] S_11_q3;
  wire   [3:0] S_11_Rq3;
  wire   [3:0] S_11_q2;
  wire   [3:0] S_11_Rq2;
  wire   [3:0] S_11_q1;
  wire   [3:0] S_11_Rq1;
  wire   [3:2] S_11_F_q3;
  wire   [3:2] S_11_F_q2;
  wire   [3:2] S_11_F_q1;
  wire   [17:0] S_11_F_CF_Reg;
  wire   [17:0] S_11_F_CF_Out;
  wire   [17:0] S_11_G_CF_Reg;
  wire   [17:0] S_11_G_CF_Out;
  wire   [3:0] S_12_G_out1;
  wire   [3:0] S_12_F_in3;
  wire   [3:0] S_12_F_in2;
  wire   [3:0] S_12_F_in1;
  wire   [3:0] S_12_q3;
  wire   [3:0] S_12_Rq3;
  wire   [3:0] S_12_q2;
  wire   [3:0] S_12_Rq2;
  wire   [3:0] S_12_q1;
  wire   [3:0] S_12_Rq1;
  wire   [3:2] S_12_F_q3;
  wire   [3:2] S_12_F_q2;
  wire   [3:2] S_12_F_q1;
  wire   [17:0] S_12_F_CF_Reg;
  wire   [17:0] S_12_F_CF_Out;
  wire   [17:0] S_12_G_CF_Reg;
  wire   [17:0] S_12_G_CF_Out;
  wire   [3:0] S_13_G_out1;
  wire   [3:0] S_13_F_in3;
  wire   [3:0] S_13_F_in2;
  wire   [3:0] S_13_F_in1;
  wire   [3:0] S_13_q3;
  wire   [3:0] S_13_Rq3;
  wire   [3:0] S_13_q2;
  wire   [3:0] S_13_Rq2;
  wire   [3:0] S_13_q1;
  wire   [3:0] S_13_Rq1;
  wire   [3:2] S_13_F_q3;
  wire   [3:2] S_13_F_q2;
  wire   [3:2] S_13_F_q1;
  wire   [17:0] S_13_F_CF_Reg;
  wire   [17:0] S_13_F_CF_Out;
  wire   [17:0] S_13_G_CF_Reg;
  wire   [17:0] S_13_G_CF_Out;
  wire   [3:0] S_14_G_out1;
  wire   [3:0] S_14_F_in3;
  wire   [3:0] S_14_F_in2;
  wire   [3:0] S_14_F_in1;
  wire   [3:0] S_14_q3;
  wire   [3:0] S_14_Rq3;
  wire   [3:0] S_14_q2;
  wire   [3:0] S_14_Rq2;
  wire   [3:0] S_14_q1;
  wire   [3:0] S_14_Rq1;
  wire   [3:2] S_14_F_q3;
  wire   [3:2] S_14_F_q2;
  wire   [3:2] S_14_F_q1;
  wire   [17:0] S_14_F_CF_Reg;
  wire   [17:0] S_14_F_CF_Out;
  wire   [17:0] S_14_G_CF_Reg;
  wire   [17:0] S_14_G_CF_Out;
  wire   [3:0] S_15_G_out1;
  wire   [3:0] S_15_F_in3;
  wire   [3:0] S_15_F_in2;
  wire   [3:0] S_15_F_in1;
  wire   [3:0] S_15_q3;
  wire   [3:0] S_15_Rq3;
  wire   [3:0] S_15_q2;
  wire   [3:0] S_15_Rq2;
  wire   [3:0] S_15_q1;
  wire   [3:0] S_15_Rq1;
  wire   [3:2] S_15_F_q3;
  wire   [3:2] S_15_F_q2;
  wire   [3:2] S_15_F_q1;
  wire   [17:0] S_15_F_CF_Reg;
  wire   [17:0] S_15_F_CF_Out;
  wire   [17:0] S_15_G_CF_Reg;
  wire   [17:0] S_15_G_CF_Out;
  wire   [63:0] KE1_KEY_PERM;
  wire   [63:0] KE2_KEY_PERM;
  wire   [63:0] KE3_KEY_PERM;

  SDFF_X1 RF1_RS_SFF_0_Q_reg ( .D(CIPHERTEXT1[0]), .SI(PLAINTEXT1[0]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[0]), .QN() );
  SDFF_X1 RF1_RS_SFF_1_Q_reg ( .D(CIPHERTEXT1[1]), .SI(PLAINTEXT1[1]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[1]), .QN() );
  SDFF_X1 RF1_RS_SFF_2_Q_reg ( .D(CIPHERTEXT1[2]), .SI(PLAINTEXT1[2]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[2]), .QN() );
  SDFF_X1 RF1_RS_SFF_3_Q_reg ( .D(CIPHERTEXT1[3]), .SI(PLAINTEXT1[3]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[3]), .QN() );
  SDFF_X1 RF1_RS_SFF_4_Q_reg ( .D(CIPHERTEXT1[4]), .SI(PLAINTEXT1[4]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[4]), .QN() );
  SDFF_X1 RF1_RS_SFF_5_Q_reg ( .D(CIPHERTEXT1[5]), .SI(PLAINTEXT1[5]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[5]), .QN() );
  SDFF_X1 RF1_RS_SFF_6_Q_reg ( .D(CIPHERTEXT1[6]), .SI(PLAINTEXT1[6]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[6]), .QN() );
  SDFF_X1 RF1_RS_SFF_7_Q_reg ( .D(CIPHERTEXT1[7]), .SI(PLAINTEXT1[7]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[7]), .QN() );
  SDFF_X1 RF1_RS_SFF_8_Q_reg ( .D(CIPHERTEXT1[8]), .SI(PLAINTEXT1[8]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[8]), .QN() );
  SDFF_X1 RF1_RS_SFF_9_Q_reg ( .D(CIPHERTEXT1[9]), .SI(PLAINTEXT1[9]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[9]), .QN() );
  SDFF_X1 RF1_RS_SFF_10_Q_reg ( .D(CIPHERTEXT1[10]), .SI(PLAINTEXT1[10]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[10]), .QN() );
  SDFF_X1 RF1_RS_SFF_11_Q_reg ( .D(CIPHERTEXT1[11]), .SI(PLAINTEXT1[11]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[11]), .QN() );
  SDFF_X1 RF1_RS_SFF_12_Q_reg ( .D(CIPHERTEXT1[12]), .SI(PLAINTEXT1[12]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[12]), .QN() );
  SDFF_X1 RF1_RS_SFF_13_Q_reg ( .D(CIPHERTEXT1[13]), .SI(PLAINTEXT1[13]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[13]), .QN() );
  SDFF_X1 RF1_RS_SFF_14_Q_reg ( .D(CIPHERTEXT1[14]), .SI(PLAINTEXT1[14]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[14]), .QN() );
  SDFF_X1 RF1_RS_SFF_15_Q_reg ( .D(CIPHERTEXT1[15]), .SI(PLAINTEXT1[15]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[15]), .QN() );
  SDFF_X1 RF1_RS_SFF_16_Q_reg ( .D(CIPHERTEXT1[16]), .SI(PLAINTEXT1[16]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[16]), .QN() );
  SDFF_X1 RF1_RS_SFF_17_Q_reg ( .D(CIPHERTEXT1[17]), .SI(PLAINTEXT1[17]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[17]), .QN() );
  SDFF_X1 RF1_RS_SFF_18_Q_reg ( .D(CIPHERTEXT1[18]), .SI(PLAINTEXT1[18]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[18]), .QN() );
  SDFF_X1 RF1_RS_SFF_19_Q_reg ( .D(CIPHERTEXT1[19]), .SI(PLAINTEXT1[19]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[19]), .QN() );
  SDFF_X1 RF1_RS_SFF_20_Q_reg ( .D(CIPHERTEXT1[20]), .SI(PLAINTEXT1[20]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[20]), .QN() );
  SDFF_X1 RF1_RS_SFF_21_Q_reg ( .D(CIPHERTEXT1[21]), .SI(PLAINTEXT1[21]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[21]), .QN() );
  SDFF_X1 RF1_RS_SFF_22_Q_reg ( .D(CIPHERTEXT1[22]), .SI(PLAINTEXT1[22]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[22]), .QN() );
  SDFF_X1 RF1_RS_SFF_23_Q_reg ( .D(CIPHERTEXT1[23]), .SI(PLAINTEXT1[23]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[23]), .QN() );
  SDFF_X1 RF1_RS_SFF_24_Q_reg ( .D(CIPHERTEXT1[24]), .SI(PLAINTEXT1[24]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[24]), .QN() );
  SDFF_X1 RF1_RS_SFF_25_Q_reg ( .D(CIPHERTEXT1[25]), .SI(PLAINTEXT1[25]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[25]), .QN() );
  SDFF_X1 RF1_RS_SFF_26_Q_reg ( .D(CIPHERTEXT1[26]), .SI(PLAINTEXT1[26]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[26]), .QN() );
  SDFF_X1 RF1_RS_SFF_27_Q_reg ( .D(CIPHERTEXT1[27]), .SI(PLAINTEXT1[27]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[27]), .QN() );
  SDFF_X1 RF1_RS_SFF_28_Q_reg ( .D(CIPHERTEXT1[28]), .SI(PLAINTEXT1[28]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[28]), .QN() );
  SDFF_X1 RF1_RS_SFF_29_Q_reg ( .D(CIPHERTEXT1[29]), .SI(PLAINTEXT1[29]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[29]), .QN() );
  SDFF_X1 RF1_RS_SFF_30_Q_reg ( .D(CIPHERTEXT1[30]), .SI(PLAINTEXT1[30]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[30]), .QN() );
  SDFF_X1 RF1_RS_SFF_31_Q_reg ( .D(CIPHERTEXT1[31]), .SI(PLAINTEXT1[31]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[31]), .QN() );
  SDFF_X1 RF1_RS_SFF_32_Q_reg ( .D(CIPHERTEXT1[32]), .SI(PLAINTEXT1[32]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[32]), .QN() );
  SDFF_X1 RF1_RS_SFF_33_Q_reg ( .D(CIPHERTEXT1[33]), .SI(PLAINTEXT1[33]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[33]), .QN() );
  SDFF_X1 RF1_RS_SFF_34_Q_reg ( .D(CIPHERTEXT1[34]), .SI(PLAINTEXT1[34]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[34]), .QN() );
  SDFF_X1 RF1_RS_SFF_35_Q_reg ( .D(CIPHERTEXT1[35]), .SI(PLAINTEXT1[35]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[35]), .QN() );
  SDFF_X1 RF1_RS_SFF_36_Q_reg ( .D(CIPHERTEXT1[36]), .SI(PLAINTEXT1[36]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[36]), .QN() );
  SDFF_X1 RF1_RS_SFF_37_Q_reg ( .D(CIPHERTEXT1[37]), .SI(PLAINTEXT1[37]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[37]), .QN() );
  SDFF_X1 RF1_RS_SFF_38_Q_reg ( .D(CIPHERTEXT1[38]), .SI(PLAINTEXT1[38]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[38]), .QN() );
  SDFF_X1 RF1_RS_SFF_39_Q_reg ( .D(CIPHERTEXT1[39]), .SI(PLAINTEXT1[39]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[39]), .QN() );
  SDFF_X1 RF1_RS_SFF_40_Q_reg ( .D(CIPHERTEXT1[40]), .SI(PLAINTEXT1[40]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[40]), .QN() );
  SDFF_X1 RF1_RS_SFF_41_Q_reg ( .D(CIPHERTEXT1[41]), .SI(PLAINTEXT1[41]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[41]), .QN() );
  SDFF_X1 RF1_RS_SFF_42_Q_reg ( .D(CIPHERTEXT1[42]), .SI(PLAINTEXT1[42]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[42]), .QN() );
  SDFF_X1 RF1_RS_SFF_43_Q_reg ( .D(CIPHERTEXT1[43]), .SI(PLAINTEXT1[43]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[43]), .QN() );
  SDFF_X1 RF1_RS_SFF_44_Q_reg ( .D(CIPHERTEXT1[44]), .SI(PLAINTEXT1[44]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[44]), .QN() );
  SDFF_X1 RF1_RS_SFF_45_Q_reg ( .D(CIPHERTEXT1[45]), .SI(PLAINTEXT1[45]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[45]), .QN() );
  SDFF_X1 RF1_RS_SFF_46_Q_reg ( .D(CIPHERTEXT1[46]), .SI(PLAINTEXT1[46]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[46]), .QN() );
  SDFF_X1 RF1_RS_SFF_47_Q_reg ( .D(CIPHERTEXT1[47]), .SI(PLAINTEXT1[47]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[47]), .QN() );
  SDFF_X1 RF1_RS_SFF_48_Q_reg ( .D(CIPHERTEXT1[48]), .SI(PLAINTEXT1[48]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[48]), .QN() );
  SDFF_X1 RF1_RS_SFF_49_Q_reg ( .D(CIPHERTEXT1[49]), .SI(PLAINTEXT1[49]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[49]), .QN() );
  SDFF_X1 RF1_RS_SFF_50_Q_reg ( .D(CIPHERTEXT1[50]), .SI(PLAINTEXT1[50]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[50]), .QN() );
  SDFF_X1 RF1_RS_SFF_51_Q_reg ( .D(CIPHERTEXT1[51]), .SI(PLAINTEXT1[51]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[51]), .QN() );
  SDFF_X1 RF1_RS_SFF_52_Q_reg ( .D(CIPHERTEXT1[52]), .SI(PLAINTEXT1[52]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[52]), .QN() );
  SDFF_X1 RF1_RS_SFF_53_Q_reg ( .D(CIPHERTEXT1[53]), .SI(PLAINTEXT1[53]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[53]), .QN() );
  SDFF_X1 RF1_RS_SFF_54_Q_reg ( .D(CIPHERTEXT1[54]), .SI(PLAINTEXT1[54]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[54]), .QN() );
  SDFF_X1 RF1_RS_SFF_55_Q_reg ( .D(CIPHERTEXT1[55]), .SI(PLAINTEXT1[55]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[55]), .QN() );
  SDFF_X1 RF1_RS_SFF_56_Q_reg ( .D(CIPHERTEXT1[56]), .SI(PLAINTEXT1[56]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[56]), .QN() );
  SDFF_X1 RF1_RS_SFF_57_Q_reg ( .D(CIPHERTEXT1[57]), .SI(PLAINTEXT1[57]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[57]), .QN() );
  SDFF_X1 RF1_RS_SFF_58_Q_reg ( .D(CIPHERTEXT1[58]), .SI(PLAINTEXT1[58]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[58]), .QN() );
  SDFF_X1 RF1_RS_SFF_59_Q_reg ( .D(CIPHERTEXT1[59]), .SI(PLAINTEXT1[59]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[59]), .QN() );
  SDFF_X1 RF1_RS_SFF_60_Q_reg ( .D(CIPHERTEXT1[60]), .SI(PLAINTEXT1[60]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[60]), .QN() );
  SDFF_X1 RF1_RS_SFF_61_Q_reg ( .D(CIPHERTEXT1[61]), .SI(PLAINTEXT1[61]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[61]), .QN() );
  SDFF_X1 RF1_RS_SFF_62_Q_reg ( .D(CIPHERTEXT1[62]), .SI(PLAINTEXT1[62]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[62]), .QN() );
  SDFF_X1 RF1_RS_SFF_63_Q_reg ( .D(CIPHERTEXT1[63]), .SI(PLAINTEXT1[63]), .SE(
        RESET), .CK(CLK), .Q(SUB_IN1[63]), .QN() );
  INV_X1 RF1_KA_U39 ( .A(SUB_OUT1[29]), .ZN(RF1_SHIFTROWS[21]) );
  XNOR2_X1 RF1_KA_U38 ( .A(RF1_KA_n18), .B(KE1_KEY_PERM[31]), .ZN(
        CIPHERTEXT1[47]) );
  XNOR2_X1 RF1_KA_U37 ( .A(ROUND_CST[3]), .B(SUB_OUT1[63]), .ZN(RF1_KA_n18) );
  XNOR2_X1 RF1_KA_U36 ( .A(RF1_KA_n17), .B(KE1_KEY_PERM[30]), .ZN(
        CIPHERTEXT1[46]) );
  XNOR2_X1 RF1_KA_U35 ( .A(ROUND_CST[2]), .B(SUB_OUT1[62]), .ZN(RF1_KA_n17) );
  XNOR2_X1 RF1_KA_U34 ( .A(RF1_KA_n16), .B(KE1_KEY_PERM[29]), .ZN(
        CIPHERTEXT1[45]) );
  XNOR2_X1 RF1_KA_U33 ( .A(ROUND_CST[1]), .B(SUB_OUT1[61]), .ZN(RF1_KA_n16) );
  XNOR2_X1 RF1_KA_U32 ( .A(RF1_KA_n15), .B(KE1_KEY_PERM[28]), .ZN(
        CIPHERTEXT1[44]) );
  XNOR2_X1 RF1_KA_U31 ( .A(ROUND_CST[0]), .B(SUB_OUT1[60]), .ZN(RF1_KA_n15) );
  XOR2_X1 RF1_KA_U30 ( .A(SUB_OUT1[59]), .B(KE1_KEY_PERM[27]), .Z(
        CIPHERTEXT1[43]) );
  XOR2_X1 RF1_KA_U29 ( .A(SUB_OUT1[58]), .B(KE1_KEY_PERM[26]), .Z(
        CIPHERTEXT1[42]) );
  XOR2_X1 RF1_KA_U28 ( .A(SUB_OUT1[57]), .B(KE1_KEY_PERM[25]), .Z(
        CIPHERTEXT1[41]) );
  XOR2_X1 RF1_KA_U27 ( .A(SUB_OUT1[56]), .B(KE1_KEY_PERM[24]), .Z(
        CIPHERTEXT1[40]) );
  XOR2_X1 RF1_KA_U26 ( .A(SUB_OUT1[55]), .B(KE1_KEY_PERM[23]), .Z(
        CIPHERTEXT1[39]) );
  XOR2_X1 RF1_KA_U25 ( .A(SUB_OUT1[54]), .B(KE1_KEY_PERM[22]), .Z(
        CIPHERTEXT1[38]) );
  XOR2_X1 RF1_KA_U24 ( .A(SUB_OUT1[53]), .B(KE1_KEY_PERM[21]), .Z(
        CIPHERTEXT1[37]) );
  XOR2_X1 RF1_KA_U23 ( .A(SUB_OUT1[52]), .B(KE1_KEY_PERM[20]), .Z(
        CIPHERTEXT1[36]) );
  XOR2_X1 RF1_KA_U22 ( .A(SUB_OUT1[51]), .B(KE1_KEY_PERM[19]), .Z(
        CIPHERTEXT1[35]) );
  XOR2_X1 RF1_KA_U21 ( .A(SUB_OUT1[50]), .B(KE1_KEY_PERM[18]), .Z(
        CIPHERTEXT1[34]) );
  XOR2_X1 RF1_KA_U20 ( .A(SUB_OUT1[49]), .B(KE1_KEY_PERM[17]), .Z(
        CIPHERTEXT1[33]) );
  XOR2_X1 RF1_KA_U19 ( .A(SUB_OUT1[48]), .B(KE1_KEY_PERM[16]), .Z(
        CIPHERTEXT1[32]) );
  XOR2_X1 RF1_KA_U18 ( .A(SUB_OUT1[47]), .B(KE1_KEY_PERM[15]), .Z(
        RF1_SHIFTROWS[43]) );
  XOR2_X1 RF1_KA_U17 ( .A(SUB_OUT1[46]), .B(KE1_KEY_PERM[14]), .Z(
        RF1_SHIFTROWS[42]) );
  XNOR2_X1 RF1_KA_U16 ( .A(RF1_KA_n14), .B(KE1_KEY_PERM[13]), .ZN(
        RF1_SHIFTROWS[41]) );
  XNOR2_X1 RF1_KA_U15 ( .A(ROUND_CST[5]), .B(SUB_OUT1[45]), .ZN(RF1_KA_n14) );
  XNOR2_X1 RF1_KA_U14 ( .A(RF1_KA_n13), .B(KE1_KEY_PERM[12]), .ZN(
        RF1_SHIFTROWS[40]) );
  XNOR2_X1 RF1_KA_U13 ( .A(ROUND_CST[4]), .B(SUB_OUT1[44]), .ZN(RF1_KA_n13) );
  XOR2_X1 RF1_KA_U12 ( .A(SUB_OUT1[43]), .B(KE1_KEY_PERM[11]), .Z(
        RF1_SHIFTROWS[39]) );
  XOR2_X1 RF1_KA_U11 ( .A(SUB_OUT1[42]), .B(KE1_KEY_PERM[10]), .Z(
        RF1_SHIFTROWS[38]) );
  XOR2_X1 RF1_KA_U10 ( .A(SUB_OUT1[41]), .B(KE1_KEY_PERM[9]), .Z(
        RF1_SHIFTROWS[37]) );
  XOR2_X1 RF1_KA_U9 ( .A(SUB_OUT1[40]), .B(KE1_KEY_PERM[8]), .Z(
        RF1_SHIFTROWS[36]) );
  XOR2_X1 RF1_KA_U8 ( .A(SUB_OUT1[39]), .B(KE1_KEY_PERM[7]), .Z(
        RF1_SHIFTROWS[35]) );
  XOR2_X1 RF1_KA_U7 ( .A(SUB_OUT1[38]), .B(KE1_KEY_PERM[6]), .Z(
        RF1_SHIFTROWS[34]) );
  XOR2_X1 RF1_KA_U6 ( .A(SUB_OUT1[37]), .B(KE1_KEY_PERM[5]), .Z(
        RF1_SHIFTROWS[33]) );
  XOR2_X1 RF1_KA_U5 ( .A(SUB_OUT1[36]), .B(KE1_KEY_PERM[4]), .Z(
        RF1_SHIFTROWS[32]) );
  XOR2_X1 RF1_KA_U4 ( .A(SUB_OUT1[35]), .B(KE1_KEY_PERM[3]), .Z(
        RF1_SHIFTROWS[47]) );
  XOR2_X1 RF1_KA_U3 ( .A(SUB_OUT1[34]), .B(KE1_KEY_PERM[2]), .Z(
        RF1_SHIFTROWS[46]) );
  XOR2_X1 RF1_KA_U2 ( .A(SUB_OUT1[33]), .B(KE1_KEY_PERM[1]), .Z(
        RF1_SHIFTROWS[45]) );
  XOR2_X1 RF1_KA_U1 ( .A(SUB_OUT1[32]), .B(KE1_KEY_PERM[0]), .Z(
        RF1_SHIFTROWS[44]) );
  XOR2_X1 RF1_MC_U48 ( .A(RF1_SHIFTROWS[15]), .B(CIPHERTEXT1[15]), .Z(
        CIPHERTEXT1[63]) );
  XOR2_X1 RF1_MC_U47 ( .A(RF1_SHIFTROWS[14]), .B(CIPHERTEXT1[14]), .Z(
        CIPHERTEXT1[62]) );
  XOR2_X1 RF1_MC_U46 ( .A(RF1_SHIFTROWS[13]), .B(CIPHERTEXT1[13]), .Z(
        CIPHERTEXT1[61]) );
  XOR2_X1 RF1_MC_U45 ( .A(RF1_SHIFTROWS[12]), .B(CIPHERTEXT1[12]), .Z(
        CIPHERTEXT1[60]) );
  XOR2_X1 RF1_MC_U44 ( .A(RF1_SHIFTROWS[11]), .B(CIPHERTEXT1[11]), .Z(
        CIPHERTEXT1[59]) );
  XOR2_X1 RF1_MC_U43 ( .A(RF1_SHIFTROWS[10]), .B(CIPHERTEXT1[10]), .Z(
        CIPHERTEXT1[58]) );
  XOR2_X1 RF1_MC_U42 ( .A(RF1_SHIFTROWS[9]), .B(CIPHERTEXT1[9]), .Z(
        CIPHERTEXT1[57]) );
  XOR2_X1 RF1_MC_U41 ( .A(CIPHERTEXT1[41]), .B(RF1_SHIFTROWS[25]), .Z(
        CIPHERTEXT1[9]) );
  XOR2_X1 RF1_MC_U40 ( .A(RF1_SHIFTROWS[8]), .B(CIPHERTEXT1[8]), .Z(
        CIPHERTEXT1[56]) );
  XOR2_X1 RF1_MC_U39 ( .A(CIPHERTEXT1[40]), .B(RF1_SHIFTROWS[24]), .Z(
        CIPHERTEXT1[8]) );
  XOR2_X1 RF1_MC_U38 ( .A(RF1_SHIFTROWS[7]), .B(CIPHERTEXT1[7]), .Z(
        CIPHERTEXT1[55]) );
  XOR2_X1 RF1_MC_U37 ( .A(CIPHERTEXT1[39]), .B(RF1_SHIFTROWS[23]), .Z(
        CIPHERTEXT1[7]) );
  XOR2_X1 RF1_MC_U36 ( .A(RF1_SHIFTROWS[6]), .B(CIPHERTEXT1[6]), .Z(
        CIPHERTEXT1[54]) );
  XOR2_X1 RF1_MC_U35 ( .A(CIPHERTEXT1[38]), .B(RF1_SHIFTROWS[22]), .Z(
        CIPHERTEXT1[6]) );
  XOR2_X1 RF1_MC_U34 ( .A(RF1_SHIFTROWS[5]), .B(CIPHERTEXT1[5]), .Z(
        CIPHERTEXT1[53]) );
  XOR2_X1 RF1_MC_U33 ( .A(CIPHERTEXT1[37]), .B(RF1_SHIFTROWS[21]), .Z(
        CIPHERTEXT1[5]) );
  XOR2_X1 RF1_MC_U32 ( .A(RF1_SHIFTROWS[4]), .B(CIPHERTEXT1[4]), .Z(
        CIPHERTEXT1[52]) );
  XOR2_X1 RF1_MC_U31 ( .A(RF1_SHIFTROWS[3]), .B(CIPHERTEXT1[3]), .Z(
        CIPHERTEXT1[51]) );
  XOR2_X1 RF1_MC_U30 ( .A(RF1_SHIFTROWS[2]), .B(CIPHERTEXT1[2]), .Z(
        CIPHERTEXT1[50]) );
  XOR2_X1 RF1_MC_U29 ( .A(CIPHERTEXT1[36]), .B(RF1_SHIFTROWS[20]), .Z(
        CIPHERTEXT1[4]) );
  XOR2_X1 RF1_MC_U28 ( .A(RF1_SHIFTROWS[1]), .B(CIPHERTEXT1[1]), .Z(
        CIPHERTEXT1[49]) );
  XOR2_X1 RF1_MC_U27 ( .A(RF1_SHIFTROWS[0]), .B(CIPHERTEXT1[0]), .Z(
        CIPHERTEXT1[48]) );
  XOR2_X1 RF1_MC_U26 ( .A(CIPHERTEXT1[35]), .B(RF1_SHIFTROWS[19]), .Z(
        CIPHERTEXT1[3]) );
  XOR2_X1 RF1_MC_U25 ( .A(RF1_SHIFTROWS[31]), .B(RF1_SHIFTROWS[47]), .Z(
        CIPHERTEXT1[31]) );
  XOR2_X1 RF1_MC_U24 ( .A(RF1_SHIFTROWS[30]), .B(RF1_SHIFTROWS[46]), .Z(
        CIPHERTEXT1[30]) );
  XOR2_X1 RF1_MC_U23 ( .A(CIPHERTEXT1[34]), .B(RF1_SHIFTROWS[18]), .Z(
        CIPHERTEXT1[2]) );
  XOR2_X1 RF1_MC_U22 ( .A(RF1_SHIFTROWS[29]), .B(RF1_SHIFTROWS[45]), .Z(
        CIPHERTEXT1[29]) );
  XOR2_X1 RF1_MC_U21 ( .A(RF1_SHIFTROWS[28]), .B(RF1_SHIFTROWS[44]), .Z(
        CIPHERTEXT1[28]) );
  XOR2_X1 RF1_MC_U20 ( .A(RF1_SHIFTROWS[27]), .B(RF1_SHIFTROWS[43]), .Z(
        CIPHERTEXT1[27]) );
  XOR2_X1 RF1_MC_U19 ( .A(RF1_SHIFTROWS[26]), .B(RF1_SHIFTROWS[42]), .Z(
        CIPHERTEXT1[26]) );
  XOR2_X1 RF1_MC_U18 ( .A(RF1_SHIFTROWS[25]), .B(RF1_SHIFTROWS[41]), .Z(
        CIPHERTEXT1[25]) );
  XOR2_X1 RF1_MC_U17 ( .A(RF1_SHIFTROWS[24]), .B(RF1_SHIFTROWS[40]), .Z(
        CIPHERTEXT1[24]) );
  XOR2_X1 RF1_MC_U16 ( .A(RF1_SHIFTROWS[23]), .B(RF1_SHIFTROWS[39]), .Z(
        CIPHERTEXT1[23]) );
  XOR2_X1 RF1_MC_U15 ( .A(RF1_SHIFTROWS[22]), .B(RF1_SHIFTROWS[38]), .Z(
        CIPHERTEXT1[22]) );
  XOR2_X1 RF1_MC_U14 ( .A(RF1_SHIFTROWS[21]), .B(RF1_SHIFTROWS[37]), .Z(
        CIPHERTEXT1[21]) );
  XOR2_X1 RF1_MC_U13 ( .A(RF1_SHIFTROWS[20]), .B(RF1_SHIFTROWS[36]), .Z(
        CIPHERTEXT1[20]) );
  XOR2_X1 RF1_MC_U12 ( .A(CIPHERTEXT1[33]), .B(RF1_SHIFTROWS[17]), .Z(
        CIPHERTEXT1[1]) );
  XOR2_X1 RF1_MC_U11 ( .A(RF1_SHIFTROWS[19]), .B(RF1_SHIFTROWS[35]), .Z(
        CIPHERTEXT1[19]) );
  XOR2_X1 RF1_MC_U10 ( .A(RF1_SHIFTROWS[18]), .B(RF1_SHIFTROWS[34]), .Z(
        CIPHERTEXT1[18]) );
  XOR2_X1 RF1_MC_U9 ( .A(RF1_SHIFTROWS[17]), .B(RF1_SHIFTROWS[33]), .Z(
        CIPHERTEXT1[17]) );
  XOR2_X1 RF1_MC_U8 ( .A(RF1_SHIFTROWS[16]), .B(RF1_SHIFTROWS[32]), .Z(
        CIPHERTEXT1[16]) );
  XOR2_X1 RF1_MC_U7 ( .A(RF1_SHIFTROWS[31]), .B(CIPHERTEXT1[47]), .Z(
        CIPHERTEXT1[15]) );
  XOR2_X1 RF1_MC_U6 ( .A(RF1_SHIFTROWS[30]), .B(CIPHERTEXT1[46]), .Z(
        CIPHERTEXT1[14]) );
  XOR2_X1 RF1_MC_U5 ( .A(RF1_SHIFTROWS[29]), .B(CIPHERTEXT1[45]), .Z(
        CIPHERTEXT1[13]) );
  XOR2_X1 RF1_MC_U4 ( .A(RF1_SHIFTROWS[28]), .B(CIPHERTEXT1[44]), .Z(
        CIPHERTEXT1[12]) );
  XOR2_X1 RF1_MC_U3 ( .A(RF1_SHIFTROWS[27]), .B(CIPHERTEXT1[43]), .Z(
        CIPHERTEXT1[11]) );
  XOR2_X1 RF1_MC_U2 ( .A(RF1_SHIFTROWS[26]), .B(CIPHERTEXT1[42]), .Z(
        CIPHERTEXT1[10]) );
  XOR2_X1 RF1_MC_U1 ( .A(RF1_SHIFTROWS[16]), .B(CIPHERTEXT1[32]), .Z(
        CIPHERTEXT1[0]) );
  SDFF_X1 RF2_RS_SFF_0_Q_reg ( .D(CIPHERTEXT2[0]), .SI(PLAINTEXT2[0]), .SE(
        RESET), .CK(CLK), .Q(S_0_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_1_Q_reg ( .D(CIPHERTEXT2[1]), .SI(PLAINTEXT2[1]), .SE(
        RESET), .CK(CLK), .Q(S_0_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_2_Q_reg ( .D(CIPHERTEXT2[2]), .SI(PLAINTEXT2[2]), .SE(
        RESET), .CK(CLK), .Q(S_0_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_3_Q_reg ( .D(CIPHERTEXT2[3]), .SI(PLAINTEXT2[3]), .SE(
        RESET), .CK(CLK), .Q(S_0_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_4_Q_reg ( .D(CIPHERTEXT2[4]), .SI(PLAINTEXT2[4]), .SE(
        RESET), .CK(CLK), .Q(S_1_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_5_Q_reg ( .D(CIPHERTEXT2[5]), .SI(PLAINTEXT2[5]), .SE(
        RESET), .CK(CLK), .Q(S_1_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_6_Q_reg ( .D(CIPHERTEXT2[6]), .SI(PLAINTEXT2[6]), .SE(
        RESET), .CK(CLK), .Q(S_1_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_7_Q_reg ( .D(CIPHERTEXT2[7]), .SI(PLAINTEXT2[7]), .SE(
        RESET), .CK(CLK), .Q(S_1_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_8_Q_reg ( .D(CIPHERTEXT2[8]), .SI(PLAINTEXT2[8]), .SE(
        RESET), .CK(CLK), .Q(S_2_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_9_Q_reg ( .D(CIPHERTEXT2[9]), .SI(PLAINTEXT2[9]), .SE(
        RESET), .CK(CLK), .Q(S_2_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_10_Q_reg ( .D(CIPHERTEXT2[10]), .SI(PLAINTEXT2[10]), .SE(
        RESET), .CK(CLK), .Q(S_2_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_11_Q_reg ( .D(CIPHERTEXT2[11]), .SI(PLAINTEXT2[11]), .SE(
        RESET), .CK(CLK), .Q(S_2_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_12_Q_reg ( .D(CIPHERTEXT2[12]), .SI(PLAINTEXT2[12]), .SE(
        RESET), .CK(CLK), .Q(S_3_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_13_Q_reg ( .D(CIPHERTEXT2[13]), .SI(PLAINTEXT2[13]), .SE(
        RESET), .CK(CLK), .Q(S_3_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_14_Q_reg ( .D(CIPHERTEXT2[14]), .SI(PLAINTEXT2[14]), .SE(
        RESET), .CK(CLK), .Q(S_3_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_15_Q_reg ( .D(CIPHERTEXT2[15]), .SI(PLAINTEXT2[15]), .SE(
        RESET), .CK(CLK), .Q(S_3_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_16_Q_reg ( .D(CIPHERTEXT2[16]), .SI(PLAINTEXT2[16]), .SE(
        RESET), .CK(CLK), .Q(S_4_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_17_Q_reg ( .D(CIPHERTEXT2[17]), .SI(PLAINTEXT2[17]), .SE(
        RESET), .CK(CLK), .Q(S_4_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_18_Q_reg ( .D(CIPHERTEXT2[18]), .SI(PLAINTEXT2[18]), .SE(
        RESET), .CK(CLK), .Q(S_4_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_19_Q_reg ( .D(CIPHERTEXT2[19]), .SI(PLAINTEXT2[19]), .SE(
        RESET), .CK(CLK), .Q(S_4_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_20_Q_reg ( .D(CIPHERTEXT2[20]), .SI(PLAINTEXT2[20]), .SE(
        RESET), .CK(CLK), .Q(S_5_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_21_Q_reg ( .D(CIPHERTEXT2[21]), .SI(PLAINTEXT2[21]), .SE(
        RESET), .CK(CLK), .Q(S_5_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_22_Q_reg ( .D(CIPHERTEXT2[22]), .SI(PLAINTEXT2[22]), .SE(
        RESET), .CK(CLK), .Q(S_5_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_23_Q_reg ( .D(CIPHERTEXT2[23]), .SI(PLAINTEXT2[23]), .SE(
        RESET), .CK(CLK), .Q(S_5_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_24_Q_reg ( .D(CIPHERTEXT2[24]), .SI(PLAINTEXT2[24]), .SE(
        RESET), .CK(CLK), .Q(S_6_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_25_Q_reg ( .D(CIPHERTEXT2[25]), .SI(PLAINTEXT2[25]), .SE(
        RESET), .CK(CLK), .Q(S_6_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_26_Q_reg ( .D(CIPHERTEXT2[26]), .SI(PLAINTEXT2[26]), .SE(
        RESET), .CK(CLK), .Q(S_6_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_27_Q_reg ( .D(CIPHERTEXT2[27]), .SI(PLAINTEXT2[27]), .SE(
        RESET), .CK(CLK), .Q(S_6_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_28_Q_reg ( .D(CIPHERTEXT2[28]), .SI(PLAINTEXT2[28]), .SE(
        RESET), .CK(CLK), .Q(S_7_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_29_Q_reg ( .D(CIPHERTEXT2[29]), .SI(PLAINTEXT2[29]), .SE(
        RESET), .CK(CLK), .Q(S_7_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_30_Q_reg ( .D(CIPHERTEXT2[30]), .SI(PLAINTEXT2[30]), .SE(
        RESET), .CK(CLK), .Q(S_7_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_31_Q_reg ( .D(CIPHERTEXT2[31]), .SI(PLAINTEXT2[31]), .SE(
        RESET), .CK(CLK), .Q(S_7_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_32_Q_reg ( .D(CIPHERTEXT2[32]), .SI(PLAINTEXT2[32]), .SE(
        RESET), .CK(CLK), .Q(S_8_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_33_Q_reg ( .D(CIPHERTEXT2[33]), .SI(PLAINTEXT2[33]), .SE(
        RESET), .CK(CLK), .Q(S_8_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_34_Q_reg ( .D(CIPHERTEXT2[34]), .SI(PLAINTEXT2[34]), .SE(
        RESET), .CK(CLK), .Q(S_8_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_35_Q_reg ( .D(CIPHERTEXT2[35]), .SI(PLAINTEXT2[35]), .SE(
        RESET), .CK(CLK), .Q(S_8_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_36_Q_reg ( .D(CIPHERTEXT2[36]), .SI(PLAINTEXT2[36]), .SE(
        RESET), .CK(CLK), .Q(S_9_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_37_Q_reg ( .D(CIPHERTEXT2[37]), .SI(PLAINTEXT2[37]), .SE(
        RESET), .CK(CLK), .Q(S_9_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_38_Q_reg ( .D(CIPHERTEXT2[38]), .SI(PLAINTEXT2[38]), .SE(
        RESET), .CK(CLK), .Q(S_9_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_39_Q_reg ( .D(CIPHERTEXT2[39]), .SI(PLAINTEXT2[39]), .SE(
        RESET), .CK(CLK), .Q(S_9_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_40_Q_reg ( .D(CIPHERTEXT2[40]), .SI(PLAINTEXT2[40]), .SE(
        RESET), .CK(CLK), .Q(S_10_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_41_Q_reg ( .D(CIPHERTEXT2[41]), .SI(PLAINTEXT2[41]), .SE(
        RESET), .CK(CLK), .Q(S_10_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_42_Q_reg ( .D(CIPHERTEXT2[42]), .SI(PLAINTEXT2[42]), .SE(
        RESET), .CK(CLK), .Q(S_10_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_43_Q_reg ( .D(CIPHERTEXT2[43]), .SI(PLAINTEXT2[43]), .SE(
        RESET), .CK(CLK), .Q(S_10_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_44_Q_reg ( .D(CIPHERTEXT2[44]), .SI(PLAINTEXT2[44]), .SE(
        RESET), .CK(CLK), .Q(S_11_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_45_Q_reg ( .D(CIPHERTEXT2[45]), .SI(PLAINTEXT2[45]), .SE(
        RESET), .CK(CLK), .Q(S_11_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_46_Q_reg ( .D(CIPHERTEXT2[46]), .SI(PLAINTEXT2[46]), .SE(
        RESET), .CK(CLK), .Q(S_11_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_47_Q_reg ( .D(CIPHERTEXT2[47]), .SI(PLAINTEXT2[47]), .SE(
        RESET), .CK(CLK), .Q(S_11_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_48_Q_reg ( .D(CIPHERTEXT2[48]), .SI(PLAINTEXT2[48]), .SE(
        RESET), .CK(CLK), .Q(S_12_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_49_Q_reg ( .D(CIPHERTEXT2[49]), .SI(PLAINTEXT2[49]), .SE(
        RESET), .CK(CLK), .Q(S_12_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_50_Q_reg ( .D(CIPHERTEXT2[50]), .SI(PLAINTEXT2[50]), .SE(
        RESET), .CK(CLK), .Q(S_12_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_51_Q_reg ( .D(CIPHERTEXT2[51]), .SI(PLAINTEXT2[51]), .SE(
        RESET), .CK(CLK), .Q(S_12_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_52_Q_reg ( .D(CIPHERTEXT2[52]), .SI(PLAINTEXT2[52]), .SE(
        RESET), .CK(CLK), .Q(S_13_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_53_Q_reg ( .D(CIPHERTEXT2[53]), .SI(PLAINTEXT2[53]), .SE(
        RESET), .CK(CLK), .Q(S_13_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_54_Q_reg ( .D(CIPHERTEXT2[54]), .SI(PLAINTEXT2[54]), .SE(
        RESET), .CK(CLK), .Q(S_13_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_55_Q_reg ( .D(CIPHERTEXT2[55]), .SI(PLAINTEXT2[55]), .SE(
        RESET), .CK(CLK), .Q(S_13_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_56_Q_reg ( .D(CIPHERTEXT2[56]), .SI(PLAINTEXT2[56]), .SE(
        RESET), .CK(CLK), .Q(S_14_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_57_Q_reg ( .D(CIPHERTEXT2[57]), .SI(PLAINTEXT2[57]), .SE(
        RESET), .CK(CLK), .Q(S_14_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_58_Q_reg ( .D(CIPHERTEXT2[58]), .SI(PLAINTEXT2[58]), .SE(
        RESET), .CK(CLK), .Q(S_14_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_59_Q_reg ( .D(CIPHERTEXT2[59]), .SI(PLAINTEXT2[59]), .SE(
        RESET), .CK(CLK), .Q(S_14_F_in2[1]), .QN() );
  SDFF_X1 RF2_RS_SFF_60_Q_reg ( .D(CIPHERTEXT2[60]), .SI(PLAINTEXT2[60]), .SE(
        RESET), .CK(CLK), .Q(S_15_F_in2[0]), .QN() );
  SDFF_X1 RF2_RS_SFF_61_Q_reg ( .D(CIPHERTEXT2[61]), .SI(PLAINTEXT2[61]), .SE(
        RESET), .CK(CLK), .Q(S_15_F_in2[2]), .QN() );
  SDFF_X1 RF2_RS_SFF_62_Q_reg ( .D(CIPHERTEXT2[62]), .SI(PLAINTEXT2[62]), .SE(
        RESET), .CK(CLK), .Q(S_15_F_in2[3]), .QN() );
  SDFF_X1 RF2_RS_SFF_63_Q_reg ( .D(CIPHERTEXT2[63]), .SI(PLAINTEXT2[63]), .SE(
        RESET), .CK(CLK), .Q(S_15_F_in2[1]), .QN() );
  INV_X1 RF2_KA_U39 ( .A(SUB_OUT2[29]), .ZN(RF2_SHIFTROWS[21]) );
  XNOR2_X1 RF2_KA_U38 ( .A(RF2_KA_n18), .B(KE2_KEY_PERM[31]), .ZN(
        CIPHERTEXT2[47]) );
  XNOR2_X1 RF2_KA_U37 ( .A(1'b0), .B(SUB_OUT2[63]), .ZN(RF2_KA_n18) );
  XNOR2_X1 RF2_KA_U36 ( .A(RF2_KA_n17), .B(KE2_KEY_PERM[30]), .ZN(
        CIPHERTEXT2[46]) );
  XNOR2_X1 RF2_KA_U35 ( .A(1'b0), .B(SUB_OUT2[62]), .ZN(RF2_KA_n17) );
  XNOR2_X1 RF2_KA_U34 ( .A(RF2_KA_n16), .B(KE2_KEY_PERM[29]), .ZN(
        CIPHERTEXT2[45]) );
  XNOR2_X1 RF2_KA_U33 ( .A(1'b0), .B(SUB_OUT2[61]), .ZN(RF2_KA_n16) );
  XNOR2_X1 RF2_KA_U32 ( .A(RF2_KA_n15), .B(KE2_KEY_PERM[28]), .ZN(
        CIPHERTEXT2[44]) );
  XNOR2_X1 RF2_KA_U31 ( .A(1'b0), .B(SUB_OUT2[60]), .ZN(RF2_KA_n15) );
  XOR2_X1 RF2_KA_U30 ( .A(SUB_OUT2[59]), .B(KE2_KEY_PERM[27]), .Z(
        CIPHERTEXT2[43]) );
  XOR2_X1 RF2_KA_U29 ( .A(SUB_OUT2[58]), .B(KE2_KEY_PERM[26]), .Z(
        CIPHERTEXT2[42]) );
  XOR2_X1 RF2_KA_U28 ( .A(SUB_OUT2[57]), .B(KE2_KEY_PERM[25]), .Z(
        CIPHERTEXT2[41]) );
  XOR2_X1 RF2_KA_U27 ( .A(SUB_OUT2[56]), .B(KE2_KEY_PERM[24]), .Z(
        CIPHERTEXT2[40]) );
  XOR2_X1 RF2_KA_U26 ( .A(SUB_OUT2[55]), .B(KE2_KEY_PERM[23]), .Z(
        CIPHERTEXT2[39]) );
  XOR2_X1 RF2_KA_U25 ( .A(SUB_OUT2[54]), .B(KE2_KEY_PERM[22]), .Z(
        CIPHERTEXT2[38]) );
  XOR2_X1 RF2_KA_U24 ( .A(SUB_OUT2[53]), .B(KE2_KEY_PERM[21]), .Z(
        CIPHERTEXT2[37]) );
  XOR2_X1 RF2_KA_U23 ( .A(SUB_OUT2[52]), .B(KE2_KEY_PERM[20]), .Z(
        CIPHERTEXT2[36]) );
  XOR2_X1 RF2_KA_U22 ( .A(SUB_OUT2[51]), .B(KE2_KEY_PERM[19]), .Z(
        CIPHERTEXT2[35]) );
  XOR2_X1 RF2_KA_U21 ( .A(SUB_OUT2[50]), .B(KE2_KEY_PERM[18]), .Z(
        CIPHERTEXT2[34]) );
  XOR2_X1 RF2_KA_U20 ( .A(SUB_OUT2[49]), .B(KE2_KEY_PERM[17]), .Z(
        CIPHERTEXT2[33]) );
  XOR2_X1 RF2_KA_U19 ( .A(SUB_OUT2[48]), .B(KE2_KEY_PERM[16]), .Z(
        CIPHERTEXT2[32]) );
  XOR2_X1 RF2_KA_U18 ( .A(SUB_OUT2[47]), .B(KE2_KEY_PERM[15]), .Z(
        RF2_SHIFTROWS[43]) );
  XOR2_X1 RF2_KA_U17 ( .A(SUB_OUT2[46]), .B(KE2_KEY_PERM[14]), .Z(
        RF2_SHIFTROWS[42]) );
  XNOR2_X1 RF2_KA_U16 ( .A(RF2_KA_n14), .B(KE2_KEY_PERM[13]), .ZN(
        RF2_SHIFTROWS[41]) );
  XNOR2_X1 RF2_KA_U15 ( .A(1'b0), .B(SUB_OUT2[45]), .ZN(RF2_KA_n14) );
  XNOR2_X1 RF2_KA_U14 ( .A(RF2_KA_n13), .B(KE2_KEY_PERM[12]), .ZN(
        RF2_SHIFTROWS[40]) );
  XNOR2_X1 RF2_KA_U13 ( .A(1'b0), .B(SUB_OUT2[44]), .ZN(RF2_KA_n13) );
  XOR2_X1 RF2_KA_U12 ( .A(SUB_OUT2[43]), .B(KE2_KEY_PERM[11]), .Z(
        RF2_SHIFTROWS[39]) );
  XOR2_X1 RF2_KA_U11 ( .A(SUB_OUT2[42]), .B(KE2_KEY_PERM[10]), .Z(
        RF2_SHIFTROWS[38]) );
  XOR2_X1 RF2_KA_U10 ( .A(SUB_OUT2[41]), .B(KE2_KEY_PERM[9]), .Z(
        RF2_SHIFTROWS[37]) );
  XOR2_X1 RF2_KA_U9 ( .A(SUB_OUT2[40]), .B(KE2_KEY_PERM[8]), .Z(
        RF2_SHIFTROWS[36]) );
  XOR2_X1 RF2_KA_U8 ( .A(SUB_OUT2[39]), .B(KE2_KEY_PERM[7]), .Z(
        RF2_SHIFTROWS[35]) );
  XOR2_X1 RF2_KA_U7 ( .A(SUB_OUT2[38]), .B(KE2_KEY_PERM[6]), .Z(
        RF2_SHIFTROWS[34]) );
  XOR2_X1 RF2_KA_U6 ( .A(SUB_OUT2[37]), .B(KE2_KEY_PERM[5]), .Z(
        RF2_SHIFTROWS[33]) );
  XOR2_X1 RF2_KA_U5 ( .A(SUB_OUT2[36]), .B(KE2_KEY_PERM[4]), .Z(
        RF2_SHIFTROWS[32]) );
  XOR2_X1 RF2_KA_U4 ( .A(SUB_OUT2[35]), .B(KE2_KEY_PERM[3]), .Z(
        RF2_SHIFTROWS[47]) );
  XOR2_X1 RF2_KA_U3 ( .A(SUB_OUT2[34]), .B(KE2_KEY_PERM[2]), .Z(
        RF2_SHIFTROWS[46]) );
  XOR2_X1 RF2_KA_U2 ( .A(SUB_OUT2[33]), .B(KE2_KEY_PERM[1]), .Z(
        RF2_SHIFTROWS[45]) );
  XOR2_X1 RF2_KA_U1 ( .A(SUB_OUT2[32]), .B(KE2_KEY_PERM[0]), .Z(
        RF2_SHIFTROWS[44]) );
  XOR2_X1 RF2_MC_U48 ( .A(RF2_SHIFTROWS[15]), .B(CIPHERTEXT2[15]), .Z(
        CIPHERTEXT2[63]) );
  XOR2_X1 RF2_MC_U47 ( .A(RF2_SHIFTROWS[14]), .B(CIPHERTEXT2[14]), .Z(
        CIPHERTEXT2[62]) );
  XOR2_X1 RF2_MC_U46 ( .A(RF2_SHIFTROWS[13]), .B(CIPHERTEXT2[13]), .Z(
        CIPHERTEXT2[61]) );
  XOR2_X1 RF2_MC_U45 ( .A(RF2_SHIFTROWS[12]), .B(CIPHERTEXT2[12]), .Z(
        CIPHERTEXT2[60]) );
  XOR2_X1 RF2_MC_U44 ( .A(RF2_SHIFTROWS[11]), .B(CIPHERTEXT2[11]), .Z(
        CIPHERTEXT2[59]) );
  XOR2_X1 RF2_MC_U43 ( .A(RF2_SHIFTROWS[10]), .B(CIPHERTEXT2[10]), .Z(
        CIPHERTEXT2[58]) );
  XOR2_X1 RF2_MC_U42 ( .A(RF2_SHIFTROWS[9]), .B(CIPHERTEXT2[9]), .Z(
        CIPHERTEXT2[57]) );
  XOR2_X1 RF2_MC_U41 ( .A(CIPHERTEXT2[41]), .B(RF2_SHIFTROWS[25]), .Z(
        CIPHERTEXT2[9]) );
  XOR2_X1 RF2_MC_U40 ( .A(RF2_SHIFTROWS[8]), .B(CIPHERTEXT2[8]), .Z(
        CIPHERTEXT2[56]) );
  XOR2_X1 RF2_MC_U39 ( .A(CIPHERTEXT2[40]), .B(RF2_SHIFTROWS[24]), .Z(
        CIPHERTEXT2[8]) );
  XOR2_X1 RF2_MC_U38 ( .A(RF2_SHIFTROWS[7]), .B(CIPHERTEXT2[7]), .Z(
        CIPHERTEXT2[55]) );
  XOR2_X1 RF2_MC_U37 ( .A(CIPHERTEXT2[39]), .B(RF2_SHIFTROWS[23]), .Z(
        CIPHERTEXT2[7]) );
  XOR2_X1 RF2_MC_U36 ( .A(RF2_SHIFTROWS[6]), .B(CIPHERTEXT2[6]), .Z(
        CIPHERTEXT2[54]) );
  XOR2_X1 RF2_MC_U35 ( .A(CIPHERTEXT2[38]), .B(RF2_SHIFTROWS[22]), .Z(
        CIPHERTEXT2[6]) );
  XOR2_X1 RF2_MC_U34 ( .A(RF2_SHIFTROWS[5]), .B(CIPHERTEXT2[5]), .Z(
        CIPHERTEXT2[53]) );
  XOR2_X1 RF2_MC_U33 ( .A(CIPHERTEXT2[37]), .B(RF2_SHIFTROWS[21]), .Z(
        CIPHERTEXT2[5]) );
  XOR2_X1 RF2_MC_U32 ( .A(RF2_SHIFTROWS[4]), .B(CIPHERTEXT2[4]), .Z(
        CIPHERTEXT2[52]) );
  XOR2_X1 RF2_MC_U31 ( .A(RF2_SHIFTROWS[3]), .B(CIPHERTEXT2[3]), .Z(
        CIPHERTEXT2[51]) );
  XOR2_X1 RF2_MC_U30 ( .A(RF2_SHIFTROWS[2]), .B(CIPHERTEXT2[2]), .Z(
        CIPHERTEXT2[50]) );
  XOR2_X1 RF2_MC_U29 ( .A(CIPHERTEXT2[36]), .B(RF2_SHIFTROWS[20]), .Z(
        CIPHERTEXT2[4]) );
  XOR2_X1 RF2_MC_U28 ( .A(RF2_SHIFTROWS[1]), .B(CIPHERTEXT2[1]), .Z(
        CIPHERTEXT2[49]) );
  XOR2_X1 RF2_MC_U27 ( .A(RF2_SHIFTROWS[0]), .B(CIPHERTEXT2[0]), .Z(
        CIPHERTEXT2[48]) );
  XOR2_X1 RF2_MC_U26 ( .A(CIPHERTEXT2[35]), .B(RF2_SHIFTROWS[19]), .Z(
        CIPHERTEXT2[3]) );
  XOR2_X1 RF2_MC_U25 ( .A(RF2_SHIFTROWS[31]), .B(RF2_SHIFTROWS[47]), .Z(
        CIPHERTEXT2[31]) );
  XOR2_X1 RF2_MC_U24 ( .A(RF2_SHIFTROWS[30]), .B(RF2_SHIFTROWS[46]), .Z(
        CIPHERTEXT2[30]) );
  XOR2_X1 RF2_MC_U23 ( .A(CIPHERTEXT2[34]), .B(RF2_SHIFTROWS[18]), .Z(
        CIPHERTEXT2[2]) );
  XOR2_X1 RF2_MC_U22 ( .A(RF2_SHIFTROWS[29]), .B(RF2_SHIFTROWS[45]), .Z(
        CIPHERTEXT2[29]) );
  XOR2_X1 RF2_MC_U21 ( .A(RF2_SHIFTROWS[28]), .B(RF2_SHIFTROWS[44]), .Z(
        CIPHERTEXT2[28]) );
  XOR2_X1 RF2_MC_U20 ( .A(RF2_SHIFTROWS[27]), .B(RF2_SHIFTROWS[43]), .Z(
        CIPHERTEXT2[27]) );
  XOR2_X1 RF2_MC_U19 ( .A(RF2_SHIFTROWS[26]), .B(RF2_SHIFTROWS[42]), .Z(
        CIPHERTEXT2[26]) );
  XOR2_X1 RF2_MC_U18 ( .A(RF2_SHIFTROWS[25]), .B(RF2_SHIFTROWS[41]), .Z(
        CIPHERTEXT2[25]) );
  XOR2_X1 RF2_MC_U17 ( .A(RF2_SHIFTROWS[24]), .B(RF2_SHIFTROWS[40]), .Z(
        CIPHERTEXT2[24]) );
  XOR2_X1 RF2_MC_U16 ( .A(RF2_SHIFTROWS[23]), .B(RF2_SHIFTROWS[39]), .Z(
        CIPHERTEXT2[23]) );
  XOR2_X1 RF2_MC_U15 ( .A(RF2_SHIFTROWS[22]), .B(RF2_SHIFTROWS[38]), .Z(
        CIPHERTEXT2[22]) );
  XOR2_X1 RF2_MC_U14 ( .A(RF2_SHIFTROWS[21]), .B(RF2_SHIFTROWS[37]), .Z(
        CIPHERTEXT2[21]) );
  XOR2_X1 RF2_MC_U13 ( .A(RF2_SHIFTROWS[20]), .B(RF2_SHIFTROWS[36]), .Z(
        CIPHERTEXT2[20]) );
  XOR2_X1 RF2_MC_U12 ( .A(CIPHERTEXT2[33]), .B(RF2_SHIFTROWS[17]), .Z(
        CIPHERTEXT2[1]) );
  XOR2_X1 RF2_MC_U11 ( .A(RF2_SHIFTROWS[19]), .B(RF2_SHIFTROWS[35]), .Z(
        CIPHERTEXT2[19]) );
  XOR2_X1 RF2_MC_U10 ( .A(RF2_SHIFTROWS[18]), .B(RF2_SHIFTROWS[34]), .Z(
        CIPHERTEXT2[18]) );
  XOR2_X1 RF2_MC_U9 ( .A(RF2_SHIFTROWS[17]), .B(RF2_SHIFTROWS[33]), .Z(
        CIPHERTEXT2[17]) );
  XOR2_X1 RF2_MC_U8 ( .A(RF2_SHIFTROWS[16]), .B(RF2_SHIFTROWS[32]), .Z(
        CIPHERTEXT2[16]) );
  XOR2_X1 RF2_MC_U7 ( .A(RF2_SHIFTROWS[31]), .B(CIPHERTEXT2[47]), .Z(
        CIPHERTEXT2[15]) );
  XOR2_X1 RF2_MC_U6 ( .A(RF2_SHIFTROWS[30]), .B(CIPHERTEXT2[46]), .Z(
        CIPHERTEXT2[14]) );
  XOR2_X1 RF2_MC_U5 ( .A(RF2_SHIFTROWS[29]), .B(CIPHERTEXT2[45]), .Z(
        CIPHERTEXT2[13]) );
  XOR2_X1 RF2_MC_U4 ( .A(RF2_SHIFTROWS[28]), .B(CIPHERTEXT2[44]), .Z(
        CIPHERTEXT2[12]) );
  XOR2_X1 RF2_MC_U3 ( .A(RF2_SHIFTROWS[27]), .B(CIPHERTEXT2[43]), .Z(
        CIPHERTEXT2[11]) );
  XOR2_X1 RF2_MC_U2 ( .A(RF2_SHIFTROWS[26]), .B(CIPHERTEXT2[42]), .Z(
        CIPHERTEXT2[10]) );
  XOR2_X1 RF2_MC_U1 ( .A(RF2_SHIFTROWS[16]), .B(CIPHERTEXT2[32]), .Z(
        CIPHERTEXT2[0]) );
  SDFF_X1 RF3_RS_SFF_0_Q_reg ( .D(CIPHERTEXT3[0]), .SI(PLAINTEXT3[0]), .SE(
        RESET), .CK(CLK), .Q(S_0_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_1_Q_reg ( .D(CIPHERTEXT3[1]), .SI(PLAINTEXT3[1]), .SE(
        RESET), .CK(CLK), .Q(S_0_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_2_Q_reg ( .D(CIPHERTEXT3[2]), .SI(PLAINTEXT3[2]), .SE(
        RESET), .CK(CLK), .Q(S_0_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_3_Q_reg ( .D(CIPHERTEXT3[3]), .SI(PLAINTEXT3[3]), .SE(
        RESET), .CK(CLK), .Q(S_0_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_4_Q_reg ( .D(CIPHERTEXT3[4]), .SI(PLAINTEXT3[4]), .SE(
        RESET), .CK(CLK), .Q(S_1_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_5_Q_reg ( .D(CIPHERTEXT3[5]), .SI(PLAINTEXT3[5]), .SE(
        RESET), .CK(CLK), .Q(S_1_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_6_Q_reg ( .D(CIPHERTEXT3[6]), .SI(PLAINTEXT3[6]), .SE(
        RESET), .CK(CLK), .Q(S_1_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_7_Q_reg ( .D(CIPHERTEXT3[7]), .SI(PLAINTEXT3[7]), .SE(
        RESET), .CK(CLK), .Q(S_1_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_8_Q_reg ( .D(CIPHERTEXT3[8]), .SI(PLAINTEXT3[8]), .SE(
        RESET), .CK(CLK), .Q(S_2_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_9_Q_reg ( .D(CIPHERTEXT3[9]), .SI(PLAINTEXT3[9]), .SE(
        RESET), .CK(CLK), .Q(S_2_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_10_Q_reg ( .D(CIPHERTEXT3[10]), .SI(PLAINTEXT3[10]), .SE(
        RESET), .CK(CLK), .Q(S_2_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_11_Q_reg ( .D(CIPHERTEXT3[11]), .SI(PLAINTEXT3[11]), .SE(
        RESET), .CK(CLK), .Q(S_2_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_12_Q_reg ( .D(CIPHERTEXT3[12]), .SI(PLAINTEXT3[12]), .SE(
        RESET), .CK(CLK), .Q(S_3_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_13_Q_reg ( .D(CIPHERTEXT3[13]), .SI(PLAINTEXT3[13]), .SE(
        RESET), .CK(CLK), .Q(S_3_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_14_Q_reg ( .D(CIPHERTEXT3[14]), .SI(PLAINTEXT3[14]), .SE(
        RESET), .CK(CLK), .Q(S_3_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_15_Q_reg ( .D(CIPHERTEXT3[15]), .SI(PLAINTEXT3[15]), .SE(
        RESET), .CK(CLK), .Q(S_3_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_16_Q_reg ( .D(CIPHERTEXT3[16]), .SI(PLAINTEXT3[16]), .SE(
        RESET), .CK(CLK), .Q(S_4_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_17_Q_reg ( .D(CIPHERTEXT3[17]), .SI(PLAINTEXT3[17]), .SE(
        RESET), .CK(CLK), .Q(S_4_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_18_Q_reg ( .D(CIPHERTEXT3[18]), .SI(PLAINTEXT3[18]), .SE(
        RESET), .CK(CLK), .Q(S_4_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_19_Q_reg ( .D(CIPHERTEXT3[19]), .SI(PLAINTEXT3[19]), .SE(
        RESET), .CK(CLK), .Q(S_4_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_20_Q_reg ( .D(CIPHERTEXT3[20]), .SI(PLAINTEXT3[20]), .SE(
        RESET), .CK(CLK), .Q(S_5_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_21_Q_reg ( .D(CIPHERTEXT3[21]), .SI(PLAINTEXT3[21]), .SE(
        RESET), .CK(CLK), .Q(S_5_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_22_Q_reg ( .D(CIPHERTEXT3[22]), .SI(PLAINTEXT3[22]), .SE(
        RESET), .CK(CLK), .Q(S_5_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_23_Q_reg ( .D(CIPHERTEXT3[23]), .SI(PLAINTEXT3[23]), .SE(
        RESET), .CK(CLK), .Q(S_5_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_24_Q_reg ( .D(CIPHERTEXT3[24]), .SI(PLAINTEXT3[24]), .SE(
        RESET), .CK(CLK), .Q(S_6_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_25_Q_reg ( .D(CIPHERTEXT3[25]), .SI(PLAINTEXT3[25]), .SE(
        RESET), .CK(CLK), .Q(S_6_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_26_Q_reg ( .D(CIPHERTEXT3[26]), .SI(PLAINTEXT3[26]), .SE(
        RESET), .CK(CLK), .Q(S_6_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_27_Q_reg ( .D(CIPHERTEXT3[27]), .SI(PLAINTEXT3[27]), .SE(
        RESET), .CK(CLK), .Q(S_6_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_28_Q_reg ( .D(CIPHERTEXT3[28]), .SI(PLAINTEXT3[28]), .SE(
        RESET), .CK(CLK), .Q(S_7_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_29_Q_reg ( .D(CIPHERTEXT3[29]), .SI(PLAINTEXT3[29]), .SE(
        RESET), .CK(CLK), .Q(S_7_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_30_Q_reg ( .D(CIPHERTEXT3[30]), .SI(PLAINTEXT3[30]), .SE(
        RESET), .CK(CLK), .Q(S_7_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_31_Q_reg ( .D(CIPHERTEXT3[31]), .SI(PLAINTEXT3[31]), .SE(
        RESET), .CK(CLK), .Q(S_7_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_32_Q_reg ( .D(CIPHERTEXT3[32]), .SI(PLAINTEXT3[32]), .SE(
        RESET), .CK(CLK), .Q(S_8_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_33_Q_reg ( .D(CIPHERTEXT3[33]), .SI(PLAINTEXT3[33]), .SE(
        RESET), .CK(CLK), .Q(S_8_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_34_Q_reg ( .D(CIPHERTEXT3[34]), .SI(PLAINTEXT3[34]), .SE(
        RESET), .CK(CLK), .Q(S_8_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_35_Q_reg ( .D(CIPHERTEXT3[35]), .SI(PLAINTEXT3[35]), .SE(
        RESET), .CK(CLK), .Q(S_8_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_36_Q_reg ( .D(CIPHERTEXT3[36]), .SI(PLAINTEXT3[36]), .SE(
        RESET), .CK(CLK), .Q(S_9_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_37_Q_reg ( .D(CIPHERTEXT3[37]), .SI(PLAINTEXT3[37]), .SE(
        RESET), .CK(CLK), .Q(S_9_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_38_Q_reg ( .D(CIPHERTEXT3[38]), .SI(PLAINTEXT3[38]), .SE(
        RESET), .CK(CLK), .Q(S_9_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_39_Q_reg ( .D(CIPHERTEXT3[39]), .SI(PLAINTEXT3[39]), .SE(
        RESET), .CK(CLK), .Q(S_9_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_40_Q_reg ( .D(CIPHERTEXT3[40]), .SI(PLAINTEXT3[40]), .SE(
        RESET), .CK(CLK), .Q(S_10_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_41_Q_reg ( .D(CIPHERTEXT3[41]), .SI(PLAINTEXT3[41]), .SE(
        RESET), .CK(CLK), .Q(S_10_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_42_Q_reg ( .D(CIPHERTEXT3[42]), .SI(PLAINTEXT3[42]), .SE(
        RESET), .CK(CLK), .Q(S_10_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_43_Q_reg ( .D(CIPHERTEXT3[43]), .SI(PLAINTEXT3[43]), .SE(
        RESET), .CK(CLK), .Q(S_10_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_44_Q_reg ( .D(CIPHERTEXT3[44]), .SI(PLAINTEXT3[44]), .SE(
        RESET), .CK(CLK), .Q(S_11_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_45_Q_reg ( .D(CIPHERTEXT3[45]), .SI(PLAINTEXT3[45]), .SE(
        RESET), .CK(CLK), .Q(S_11_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_46_Q_reg ( .D(CIPHERTEXT3[46]), .SI(PLAINTEXT3[46]), .SE(
        RESET), .CK(CLK), .Q(S_11_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_47_Q_reg ( .D(CIPHERTEXT3[47]), .SI(PLAINTEXT3[47]), .SE(
        RESET), .CK(CLK), .Q(S_11_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_48_Q_reg ( .D(CIPHERTEXT3[48]), .SI(PLAINTEXT3[48]), .SE(
        RESET), .CK(CLK), .Q(S_12_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_49_Q_reg ( .D(CIPHERTEXT3[49]), .SI(PLAINTEXT3[49]), .SE(
        RESET), .CK(CLK), .Q(S_12_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_50_Q_reg ( .D(CIPHERTEXT3[50]), .SI(PLAINTEXT3[50]), .SE(
        RESET), .CK(CLK), .Q(S_12_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_51_Q_reg ( .D(CIPHERTEXT3[51]), .SI(PLAINTEXT3[51]), .SE(
        RESET), .CK(CLK), .Q(S_12_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_52_Q_reg ( .D(CIPHERTEXT3[52]), .SI(PLAINTEXT3[52]), .SE(
        RESET), .CK(CLK), .Q(S_13_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_53_Q_reg ( .D(CIPHERTEXT3[53]), .SI(PLAINTEXT3[53]), .SE(
        RESET), .CK(CLK), .Q(S_13_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_54_Q_reg ( .D(CIPHERTEXT3[54]), .SI(PLAINTEXT3[54]), .SE(
        RESET), .CK(CLK), .Q(S_13_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_55_Q_reg ( .D(CIPHERTEXT3[55]), .SI(PLAINTEXT3[55]), .SE(
        RESET), .CK(CLK), .Q(S_13_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_56_Q_reg ( .D(CIPHERTEXT3[56]), .SI(PLAINTEXT3[56]), .SE(
        RESET), .CK(CLK), .Q(S_14_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_57_Q_reg ( .D(CIPHERTEXT3[57]), .SI(PLAINTEXT3[57]), .SE(
        RESET), .CK(CLK), .Q(S_14_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_58_Q_reg ( .D(CIPHERTEXT3[58]), .SI(PLAINTEXT3[58]), .SE(
        RESET), .CK(CLK), .Q(S_14_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_59_Q_reg ( .D(CIPHERTEXT3[59]), .SI(PLAINTEXT3[59]), .SE(
        RESET), .CK(CLK), .Q(S_14_F_in3[1]), .QN() );
  SDFF_X1 RF3_RS_SFF_60_Q_reg ( .D(CIPHERTEXT3[60]), .SI(PLAINTEXT3[60]), .SE(
        RESET), .CK(CLK), .Q(S_15_F_in3[0]), .QN() );
  SDFF_X1 RF3_RS_SFF_61_Q_reg ( .D(CIPHERTEXT3[61]), .SI(PLAINTEXT3[61]), .SE(
        RESET), .CK(CLK), .Q(S_15_F_in3[2]), .QN() );
  SDFF_X1 RF3_RS_SFF_62_Q_reg ( .D(CIPHERTEXT3[62]), .SI(PLAINTEXT3[62]), .SE(
        RESET), .CK(CLK), .Q(S_15_F_in3[3]), .QN() );
  SDFF_X1 RF3_RS_SFF_63_Q_reg ( .D(CIPHERTEXT3[63]), .SI(PLAINTEXT3[63]), .SE(
        RESET), .CK(CLK), .Q(S_15_F_in3[1]), .QN() );
  INV_X1 RF3_KA_U39 ( .A(SUB_OUT3[29]), .ZN(RF3_SHIFTROWS[21]) );
  XNOR2_X1 RF3_KA_U38 ( .A(RF3_KA_n18), .B(KE3_KEY_PERM[31]), .ZN(
        CIPHERTEXT3[47]) );
  XNOR2_X1 RF3_KA_U37 ( .A(1'b0), .B(SUB_OUT3[63]), .ZN(RF3_KA_n18) );
  XNOR2_X1 RF3_KA_U36 ( .A(RF3_KA_n17), .B(KE3_KEY_PERM[30]), .ZN(
        CIPHERTEXT3[46]) );
  XNOR2_X1 RF3_KA_U35 ( .A(1'b0), .B(SUB_OUT3[62]), .ZN(RF3_KA_n17) );
  XNOR2_X1 RF3_KA_U34 ( .A(RF3_KA_n16), .B(KE3_KEY_PERM[29]), .ZN(
        CIPHERTEXT3[45]) );
  XNOR2_X1 RF3_KA_U33 ( .A(1'b0), .B(SUB_OUT3[61]), .ZN(RF3_KA_n16) );
  XNOR2_X1 RF3_KA_U32 ( .A(RF3_KA_n15), .B(KE3_KEY_PERM[28]), .ZN(
        CIPHERTEXT3[44]) );
  XNOR2_X1 RF3_KA_U31 ( .A(1'b0), .B(SUB_OUT3[60]), .ZN(RF3_KA_n15) );
  XOR2_X1 RF3_KA_U30 ( .A(SUB_OUT3[59]), .B(KE3_KEY_PERM[27]), .Z(
        CIPHERTEXT3[43]) );
  XOR2_X1 RF3_KA_U29 ( .A(SUB_OUT3[58]), .B(KE3_KEY_PERM[26]), .Z(
        CIPHERTEXT3[42]) );
  XOR2_X1 RF3_KA_U28 ( .A(SUB_OUT3[57]), .B(KE3_KEY_PERM[25]), .Z(
        CIPHERTEXT3[41]) );
  XOR2_X1 RF3_KA_U27 ( .A(SUB_OUT3[56]), .B(KE3_KEY_PERM[24]), .Z(
        CIPHERTEXT3[40]) );
  XOR2_X1 RF3_KA_U26 ( .A(SUB_OUT3[55]), .B(KE3_KEY_PERM[23]), .Z(
        CIPHERTEXT3[39]) );
  XOR2_X1 RF3_KA_U25 ( .A(SUB_OUT3[54]), .B(KE3_KEY_PERM[22]), .Z(
        CIPHERTEXT3[38]) );
  XOR2_X1 RF3_KA_U24 ( .A(SUB_OUT3[53]), .B(KE3_KEY_PERM[21]), .Z(
        CIPHERTEXT3[37]) );
  XOR2_X1 RF3_KA_U23 ( .A(SUB_OUT3[52]), .B(KE3_KEY_PERM[20]), .Z(
        CIPHERTEXT3[36]) );
  XOR2_X1 RF3_KA_U22 ( .A(SUB_OUT3[51]), .B(KE3_KEY_PERM[19]), .Z(
        CIPHERTEXT3[35]) );
  XOR2_X1 RF3_KA_U21 ( .A(SUB_OUT3[50]), .B(KE3_KEY_PERM[18]), .Z(
        CIPHERTEXT3[34]) );
  XOR2_X1 RF3_KA_U20 ( .A(SUB_OUT3[49]), .B(KE3_KEY_PERM[17]), .Z(
        CIPHERTEXT3[33]) );
  XOR2_X1 RF3_KA_U19 ( .A(SUB_OUT3[48]), .B(KE3_KEY_PERM[16]), .Z(
        CIPHERTEXT3[32]) );
  XOR2_X1 RF3_KA_U18 ( .A(SUB_OUT3[47]), .B(KE3_KEY_PERM[15]), .Z(
        RF3_SHIFTROWS[43]) );
  XOR2_X1 RF3_KA_U17 ( .A(SUB_OUT3[46]), .B(KE3_KEY_PERM[14]), .Z(
        RF3_SHIFTROWS[42]) );
  XNOR2_X1 RF3_KA_U16 ( .A(RF3_KA_n14), .B(KE3_KEY_PERM[13]), .ZN(
        RF3_SHIFTROWS[41]) );
  XNOR2_X1 RF3_KA_U15 ( .A(1'b0), .B(SUB_OUT3[45]), .ZN(RF3_KA_n14) );
  XNOR2_X1 RF3_KA_U14 ( .A(RF3_KA_n13), .B(KE3_KEY_PERM[12]), .ZN(
        RF3_SHIFTROWS[40]) );
  XNOR2_X1 RF3_KA_U13 ( .A(1'b0), .B(SUB_OUT3[44]), .ZN(RF3_KA_n13) );
  XOR2_X1 RF3_KA_U12 ( .A(SUB_OUT3[43]), .B(KE3_KEY_PERM[11]), .Z(
        RF3_SHIFTROWS[39]) );
  XOR2_X1 RF3_KA_U11 ( .A(SUB_OUT3[42]), .B(KE3_KEY_PERM[10]), .Z(
        RF3_SHIFTROWS[38]) );
  XOR2_X1 RF3_KA_U10 ( .A(SUB_OUT3[41]), .B(KE3_KEY_PERM[9]), .Z(
        RF3_SHIFTROWS[37]) );
  XOR2_X1 RF3_KA_U9 ( .A(SUB_OUT3[40]), .B(KE3_KEY_PERM[8]), .Z(
        RF3_SHIFTROWS[36]) );
  XOR2_X1 RF3_KA_U8 ( .A(SUB_OUT3[39]), .B(KE3_KEY_PERM[7]), .Z(
        RF3_SHIFTROWS[35]) );
  XOR2_X1 RF3_KA_U7 ( .A(SUB_OUT3[38]), .B(KE3_KEY_PERM[6]), .Z(
        RF3_SHIFTROWS[34]) );
  XOR2_X1 RF3_KA_U6 ( .A(SUB_OUT3[37]), .B(KE3_KEY_PERM[5]), .Z(
        RF3_SHIFTROWS[33]) );
  XOR2_X1 RF3_KA_U5 ( .A(SUB_OUT3[36]), .B(KE3_KEY_PERM[4]), .Z(
        RF3_SHIFTROWS[32]) );
  XOR2_X1 RF3_KA_U4 ( .A(SUB_OUT3[35]), .B(KE3_KEY_PERM[3]), .Z(
        RF3_SHIFTROWS[47]) );
  XOR2_X1 RF3_KA_U3 ( .A(SUB_OUT3[34]), .B(KE3_KEY_PERM[2]), .Z(
        RF3_SHIFTROWS[46]) );
  XOR2_X1 RF3_KA_U2 ( .A(SUB_OUT3[33]), .B(KE3_KEY_PERM[1]), .Z(
        RF3_SHIFTROWS[45]) );
  XOR2_X1 RF3_KA_U1 ( .A(SUB_OUT3[32]), .B(KE3_KEY_PERM[0]), .Z(
        RF3_SHIFTROWS[44]) );
  XOR2_X1 RF3_MC_U48 ( .A(RF3_SHIFTROWS[15]), .B(CIPHERTEXT3[15]), .Z(
        CIPHERTEXT3[63]) );
  XOR2_X1 RF3_MC_U47 ( .A(RF3_SHIFTROWS[14]), .B(CIPHERTEXT3[14]), .Z(
        CIPHERTEXT3[62]) );
  XOR2_X1 RF3_MC_U46 ( .A(RF3_SHIFTROWS[13]), .B(CIPHERTEXT3[13]), .Z(
        CIPHERTEXT3[61]) );
  XOR2_X1 RF3_MC_U45 ( .A(RF3_SHIFTROWS[12]), .B(CIPHERTEXT3[12]), .Z(
        CIPHERTEXT3[60]) );
  XOR2_X1 RF3_MC_U44 ( .A(RF3_SHIFTROWS[11]), .B(CIPHERTEXT3[11]), .Z(
        CIPHERTEXT3[59]) );
  XOR2_X1 RF3_MC_U43 ( .A(RF3_SHIFTROWS[10]), .B(CIPHERTEXT3[10]), .Z(
        CIPHERTEXT3[58]) );
  XOR2_X1 RF3_MC_U42 ( .A(RF3_SHIFTROWS[9]), .B(CIPHERTEXT3[9]), .Z(
        CIPHERTEXT3[57]) );
  XOR2_X1 RF3_MC_U41 ( .A(CIPHERTEXT3[41]), .B(RF3_SHIFTROWS[25]), .Z(
        CIPHERTEXT3[9]) );
  XOR2_X1 RF3_MC_U40 ( .A(RF3_SHIFTROWS[8]), .B(CIPHERTEXT3[8]), .Z(
        CIPHERTEXT3[56]) );
  XOR2_X1 RF3_MC_U39 ( .A(CIPHERTEXT3[40]), .B(RF3_SHIFTROWS[24]), .Z(
        CIPHERTEXT3[8]) );
  XOR2_X1 RF3_MC_U38 ( .A(RF3_SHIFTROWS[7]), .B(CIPHERTEXT3[7]), .Z(
        CIPHERTEXT3[55]) );
  XOR2_X1 RF3_MC_U37 ( .A(CIPHERTEXT3[39]), .B(RF3_SHIFTROWS[23]), .Z(
        CIPHERTEXT3[7]) );
  XOR2_X1 RF3_MC_U36 ( .A(RF3_SHIFTROWS[6]), .B(CIPHERTEXT3[6]), .Z(
        CIPHERTEXT3[54]) );
  XOR2_X1 RF3_MC_U35 ( .A(CIPHERTEXT3[38]), .B(RF3_SHIFTROWS[22]), .Z(
        CIPHERTEXT3[6]) );
  XOR2_X1 RF3_MC_U34 ( .A(RF3_SHIFTROWS[5]), .B(CIPHERTEXT3[5]), .Z(
        CIPHERTEXT3[53]) );
  XOR2_X1 RF3_MC_U33 ( .A(CIPHERTEXT3[37]), .B(RF3_SHIFTROWS[21]), .Z(
        CIPHERTEXT3[5]) );
  XOR2_X1 RF3_MC_U32 ( .A(RF3_SHIFTROWS[4]), .B(CIPHERTEXT3[4]), .Z(
        CIPHERTEXT3[52]) );
  XOR2_X1 RF3_MC_U31 ( .A(RF3_SHIFTROWS[3]), .B(CIPHERTEXT3[3]), .Z(
        CIPHERTEXT3[51]) );
  XOR2_X1 RF3_MC_U30 ( .A(RF3_SHIFTROWS[2]), .B(CIPHERTEXT3[2]), .Z(
        CIPHERTEXT3[50]) );
  XOR2_X1 RF3_MC_U29 ( .A(CIPHERTEXT3[36]), .B(RF3_SHIFTROWS[20]), .Z(
        CIPHERTEXT3[4]) );
  XOR2_X1 RF3_MC_U28 ( .A(RF3_SHIFTROWS[1]), .B(CIPHERTEXT3[1]), .Z(
        CIPHERTEXT3[49]) );
  XOR2_X1 RF3_MC_U27 ( .A(RF3_SHIFTROWS[0]), .B(CIPHERTEXT3[0]), .Z(
        CIPHERTEXT3[48]) );
  XOR2_X1 RF3_MC_U26 ( .A(CIPHERTEXT3[35]), .B(RF3_SHIFTROWS[19]), .Z(
        CIPHERTEXT3[3]) );
  XOR2_X1 RF3_MC_U25 ( .A(RF3_SHIFTROWS[31]), .B(RF3_SHIFTROWS[47]), .Z(
        CIPHERTEXT3[31]) );
  XOR2_X1 RF3_MC_U24 ( .A(RF3_SHIFTROWS[30]), .B(RF3_SHIFTROWS[46]), .Z(
        CIPHERTEXT3[30]) );
  XOR2_X1 RF3_MC_U23 ( .A(CIPHERTEXT3[34]), .B(RF3_SHIFTROWS[18]), .Z(
        CIPHERTEXT3[2]) );
  XOR2_X1 RF3_MC_U22 ( .A(RF3_SHIFTROWS[29]), .B(RF3_SHIFTROWS[45]), .Z(
        CIPHERTEXT3[29]) );
  XOR2_X1 RF3_MC_U21 ( .A(RF3_SHIFTROWS[28]), .B(RF3_SHIFTROWS[44]), .Z(
        CIPHERTEXT3[28]) );
  XOR2_X1 RF3_MC_U20 ( .A(RF3_SHIFTROWS[27]), .B(RF3_SHIFTROWS[43]), .Z(
        CIPHERTEXT3[27]) );
  XOR2_X1 RF3_MC_U19 ( .A(RF3_SHIFTROWS[26]), .B(RF3_SHIFTROWS[42]), .Z(
        CIPHERTEXT3[26]) );
  XOR2_X1 RF3_MC_U18 ( .A(RF3_SHIFTROWS[25]), .B(RF3_SHIFTROWS[41]), .Z(
        CIPHERTEXT3[25]) );
  XOR2_X1 RF3_MC_U17 ( .A(RF3_SHIFTROWS[24]), .B(RF3_SHIFTROWS[40]), .Z(
        CIPHERTEXT3[24]) );
  XOR2_X1 RF3_MC_U16 ( .A(RF3_SHIFTROWS[23]), .B(RF3_SHIFTROWS[39]), .Z(
        CIPHERTEXT3[23]) );
  XOR2_X1 RF3_MC_U15 ( .A(RF3_SHIFTROWS[22]), .B(RF3_SHIFTROWS[38]), .Z(
        CIPHERTEXT3[22]) );
  XOR2_X1 RF3_MC_U14 ( .A(RF3_SHIFTROWS[21]), .B(RF3_SHIFTROWS[37]), .Z(
        CIPHERTEXT3[21]) );
  XOR2_X1 RF3_MC_U13 ( .A(RF3_SHIFTROWS[20]), .B(RF3_SHIFTROWS[36]), .Z(
        CIPHERTEXT3[20]) );
  XOR2_X1 RF3_MC_U12 ( .A(CIPHERTEXT3[33]), .B(RF3_SHIFTROWS[17]), .Z(
        CIPHERTEXT3[1]) );
  XOR2_X1 RF3_MC_U11 ( .A(RF3_SHIFTROWS[19]), .B(RF3_SHIFTROWS[35]), .Z(
        CIPHERTEXT3[19]) );
  XOR2_X1 RF3_MC_U10 ( .A(RF3_SHIFTROWS[18]), .B(RF3_SHIFTROWS[34]), .Z(
        CIPHERTEXT3[18]) );
  XOR2_X1 RF3_MC_U9 ( .A(RF3_SHIFTROWS[17]), .B(RF3_SHIFTROWS[33]), .Z(
        CIPHERTEXT3[17]) );
  XOR2_X1 RF3_MC_U8 ( .A(RF3_SHIFTROWS[16]), .B(RF3_SHIFTROWS[32]), .Z(
        CIPHERTEXT3[16]) );
  XOR2_X1 RF3_MC_U7 ( .A(RF3_SHIFTROWS[31]), .B(CIPHERTEXT3[47]), .Z(
        CIPHERTEXT3[15]) );
  XOR2_X1 RF3_MC_U6 ( .A(RF3_SHIFTROWS[30]), .B(CIPHERTEXT3[46]), .Z(
        CIPHERTEXT3[14]) );
  XOR2_X1 RF3_MC_U5 ( .A(RF3_SHIFTROWS[29]), .B(CIPHERTEXT3[45]), .Z(
        CIPHERTEXT3[13]) );
  XOR2_X1 RF3_MC_U4 ( .A(RF3_SHIFTROWS[28]), .B(CIPHERTEXT3[44]), .Z(
        CIPHERTEXT3[12]) );
  XOR2_X1 RF3_MC_U3 ( .A(RF3_SHIFTROWS[27]), .B(CIPHERTEXT3[43]), .Z(
        CIPHERTEXT3[11]) );
  XOR2_X1 RF3_MC_U2 ( .A(RF3_SHIFTROWS[26]), .B(CIPHERTEXT3[42]), .Z(
        CIPHERTEXT3[10]) );
  XOR2_X1 RF3_MC_U1 ( .A(RF3_SHIFTROWS[16]), .B(CIPHERTEXT3[32]), .Z(
        CIPHERTEXT3[0]) );
  DFF_X1 S_0_Rq3_reg_0_ ( .D(S_0_q3[0]), .CK(CLK), .Q(S_0_Rq3[0]), .QN() );
  DFF_X1 S_0_Rq3_reg_1_ ( .D(S_0_q3[1]), .CK(CLK), .Q(S_0_Rq3[1]), .QN() );
  DFF_X1 S_0_Rq3_reg_2_ ( .D(S_0_q3[2]), .CK(CLK), .Q(S_0_Rq3[2]), .QN() );
  DFF_X1 S_0_Rq3_reg_3_ ( .D(S_0_q3[3]), .CK(CLK), .Q(S_0_Rq3[3]), .QN() );
  DFF_X1 S_0_Rq2_reg_0_ ( .D(S_0_q2[0]), .CK(CLK), .Q(S_0_Rq2[0]), .QN() );
  DFF_X1 S_0_Rq2_reg_1_ ( .D(S_0_q2[1]), .CK(CLK), .Q(S_0_Rq2[1]), .QN() );
  DFF_X1 S_0_Rq2_reg_2_ ( .D(S_0_q2[2]), .CK(CLK), .Q(S_0_Rq2[2]), .QN() );
  DFF_X1 S_0_Rq2_reg_3_ ( .D(S_0_q2[3]), .CK(CLK), .Q(S_0_Rq2[3]), .QN() );
  DFF_X1 S_0_Rq1_reg_0_ ( .D(S_0_q1[0]), .CK(CLK), .Q(S_0_Rq1[0]), .QN() );
  DFF_X1 S_0_Rq1_reg_1_ ( .D(S_0_q1[1]), .CK(CLK), .Q(S_0_Rq1[1]), .QN() );
  DFF_X1 S_0_Rq1_reg_2_ ( .D(S_0_q1[2]), .CK(CLK), .Q(S_0_Rq1[2]), .QN() );
  DFF_X1 S_0_Rq1_reg_3_ ( .D(S_0_q1[3]), .CK(CLK), .Q(S_0_Rq1[3]), .QN() );
  INV_X1 S_0_InputAffine_U4 ( .A(SUB_IN1[0]), .ZN(S_0_F_in1[0]) );
  INV_X1 S_0_InputAffine_U3 ( .A(SUB_IN1[2]), .ZN(S_0_F_in1[3]) );
  INV_X1 S_0_InputAffine_U2 ( .A(SUB_IN1[3]), .ZN(S_0_F_in1[1]) );
  INV_X1 S_0_InputAffine_U1 ( .A(SUB_IN1[1]), .ZN(S_0_F_in1[2]) );
  XNOR2_X1 S_0_F_U18 ( .A(S_0_F_n4), .B(FRESH[3]), .ZN(S_0_q3[3]) );
  XNOR2_X1 S_0_F_U17 ( .A(FRESH[2]), .B(S_0_F_q3[3]), .ZN(S_0_F_n4) );
  XNOR2_X1 S_0_F_U16 ( .A(S_0_F_n3), .B(FRESH[1]), .ZN(S_0_q3[2]) );
  XNOR2_X1 S_0_F_U15 ( .A(FRESH[0]), .B(S_0_F_q3[2]), .ZN(S_0_F_n3) );
  XOR2_X1 S_0_F_U14 ( .A(FRESH[3]), .B(S_0_F_q2[3]), .Z(S_0_q2[3]) );
  XOR2_X1 S_0_F_U13 ( .A(FRESH[1]), .B(S_0_F_q2[2]), .Z(S_0_q2[2]) );
  XOR2_X1 S_0_F_U12 ( .A(FRESH[2]), .B(S_0_F_q1[3]), .Z(S_0_q1[3]) );
  XOR2_X1 S_0_F_U11 ( .A(FRESH[0]), .B(S_0_F_q1[2]), .Z(S_0_q1[2]) );
  XNOR2_X1 S_0_F_U10 ( .A(S_0_F_n2), .B(FRESH[5]), .ZN(S_0_F_N5) );
  XNOR2_X1 S_0_F_U9 ( .A(S_0_F_in3[3]), .B(FRESH[4]), .ZN(S_0_F_n2) );
  XOR2_X1 S_0_F_U8 ( .A(FRESH[5]), .B(S_0_F_in2[3]), .Z(S_0_F_N4) );
  XOR2_X1 S_0_F_U7 ( .A(FRESH[4]), .B(S_0_F_in1[3]), .Z(S_0_F_N3) );
  XNOR2_X1 S_0_F_U6 ( .A(S_0_F_n1), .B(FRESH[7]), .ZN(S_0_F_N2) );
  XNOR2_X1 S_0_F_U5 ( .A(S_0_F_in3[2]), .B(FRESH[6]), .ZN(S_0_F_n1) );
  XOR2_X1 S_0_F_U4 ( .A(FRESH[7]), .B(S_0_F_in2[2]), .Z(S_0_F_N1) );
  XOR2_X1 S_0_F_U3 ( .A(FRESH[6]), .B(S_0_F_in1[2]), .Z(S_0_F_N0) );
  DFF_X1 S_0_F_CF_Reg_reg_0_ ( .D(S_0_F_CF_Out[0]), .CK(CLK), .Q(
        S_0_F_CF_Reg[0]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_1_ ( .D(S_0_F_CF_Out[1]), .CK(CLK), .Q(
        S_0_F_CF_Reg[1]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_2_ ( .D(S_0_F_CF_Out[2]), .CK(CLK), .Q(
        S_0_F_CF_Reg[2]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_3_ ( .D(S_0_F_CF_Out[3]), .CK(CLK), .Q(
        S_0_F_CF_Reg[3]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_4_ ( .D(S_0_F_CF_Out[4]), .CK(CLK), .Q(
        S_0_F_CF_Reg[4]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_5_ ( .D(S_0_F_CF_Out[5]), .CK(CLK), .Q(
        S_0_F_CF_Reg[5]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_6_ ( .D(S_0_F_CF_Out[6]), .CK(CLK), .Q(
        S_0_F_CF_Reg[6]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_7_ ( .D(S_0_F_CF_Out[7]), .CK(CLK), .Q(
        S_0_F_CF_Reg[7]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_8_ ( .D(S_0_F_CF_Out[8]), .CK(CLK), .Q(
        S_0_F_CF_Reg[8]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_9_ ( .D(S_0_F_CF_Out[9]), .CK(CLK), .Q(
        S_0_F_CF_Reg[9]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_10_ ( .D(S_0_F_CF_Out[10]), .CK(CLK), .Q(
        S_0_F_CF_Reg[10]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_11_ ( .D(S_0_F_CF_Out[11]), .CK(CLK), .Q(
        S_0_F_CF_Reg[11]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_12_ ( .D(S_0_F_CF_Out[12]), .CK(CLK), .Q(
        S_0_F_CF_Reg[12]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_13_ ( .D(S_0_F_CF_Out[13]), .CK(CLK), .Q(
        S_0_F_CF_Reg[13]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_14_ ( .D(S_0_F_CF_Out[14]), .CK(CLK), .Q(
        S_0_F_CF_Reg[14]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_15_ ( .D(S_0_F_CF_Out[15]), .CK(CLK), .Q(
        S_0_F_CF_Reg[15]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_16_ ( .D(S_0_F_CF_Out[16]), .CK(CLK), .Q(
        S_0_F_CF_Reg[16]), .QN() );
  DFF_X1 S_0_F_CF_Reg_reg_17_ ( .D(S_0_F_CF_Out[17]), .CK(CLK), .Q(
        S_0_F_CF_Reg[17]), .QN() );
  DFF_X1 S_0_F_out2_reg_0_ ( .D(S_0_F_N4), .CK(CLK), .Q(S_0_q2[0]), .QN() );
  DFF_X1 S_0_F_out2_reg_1_ ( .D(S_0_F_N1), .CK(CLK), .Q(S_0_q2[1]), .QN() );
  DFF_X1 S_0_F_out3_reg_0_ ( .D(S_0_F_N5), .CK(CLK), .Q(S_0_q3[0]), .QN() );
  DFF_X1 S_0_F_out3_reg_1_ ( .D(S_0_F_N2), .CK(CLK), .Q(S_0_q3[1]), .QN() );
  DFF_X1 S_0_F_out1_reg_0_ ( .D(S_0_F_N3), .CK(CLK), .Q(S_0_q1[0]), .QN() );
  DFF_X1 S_0_F_out1_reg_1_ ( .D(S_0_F_N0), .CK(CLK), .Q(S_0_q1[1]), .QN() );
  NOR2_X1 S_0_F_Inst_0__CF_Inst_U2 ( .A1(S_0_F_in1[2]), .A2(
        S_0_F_Inst_0__CF_Inst_n3), .ZN(S_0_F_CF_Out[0]) );
  INV_X1 S_0_F_Inst_0__CF_Inst_U1 ( .A(S_0_F_in1[3]), .ZN(
        S_0_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_0_F_Inst_1__CF_Inst_U2 ( .A(S_0_F_Inst_1__CF_Inst_n3), .B(
        S_0_F_in1[1]), .ZN(S_0_F_CF_Out[1]) );
  NAND2_X1 S_0_F_Inst_1__CF_Inst_U1 ( .A1(S_0_F_in2[2]), .A2(S_0_F_in1[3]), 
        .ZN(S_0_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_0_F_Inst_2__CF_Inst_U1 ( .A1(S_0_F_in1[3]), .A2(S_0_F_in3[2]), .ZN(
        S_0_F_CF_Out[2]) );
  NOR2_X1 S_0_F_Inst_3__CF_Inst_U2 ( .A1(S_0_F_in2[3]), .A2(
        S_0_F_Inst_3__CF_Inst_n3), .ZN(S_0_F_CF_Out[3]) );
  INV_X1 S_0_F_Inst_3__CF_Inst_U1 ( .A(S_0_F_in1[2]), .ZN(
        S_0_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_0_F_Inst_4__CF_Inst_U2 ( .A(S_0_F_Inst_4__CF_Inst_n3), .B(
        S_0_F_in2[1]), .ZN(S_0_F_CF_Out[4]) );
  NAND2_X1 S_0_F_Inst_4__CF_Inst_U1 ( .A1(S_0_F_in2[2]), .A2(S_0_F_in2[3]), 
        .ZN(S_0_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_0_F_Inst_5__CF_Inst_U1 ( .A1(S_0_F_in3[2]), .A2(S_0_F_in2[3]), 
        .ZN(S_0_F_CF_Out[5]) );
  XNOR2_X1 S_0_F_Inst_6__CF_Inst_U2 ( .A(S_0_F_Inst_6__CF_Inst_n7), .B(
        S_0_F_in3[1]), .ZN(S_0_F_CF_Out[6]) );
  NOR2_X1 S_0_F_Inst_6__CF_Inst_U1 ( .A1(S_0_F_in1[2]), .A2(S_0_F_in3[3]), 
        .ZN(S_0_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_0_F_Inst_7__CF_Inst_U1 ( .A1(S_0_F_in2[2]), .A2(S_0_F_in3[3]), 
        .ZN(S_0_F_CF_Out[7]) );
  OR2_X1 S_0_F_Inst_8__CF_Inst_U1 ( .A1(S_0_F_in3[3]), .A2(S_0_F_in3[2]), .ZN(
        S_0_F_CF_Out[8]) );
  NOR2_X1 S_0_F_Inst_9__CF_Inst_U2 ( .A1(S_0_F_in1[3]), .A2(
        S_0_F_Inst_9__CF_Inst_n3), .ZN(S_0_F_CF_Out[9]) );
  INV_X1 S_0_F_Inst_9__CF_Inst_U1 ( .A(S_0_F_in1[1]), .ZN(
        S_0_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_0_F_Inst_10__CF_Inst_U1 ( .A1(S_0_F_in2[1]), .A2(S_0_F_in1[3]), 
        .ZN(S_0_F_CF_Out[10]) );
  XNOR2_X1 S_0_F_Inst_11__CF_Inst_U2 ( .A(S_0_F_Inst_11__CF_Inst_n3), .B(
        S_0_F_in1[0]), .ZN(S_0_F_CF_Out[11]) );
  NAND2_X1 S_0_F_Inst_11__CF_Inst_U1 ( .A1(S_0_F_in3[1]), .A2(S_0_F_in1[3]), 
        .ZN(S_0_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_0_F_Inst_12__CF_Inst_U2 ( .A(S_0_F_Inst_12__CF_Inst_n3), .B(
        S_0_F_in2[0]), .ZN(S_0_F_CF_Out[12]) );
  NAND2_X1 S_0_F_Inst_12__CF_Inst_U1 ( .A1(S_0_F_in1[1]), .A2(S_0_F_in2[3]), 
        .ZN(S_0_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_0_F_Inst_13__CF_Inst_U2 ( .A1(S_0_F_in2[3]), .A2(
        S_0_F_Inst_13__CF_Inst_n3), .ZN(S_0_F_CF_Out[13]) );
  INV_X1 S_0_F_Inst_13__CF_Inst_U1 ( .A(S_0_F_in2[1]), .ZN(
        S_0_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_0_F_Inst_14__CF_Inst_U1 ( .A1(S_0_F_in3[1]), .A2(S_0_F_in2[3]), 
        .ZN(S_0_F_CF_Out[14]) );
  XNOR2_X1 S_0_F_Inst_15__CF_Inst_U2 ( .A(S_0_F_Inst_15__CF_Inst_n7), .B(
        S_0_F_in3[0]), .ZN(S_0_F_CF_Out[15]) );
  NOR2_X1 S_0_F_Inst_15__CF_Inst_U1 ( .A1(S_0_F_in1[1]), .A2(S_0_F_in3[3]), 
        .ZN(S_0_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_0_F_Inst_16__CF_Inst_U2 ( .A1(S_0_F_in3[3]), .A2(
        S_0_F_Inst_16__CF_Inst_n3), .ZN(S_0_F_CF_Out[16]) );
  INV_X1 S_0_F_Inst_16__CF_Inst_U1 ( .A(S_0_F_in2[1]), .ZN(
        S_0_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_0_F_Inst_17__CF_Inst_U2 ( .A1(S_0_F_in3[1]), .A2(
        S_0_F_Inst_17__CF_Inst_n3), .ZN(S_0_F_CF_Out[17]) );
  INV_X1 S_0_F_Inst_17__CF_Inst_U1 ( .A(S_0_F_in3[3]), .ZN(
        S_0_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_0_F_InstXOR_0__Compression1_U2 ( .A(
        S_0_F_InstXOR_0__Compression1_n3), .B(S_0_F_CF_Reg[2]), .ZN(
        S_0_F_q1[2]) );
  XNOR2_X1 S_0_F_InstXOR_0__Compression1_U1 ( .A(S_0_F_CF_Reg[0]), .B(
        S_0_F_CF_Reg[1]), .ZN(S_0_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_0_F_InstXOR_0__Compression2_U2 ( .A(
        S_0_F_InstXOR_0__Compression2_n3), .B(S_0_F_CF_Reg[5]), .ZN(
        S_0_F_q2[2]) );
  XNOR2_X1 S_0_F_InstXOR_0__Compression2_U1 ( .A(S_0_F_CF_Reg[3]), .B(
        S_0_F_CF_Reg[4]), .ZN(S_0_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_0_F_InstXOR_0__Compression3_U2 ( .A(
        S_0_F_InstXOR_0__Compression3_n3), .B(S_0_F_CF_Reg[8]), .ZN(
        S_0_F_q3[2]) );
  XNOR2_X1 S_0_F_InstXOR_0__Compression3_U1 ( .A(S_0_F_CF_Reg[6]), .B(
        S_0_F_CF_Reg[7]), .ZN(S_0_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_0_F_InstXOR_1__Compression1_U2 ( .A(
        S_0_F_InstXOR_1__Compression1_n3), .B(S_0_F_CF_Reg[11]), .ZN(
        S_0_F_q1[3]) );
  XNOR2_X1 S_0_F_InstXOR_1__Compression1_U1 ( .A(S_0_F_CF_Reg[9]), .B(
        S_0_F_CF_Reg[10]), .ZN(S_0_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_0_F_InstXOR_1__Compression2_U2 ( .A(
        S_0_F_InstXOR_1__Compression2_n3), .B(S_0_F_CF_Reg[14]), .ZN(
        S_0_F_q2[3]) );
  XNOR2_X1 S_0_F_InstXOR_1__Compression2_U1 ( .A(S_0_F_CF_Reg[12]), .B(
        S_0_F_CF_Reg[13]), .ZN(S_0_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_0_F_InstXOR_1__Compression3_U2 ( .A(
        S_0_F_InstXOR_1__Compression3_n3), .B(S_0_F_CF_Reg[17]), .ZN(
        S_0_F_q3[3]) );
  XNOR2_X1 S_0_F_InstXOR_1__Compression3_U1 ( .A(S_0_F_CF_Reg[15]), .B(
        S_0_F_CF_Reg[16]), .ZN(S_0_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_0_G_CF_Reg_reg_0_ ( .D(S_0_G_CF_Out[0]), .CK(CLK), .Q(
        S_0_G_CF_Reg[0]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_1_ ( .D(S_0_G_CF_Out[1]), .CK(CLK), .Q(
        S_0_G_CF_Reg[1]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_2_ ( .D(S_0_G_CF_Out[2]), .CK(CLK), .Q(
        S_0_G_CF_Reg[2]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_3_ ( .D(S_0_G_CF_Out[3]), .CK(CLK), .Q(
        S_0_G_CF_Reg[3]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_4_ ( .D(S_0_G_CF_Out[4]), .CK(CLK), .Q(
        S_0_G_CF_Reg[4]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_5_ ( .D(S_0_G_CF_Out[5]), .CK(CLK), .Q(
        S_0_G_CF_Reg[5]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_6_ ( .D(S_0_G_CF_Out[6]), .CK(CLK), .Q(
        S_0_G_CF_Reg[6]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_7_ ( .D(S_0_G_CF_Out[7]), .CK(CLK), .Q(
        S_0_G_CF_Reg[7]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_8_ ( .D(S_0_G_CF_Out[8]), .CK(CLK), .Q(
        S_0_G_CF_Reg[8]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_9_ ( .D(S_0_G_CF_Out[9]), .CK(CLK), .Q(
        S_0_G_CF_Reg[9]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_10_ ( .D(S_0_G_CF_Out[10]), .CK(CLK), .Q(
        S_0_G_CF_Reg[10]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_11_ ( .D(S_0_G_CF_Out[11]), .CK(CLK), .Q(
        S_0_G_CF_Reg[11]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_12_ ( .D(S_0_G_CF_Out[12]), .CK(CLK), .Q(
        S_0_G_CF_Reg[12]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_13_ ( .D(S_0_G_CF_Out[13]), .CK(CLK), .Q(
        S_0_G_CF_Reg[13]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_14_ ( .D(S_0_G_CF_Out[14]), .CK(CLK), .Q(
        S_0_G_CF_Reg[14]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_15_ ( .D(S_0_G_CF_Out[15]), .CK(CLK), .Q(
        S_0_G_CF_Reg[15]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_16_ ( .D(S_0_G_CF_Out[16]), .CK(CLK), .Q(
        S_0_G_CF_Reg[16]), .QN() );
  DFF_X1 S_0_G_CF_Reg_reg_17_ ( .D(S_0_G_CF_Out[17]), .CK(CLK), .Q(
        S_0_G_CF_Reg[17]), .QN() );
  DFF_X1 S_0_G_out1_reg_2_ ( .D(S_0_Rq1[2]), .CK(CLK), .Q(S_0_G_out1[2]), 
        .QN() );
  DFF_X1 S_0_G_out1_reg_3_ ( .D(S_0_Rq1[3]), .CK(CLK), .Q(S_0_G_out1[3]), 
        .QN() );
  DFF_X1 S_0_G_out2_reg_2_ ( .D(S_0_Rq2[2]), .CK(CLK), .Q(RF2_SHIFTROWS[6]), 
        .QN() );
  DFF_X1 S_0_G_out2_reg_3_ ( .D(S_0_Rq2[3]), .CK(CLK), .Q(RF2_SHIFTROWS[7]), 
        .QN() );
  DFF_X1 S_0_G_out3_reg_2_ ( .D(S_0_Rq3[2]), .CK(CLK), .Q(RF3_SHIFTROWS[6]), 
        .QN() );
  DFF_X1 S_0_G_out3_reg_3_ ( .D(S_0_Rq3[3]), .CK(CLK), .Q(RF3_SHIFTROWS[7]), 
        .QN() );
  AND2_X1 S_0_G_Inst_0__CF_Inst_U1 ( .A1(S_0_Rq1[1]), .A2(S_0_Rq1[3]), .ZN(
        S_0_G_CF_Out[0]) );
  NOR2_X1 S_0_G_Inst_1__CF_Inst_U2 ( .A1(S_0_Rq1[3]), .A2(
        S_0_G_Inst_1__CF_Inst_n3), .ZN(S_0_G_CF_Out[1]) );
  INV_X1 S_0_G_Inst_1__CF_Inst_U1 ( .A(S_0_Rq2[1]), .ZN(
        S_0_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_0_G_Inst_2__CF_Inst_U2 ( .A(S_0_G_Inst_2__CF_Inst_n3), .B(
        S_0_Rq2[0]), .ZN(S_0_G_CF_Out[2]) );
  NAND2_X1 S_0_G_Inst_2__CF_Inst_U1 ( .A1(S_0_Rq1[1]), .A2(S_0_Rq2[3]), .ZN(
        S_0_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_0_G_Inst_3__CF_Inst_U3 ( .A(S_0_Rq1[0]), .B(
        S_0_G_Inst_3__CF_Inst_n6), .ZN(S_0_G_CF_Out[3]) );
  NAND2_X1 S_0_G_Inst_3__CF_Inst_U2 ( .A1(S_0_Rq3[1]), .A2(
        S_0_G_Inst_3__CF_Inst_n5), .ZN(S_0_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_0_G_Inst_3__CF_Inst_U1 ( .A(S_0_Rq1[3]), .ZN(
        S_0_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_0_G_Inst_4__CF_Inst_U1 ( .A1(S_0_Rq2[1]), .A2(S_0_Rq2[3]), .ZN(
        S_0_G_CF_Out[4]) );
  OR2_X1 S_0_G_Inst_5__CF_Inst_U1 ( .A1(S_0_Rq3[3]), .A2(S_0_Rq2[1]), .ZN(
        S_0_G_CF_Out[5]) );
  AND2_X1 S_0_G_Inst_6__CF_Inst_U1 ( .A1(S_0_Rq3[1]), .A2(S_0_Rq2[3]), .ZN(
        S_0_G_CF_Out[6]) );
  XNOR2_X1 S_0_G_Inst_7__CF_Inst_U2 ( .A(S_0_G_Inst_7__CF_Inst_n3), .B(
        S_0_Rq3[0]), .ZN(S_0_G_CF_Out[7]) );
  NAND2_X1 S_0_G_Inst_7__CF_Inst_U1 ( .A1(S_0_Rq1[1]), .A2(S_0_Rq3[3]), .ZN(
        S_0_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_0_G_Inst_8__CF_Inst_U1 ( .A1(S_0_Rq3[3]), .A2(S_0_Rq3[1]), .ZN(
        S_0_G_CF_Out[8]) );
  NOR2_X1 S_0_G_Inst_9__CF_Inst_U2 ( .A1(S_0_Rq1[3]), .A2(
        S_0_G_Inst_9__CF_Inst_n3), .ZN(S_0_G_CF_Out[9]) );
  INV_X1 S_0_G_Inst_9__CF_Inst_U1 ( .A(S_0_Rq1[2]), .ZN(
        S_0_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_0_G_Inst_10__CF_Inst_U2 ( .A1(S_0_Rq2[2]), .A2(
        S_0_G_Inst_10__CF_Inst_n3), .ZN(S_0_G_CF_Out[10]) );
  INV_X1 S_0_G_Inst_10__CF_Inst_U1 ( .A(S_0_Rq1[3]), .ZN(
        S_0_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_0_G_Inst_11__CF_Inst_U3 ( .A(S_0_Rq1[1]), .B(
        S_0_G_Inst_11__CF_Inst_n6), .ZN(S_0_G_CF_Out[11]) );
  NAND2_X1 S_0_G_Inst_11__CF_Inst_U2 ( .A1(S_0_Rq1[3]), .A2(
        S_0_G_Inst_11__CF_Inst_n5), .ZN(S_0_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_0_G_Inst_11__CF_Inst_U1 ( .A(S_0_Rq3[2]), .ZN(
        S_0_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_0_G_Inst_12__CF_Inst_U2 ( .A1(S_0_Rq2[3]), .A2(
        S_0_G_Inst_12__CF_Inst_n3), .ZN(S_0_G_CF_Out[12]) );
  INV_X1 S_0_G_Inst_12__CF_Inst_U1 ( .A(S_0_Rq1[2]), .ZN(
        S_0_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_0_G_Inst_13__CF_Inst_U1 ( .A1(S_0_Rq2[2]), .A2(S_0_Rq2[3]), .ZN(
        S_0_G_CF_Out[13]) );
  XNOR2_X1 S_0_G_Inst_14__CF_Inst_U3 ( .A(S_0_Rq2[1]), .B(
        S_0_G_Inst_14__CF_Inst_n6), .ZN(S_0_G_CF_Out[14]) );
  NAND2_X1 S_0_G_Inst_14__CF_Inst_U2 ( .A1(S_0_Rq3[2]), .A2(
        S_0_G_Inst_14__CF_Inst_n5), .ZN(S_0_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_0_G_Inst_14__CF_Inst_U1 ( .A(S_0_Rq2[3]), .ZN(
        S_0_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_0_G_Inst_15__CF_Inst_U2 ( .A(S_0_G_Inst_15__CF_Inst_n3), .B(
        S_0_Rq3[1]), .ZN(S_0_G_CF_Out[15]) );
  NAND2_X1 S_0_G_Inst_15__CF_Inst_U1 ( .A1(S_0_Rq1[2]), .A2(S_0_Rq3[3]), .ZN(
        S_0_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_0_G_Inst_16__CF_Inst_U1 ( .A1(S_0_Rq2[2]), .A2(S_0_Rq3[3]), .ZN(
        S_0_G_CF_Out[16]) );
  NOR2_X1 S_0_G_Inst_17__CF_Inst_U2 ( .A1(S_0_Rq3[3]), .A2(
        S_0_G_Inst_17__CF_Inst_n3), .ZN(S_0_G_CF_Out[17]) );
  INV_X1 S_0_G_Inst_17__CF_Inst_U1 ( .A(S_0_Rq3[2]), .ZN(
        S_0_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_0_G_InstXOR_0__Compression1_U2 ( .A(
        S_0_G_InstXOR_0__Compression1_n3), .B(S_0_G_CF_Reg[2]), .ZN(
        S_0_G_out1[0]) );
  XNOR2_X1 S_0_G_InstXOR_0__Compression1_U1 ( .A(S_0_G_CF_Reg[0]), .B(
        S_0_G_CF_Reg[1]), .ZN(S_0_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_0_G_InstXOR_0__Compression2_U2 ( .A(
        S_0_G_InstXOR_0__Compression2_n3), .B(S_0_G_CF_Reg[5]), .ZN(
        RF2_SHIFTROWS[5]) );
  XNOR2_X1 S_0_G_InstXOR_0__Compression2_U1 ( .A(S_0_G_CF_Reg[3]), .B(
        S_0_G_CF_Reg[4]), .ZN(S_0_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_0_G_InstXOR_0__Compression3_U2 ( .A(
        S_0_G_InstXOR_0__Compression3_n3), .B(S_0_G_CF_Reg[8]), .ZN(
        RF3_SHIFTROWS[5]) );
  XNOR2_X1 S_0_G_InstXOR_0__Compression3_U1 ( .A(S_0_G_CF_Reg[6]), .B(
        S_0_G_CF_Reg[7]), .ZN(S_0_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_0_G_InstXOR_1__Compression1_U2 ( .A(
        S_0_G_InstXOR_1__Compression1_n3), .B(S_0_G_CF_Reg[11]), .ZN(
        S_0_G_out1[1]) );
  XNOR2_X1 S_0_G_InstXOR_1__Compression1_U1 ( .A(S_0_G_CF_Reg[9]), .B(
        S_0_G_CF_Reg[10]), .ZN(S_0_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_0_G_InstXOR_1__Compression2_U2 ( .A(
        S_0_G_InstXOR_1__Compression2_n3), .B(S_0_G_CF_Reg[14]), .ZN(
        RF2_SHIFTROWS[4]) );
  XNOR2_X1 S_0_G_InstXOR_1__Compression2_U1 ( .A(S_0_G_CF_Reg[12]), .B(
        S_0_G_CF_Reg[13]), .ZN(S_0_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_0_G_InstXOR_1__Compression3_U2 ( .A(
        S_0_G_InstXOR_1__Compression3_n3), .B(S_0_G_CF_Reg[17]), .ZN(
        RF3_SHIFTROWS[4]) );
  XNOR2_X1 S_0_G_InstXOR_1__Compression3_U1 ( .A(S_0_G_CF_Reg[15]), .B(
        S_0_G_CF_Reg[16]), .ZN(S_0_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_0_OutputAffine_U4 ( .A(S_0_G_out1[3]), .ZN(RF1_SHIFTROWS[7]) );
  INV_X1 S_0_OutputAffine_U3 ( .A(S_0_G_out1[2]), .ZN(RF1_SHIFTROWS[6]) );
  INV_X1 S_0_OutputAffine_U2 ( .A(S_0_G_out1[1]), .ZN(RF1_SHIFTROWS[4]) );
  INV_X1 S_0_OutputAffine_U1 ( .A(S_0_G_out1[0]), .ZN(RF1_SHIFTROWS[5]) );
  DFF_X1 S_1_Rq3_reg_0_ ( .D(S_1_q3[0]), .CK(CLK), .Q(S_1_Rq3[0]), .QN() );
  DFF_X1 S_1_Rq3_reg_1_ ( .D(S_1_q3[1]), .CK(CLK), .Q(S_1_Rq3[1]), .QN() );
  DFF_X1 S_1_Rq3_reg_2_ ( .D(S_1_q3[2]), .CK(CLK), .Q(S_1_Rq3[2]), .QN() );
  DFF_X1 S_1_Rq3_reg_3_ ( .D(S_1_q3[3]), .CK(CLK), .Q(S_1_Rq3[3]), .QN() );
  DFF_X1 S_1_Rq2_reg_0_ ( .D(S_1_q2[0]), .CK(CLK), .Q(S_1_Rq2[0]), .QN() );
  DFF_X1 S_1_Rq2_reg_1_ ( .D(S_1_q2[1]), .CK(CLK), .Q(S_1_Rq2[1]), .QN() );
  DFF_X1 S_1_Rq2_reg_2_ ( .D(S_1_q2[2]), .CK(CLK), .Q(S_1_Rq2[2]), .QN() );
  DFF_X1 S_1_Rq2_reg_3_ ( .D(S_1_q2[3]), .CK(CLK), .Q(S_1_Rq2[3]), .QN() );
  DFF_X1 S_1_Rq1_reg_0_ ( .D(S_1_q1[0]), .CK(CLK), .Q(S_1_Rq1[0]), .QN() );
  DFF_X1 S_1_Rq1_reg_1_ ( .D(S_1_q1[1]), .CK(CLK), .Q(S_1_Rq1[1]), .QN() );
  DFF_X1 S_1_Rq1_reg_2_ ( .D(S_1_q1[2]), .CK(CLK), .Q(S_1_Rq1[2]), .QN() );
  DFF_X1 S_1_Rq1_reg_3_ ( .D(S_1_q1[3]), .CK(CLK), .Q(S_1_Rq1[3]), .QN() );
  INV_X1 S_1_InputAffine_U4 ( .A(SUB_IN1[4]), .ZN(S_1_F_in1[0]) );
  INV_X1 S_1_InputAffine_U3 ( .A(SUB_IN1[6]), .ZN(S_1_F_in1[3]) );
  INV_X1 S_1_InputAffine_U2 ( .A(SUB_IN1[7]), .ZN(S_1_F_in1[1]) );
  INV_X1 S_1_InputAffine_U1 ( .A(SUB_IN1[5]), .ZN(S_1_F_in1[2]) );
  XNOR2_X1 S_1_F_U18 ( .A(S_1_F_n12), .B(FRESH[11]), .ZN(S_1_q3[3]) );
  XNOR2_X1 S_1_F_U17 ( .A(FRESH[10]), .B(S_1_F_q3[3]), .ZN(S_1_F_n12) );
  XNOR2_X1 S_1_F_U16 ( .A(S_1_F_n11), .B(FRESH[9]), .ZN(S_1_q3[2]) );
  XNOR2_X1 S_1_F_U15 ( .A(FRESH[8]), .B(S_1_F_q3[2]), .ZN(S_1_F_n11) );
  XOR2_X1 S_1_F_U14 ( .A(FRESH[11]), .B(S_1_F_q2[3]), .Z(S_1_q2[3]) );
  XOR2_X1 S_1_F_U13 ( .A(FRESH[9]), .B(S_1_F_q2[2]), .Z(S_1_q2[2]) );
  XOR2_X1 S_1_F_U12 ( .A(FRESH[10]), .B(S_1_F_q1[3]), .Z(S_1_q1[3]) );
  XOR2_X1 S_1_F_U11 ( .A(FRESH[8]), .B(S_1_F_q1[2]), .Z(S_1_q1[2]) );
  XNOR2_X1 S_1_F_U10 ( .A(S_1_F_n10), .B(FRESH[13]), .ZN(S_1_F_N5) );
  XNOR2_X1 S_1_F_U9 ( .A(S_1_F_in3[3]), .B(FRESH[12]), .ZN(S_1_F_n10) );
  XOR2_X1 S_1_F_U8 ( .A(FRESH[13]), .B(S_1_F_in2[3]), .Z(S_1_F_N4) );
  XOR2_X1 S_1_F_U7 ( .A(FRESH[12]), .B(S_1_F_in1[3]), .Z(S_1_F_N3) );
  XNOR2_X1 S_1_F_U6 ( .A(S_1_F_n9), .B(FRESH[15]), .ZN(S_1_F_N2) );
  XNOR2_X1 S_1_F_U5 ( .A(S_1_F_in3[2]), .B(FRESH[14]), .ZN(S_1_F_n9) );
  XOR2_X1 S_1_F_U4 ( .A(FRESH[15]), .B(S_1_F_in2[2]), .Z(S_1_F_N1) );
  XOR2_X1 S_1_F_U3 ( .A(FRESH[14]), .B(S_1_F_in1[2]), .Z(S_1_F_N0) );
  DFF_X1 S_1_F_CF_Reg_reg_0_ ( .D(S_1_F_CF_Out[0]), .CK(CLK), .Q(
        S_1_F_CF_Reg[0]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_1_ ( .D(S_1_F_CF_Out[1]), .CK(CLK), .Q(
        S_1_F_CF_Reg[1]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_2_ ( .D(S_1_F_CF_Out[2]), .CK(CLK), .Q(
        S_1_F_CF_Reg[2]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_3_ ( .D(S_1_F_CF_Out[3]), .CK(CLK), .Q(
        S_1_F_CF_Reg[3]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_4_ ( .D(S_1_F_CF_Out[4]), .CK(CLK), .Q(
        S_1_F_CF_Reg[4]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_5_ ( .D(S_1_F_CF_Out[5]), .CK(CLK), .Q(
        S_1_F_CF_Reg[5]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_6_ ( .D(S_1_F_CF_Out[6]), .CK(CLK), .Q(
        S_1_F_CF_Reg[6]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_7_ ( .D(S_1_F_CF_Out[7]), .CK(CLK), .Q(
        S_1_F_CF_Reg[7]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_8_ ( .D(S_1_F_CF_Out[8]), .CK(CLK), .Q(
        S_1_F_CF_Reg[8]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_9_ ( .D(S_1_F_CF_Out[9]), .CK(CLK), .Q(
        S_1_F_CF_Reg[9]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_10_ ( .D(S_1_F_CF_Out[10]), .CK(CLK), .Q(
        S_1_F_CF_Reg[10]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_11_ ( .D(S_1_F_CF_Out[11]), .CK(CLK), .Q(
        S_1_F_CF_Reg[11]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_12_ ( .D(S_1_F_CF_Out[12]), .CK(CLK), .Q(
        S_1_F_CF_Reg[12]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_13_ ( .D(S_1_F_CF_Out[13]), .CK(CLK), .Q(
        S_1_F_CF_Reg[13]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_14_ ( .D(S_1_F_CF_Out[14]), .CK(CLK), .Q(
        S_1_F_CF_Reg[14]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_15_ ( .D(S_1_F_CF_Out[15]), .CK(CLK), .Q(
        S_1_F_CF_Reg[15]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_16_ ( .D(S_1_F_CF_Out[16]), .CK(CLK), .Q(
        S_1_F_CF_Reg[16]), .QN() );
  DFF_X1 S_1_F_CF_Reg_reg_17_ ( .D(S_1_F_CF_Out[17]), .CK(CLK), .Q(
        S_1_F_CF_Reg[17]), .QN() );
  DFF_X1 S_1_F_out2_reg_0_ ( .D(S_1_F_N4), .CK(CLK), .Q(S_1_q2[0]), .QN() );
  DFF_X1 S_1_F_out2_reg_1_ ( .D(S_1_F_N1), .CK(CLK), .Q(S_1_q2[1]), .QN() );
  DFF_X1 S_1_F_out3_reg_0_ ( .D(S_1_F_N5), .CK(CLK), .Q(S_1_q3[0]), .QN() );
  DFF_X1 S_1_F_out3_reg_1_ ( .D(S_1_F_N2), .CK(CLK), .Q(S_1_q3[1]), .QN() );
  DFF_X1 S_1_F_out1_reg_0_ ( .D(S_1_F_N3), .CK(CLK), .Q(S_1_q1[0]), .QN() );
  DFF_X1 S_1_F_out1_reg_1_ ( .D(S_1_F_N0), .CK(CLK), .Q(S_1_q1[1]), .QN() );
  NOR2_X1 S_1_F_Inst_0__CF_Inst_U2 ( .A1(S_1_F_in1[2]), .A2(
        S_1_F_Inst_0__CF_Inst_n3), .ZN(S_1_F_CF_Out[0]) );
  INV_X1 S_1_F_Inst_0__CF_Inst_U1 ( .A(S_1_F_in1[3]), .ZN(
        S_1_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_1_F_Inst_1__CF_Inst_U2 ( .A(S_1_F_Inst_1__CF_Inst_n3), .B(
        S_1_F_in1[1]), .ZN(S_1_F_CF_Out[1]) );
  NAND2_X1 S_1_F_Inst_1__CF_Inst_U1 ( .A1(S_1_F_in2[2]), .A2(S_1_F_in1[3]), 
        .ZN(S_1_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_1_F_Inst_2__CF_Inst_U1 ( .A1(S_1_F_in1[3]), .A2(S_1_F_in3[2]), .ZN(
        S_1_F_CF_Out[2]) );
  NOR2_X1 S_1_F_Inst_3__CF_Inst_U2 ( .A1(S_1_F_in2[3]), .A2(
        S_1_F_Inst_3__CF_Inst_n3), .ZN(S_1_F_CF_Out[3]) );
  INV_X1 S_1_F_Inst_3__CF_Inst_U1 ( .A(S_1_F_in1[2]), .ZN(
        S_1_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_1_F_Inst_4__CF_Inst_U2 ( .A(S_1_F_Inst_4__CF_Inst_n3), .B(
        S_1_F_in2[1]), .ZN(S_1_F_CF_Out[4]) );
  NAND2_X1 S_1_F_Inst_4__CF_Inst_U1 ( .A1(S_1_F_in2[2]), .A2(S_1_F_in2[3]), 
        .ZN(S_1_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_1_F_Inst_5__CF_Inst_U1 ( .A1(S_1_F_in3[2]), .A2(S_1_F_in2[3]), 
        .ZN(S_1_F_CF_Out[5]) );
  XNOR2_X1 S_1_F_Inst_6__CF_Inst_U2 ( .A(S_1_F_Inst_6__CF_Inst_n7), .B(
        S_1_F_in3[1]), .ZN(S_1_F_CF_Out[6]) );
  NOR2_X1 S_1_F_Inst_6__CF_Inst_U1 ( .A1(S_1_F_in1[2]), .A2(S_1_F_in3[3]), 
        .ZN(S_1_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_1_F_Inst_7__CF_Inst_U1 ( .A1(S_1_F_in2[2]), .A2(S_1_F_in3[3]), 
        .ZN(S_1_F_CF_Out[7]) );
  OR2_X1 S_1_F_Inst_8__CF_Inst_U1 ( .A1(S_1_F_in3[3]), .A2(S_1_F_in3[2]), .ZN(
        S_1_F_CF_Out[8]) );
  NOR2_X1 S_1_F_Inst_9__CF_Inst_U2 ( .A1(S_1_F_in1[3]), .A2(
        S_1_F_Inst_9__CF_Inst_n3), .ZN(S_1_F_CF_Out[9]) );
  INV_X1 S_1_F_Inst_9__CF_Inst_U1 ( .A(S_1_F_in1[1]), .ZN(
        S_1_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_1_F_Inst_10__CF_Inst_U1 ( .A1(S_1_F_in2[1]), .A2(S_1_F_in1[3]), 
        .ZN(S_1_F_CF_Out[10]) );
  XNOR2_X1 S_1_F_Inst_11__CF_Inst_U2 ( .A(S_1_F_Inst_11__CF_Inst_n3), .B(
        S_1_F_in1[0]), .ZN(S_1_F_CF_Out[11]) );
  NAND2_X1 S_1_F_Inst_11__CF_Inst_U1 ( .A1(S_1_F_in3[1]), .A2(S_1_F_in1[3]), 
        .ZN(S_1_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_1_F_Inst_12__CF_Inst_U2 ( .A(S_1_F_Inst_12__CF_Inst_n3), .B(
        S_1_F_in2[0]), .ZN(S_1_F_CF_Out[12]) );
  NAND2_X1 S_1_F_Inst_12__CF_Inst_U1 ( .A1(S_1_F_in1[1]), .A2(S_1_F_in2[3]), 
        .ZN(S_1_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_1_F_Inst_13__CF_Inst_U2 ( .A1(S_1_F_in2[3]), .A2(
        S_1_F_Inst_13__CF_Inst_n3), .ZN(S_1_F_CF_Out[13]) );
  INV_X1 S_1_F_Inst_13__CF_Inst_U1 ( .A(S_1_F_in2[1]), .ZN(
        S_1_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_1_F_Inst_14__CF_Inst_U1 ( .A1(S_1_F_in3[1]), .A2(S_1_F_in2[3]), 
        .ZN(S_1_F_CF_Out[14]) );
  XNOR2_X1 S_1_F_Inst_15__CF_Inst_U2 ( .A(S_1_F_Inst_15__CF_Inst_n7), .B(
        S_1_F_in3[0]), .ZN(S_1_F_CF_Out[15]) );
  NOR2_X1 S_1_F_Inst_15__CF_Inst_U1 ( .A1(S_1_F_in1[1]), .A2(S_1_F_in3[3]), 
        .ZN(S_1_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_1_F_Inst_16__CF_Inst_U2 ( .A1(S_1_F_in3[3]), .A2(
        S_1_F_Inst_16__CF_Inst_n3), .ZN(S_1_F_CF_Out[16]) );
  INV_X1 S_1_F_Inst_16__CF_Inst_U1 ( .A(S_1_F_in2[1]), .ZN(
        S_1_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_1_F_Inst_17__CF_Inst_U2 ( .A1(S_1_F_in3[1]), .A2(
        S_1_F_Inst_17__CF_Inst_n3), .ZN(S_1_F_CF_Out[17]) );
  INV_X1 S_1_F_Inst_17__CF_Inst_U1 ( .A(S_1_F_in3[3]), .ZN(
        S_1_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_1_F_InstXOR_0__Compression1_U2 ( .A(
        S_1_F_InstXOR_0__Compression1_n3), .B(S_1_F_CF_Reg[2]), .ZN(
        S_1_F_q1[2]) );
  XNOR2_X1 S_1_F_InstXOR_0__Compression1_U1 ( .A(S_1_F_CF_Reg[0]), .B(
        S_1_F_CF_Reg[1]), .ZN(S_1_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_1_F_InstXOR_0__Compression2_U2 ( .A(
        S_1_F_InstXOR_0__Compression2_n3), .B(S_1_F_CF_Reg[5]), .ZN(
        S_1_F_q2[2]) );
  XNOR2_X1 S_1_F_InstXOR_0__Compression2_U1 ( .A(S_1_F_CF_Reg[3]), .B(
        S_1_F_CF_Reg[4]), .ZN(S_1_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_1_F_InstXOR_0__Compression3_U2 ( .A(
        S_1_F_InstXOR_0__Compression3_n3), .B(S_1_F_CF_Reg[8]), .ZN(
        S_1_F_q3[2]) );
  XNOR2_X1 S_1_F_InstXOR_0__Compression3_U1 ( .A(S_1_F_CF_Reg[6]), .B(
        S_1_F_CF_Reg[7]), .ZN(S_1_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_1_F_InstXOR_1__Compression1_U2 ( .A(
        S_1_F_InstXOR_1__Compression1_n3), .B(S_1_F_CF_Reg[11]), .ZN(
        S_1_F_q1[3]) );
  XNOR2_X1 S_1_F_InstXOR_1__Compression1_U1 ( .A(S_1_F_CF_Reg[9]), .B(
        S_1_F_CF_Reg[10]), .ZN(S_1_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_1_F_InstXOR_1__Compression2_U2 ( .A(
        S_1_F_InstXOR_1__Compression2_n3), .B(S_1_F_CF_Reg[14]), .ZN(
        S_1_F_q2[3]) );
  XNOR2_X1 S_1_F_InstXOR_1__Compression2_U1 ( .A(S_1_F_CF_Reg[12]), .B(
        S_1_F_CF_Reg[13]), .ZN(S_1_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_1_F_InstXOR_1__Compression3_U2 ( .A(
        S_1_F_InstXOR_1__Compression3_n3), .B(S_1_F_CF_Reg[17]), .ZN(
        S_1_F_q3[3]) );
  XNOR2_X1 S_1_F_InstXOR_1__Compression3_U1 ( .A(S_1_F_CF_Reg[15]), .B(
        S_1_F_CF_Reg[16]), .ZN(S_1_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_1_G_CF_Reg_reg_0_ ( .D(S_1_G_CF_Out[0]), .CK(CLK), .Q(
        S_1_G_CF_Reg[0]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_1_ ( .D(S_1_G_CF_Out[1]), .CK(CLK), .Q(
        S_1_G_CF_Reg[1]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_2_ ( .D(S_1_G_CF_Out[2]), .CK(CLK), .Q(
        S_1_G_CF_Reg[2]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_3_ ( .D(S_1_G_CF_Out[3]), .CK(CLK), .Q(
        S_1_G_CF_Reg[3]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_4_ ( .D(S_1_G_CF_Out[4]), .CK(CLK), .Q(
        S_1_G_CF_Reg[4]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_5_ ( .D(S_1_G_CF_Out[5]), .CK(CLK), .Q(
        S_1_G_CF_Reg[5]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_6_ ( .D(S_1_G_CF_Out[6]), .CK(CLK), .Q(
        S_1_G_CF_Reg[6]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_7_ ( .D(S_1_G_CF_Out[7]), .CK(CLK), .Q(
        S_1_G_CF_Reg[7]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_8_ ( .D(S_1_G_CF_Out[8]), .CK(CLK), .Q(
        S_1_G_CF_Reg[8]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_9_ ( .D(S_1_G_CF_Out[9]), .CK(CLK), .Q(
        S_1_G_CF_Reg[9]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_10_ ( .D(S_1_G_CF_Out[10]), .CK(CLK), .Q(
        S_1_G_CF_Reg[10]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_11_ ( .D(S_1_G_CF_Out[11]), .CK(CLK), .Q(
        S_1_G_CF_Reg[11]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_12_ ( .D(S_1_G_CF_Out[12]), .CK(CLK), .Q(
        S_1_G_CF_Reg[12]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_13_ ( .D(S_1_G_CF_Out[13]), .CK(CLK), .Q(
        S_1_G_CF_Reg[13]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_14_ ( .D(S_1_G_CF_Out[14]), .CK(CLK), .Q(
        S_1_G_CF_Reg[14]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_15_ ( .D(S_1_G_CF_Out[15]), .CK(CLK), .Q(
        S_1_G_CF_Reg[15]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_16_ ( .D(S_1_G_CF_Out[16]), .CK(CLK), .Q(
        S_1_G_CF_Reg[16]), .QN() );
  DFF_X1 S_1_G_CF_Reg_reg_17_ ( .D(S_1_G_CF_Out[17]), .CK(CLK), .Q(
        S_1_G_CF_Reg[17]), .QN() );
  DFF_X1 S_1_G_out1_reg_2_ ( .D(S_1_Rq1[2]), .CK(CLK), .Q(S_1_G_out1[2]), 
        .QN() );
  DFF_X1 S_1_G_out1_reg_3_ ( .D(S_1_Rq1[3]), .CK(CLK), .Q(S_1_G_out1[3]), 
        .QN() );
  DFF_X1 S_1_G_out2_reg_2_ ( .D(S_1_Rq2[2]), .CK(CLK), .Q(RF2_SHIFTROWS[10]), 
        .QN() );
  DFF_X1 S_1_G_out2_reg_3_ ( .D(S_1_Rq2[3]), .CK(CLK), .Q(RF2_SHIFTROWS[11]), 
        .QN() );
  DFF_X1 S_1_G_out3_reg_2_ ( .D(S_1_Rq3[2]), .CK(CLK), .Q(RF3_SHIFTROWS[10]), 
        .QN() );
  DFF_X1 S_1_G_out3_reg_3_ ( .D(S_1_Rq3[3]), .CK(CLK), .Q(RF3_SHIFTROWS[11]), 
        .QN() );
  AND2_X1 S_1_G_Inst_0__CF_Inst_U1 ( .A1(S_1_Rq1[1]), .A2(S_1_Rq1[3]), .ZN(
        S_1_G_CF_Out[0]) );
  NOR2_X1 S_1_G_Inst_1__CF_Inst_U2 ( .A1(S_1_Rq1[3]), .A2(
        S_1_G_Inst_1__CF_Inst_n3), .ZN(S_1_G_CF_Out[1]) );
  INV_X1 S_1_G_Inst_1__CF_Inst_U1 ( .A(S_1_Rq2[1]), .ZN(
        S_1_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_1_G_Inst_2__CF_Inst_U2 ( .A(S_1_G_Inst_2__CF_Inst_n3), .B(
        S_1_Rq2[0]), .ZN(S_1_G_CF_Out[2]) );
  NAND2_X1 S_1_G_Inst_2__CF_Inst_U1 ( .A1(S_1_Rq1[1]), .A2(S_1_Rq2[3]), .ZN(
        S_1_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_1_G_Inst_3__CF_Inst_U3 ( .A(S_1_Rq1[0]), .B(
        S_1_G_Inst_3__CF_Inst_n6), .ZN(S_1_G_CF_Out[3]) );
  NAND2_X1 S_1_G_Inst_3__CF_Inst_U2 ( .A1(S_1_Rq3[1]), .A2(
        S_1_G_Inst_3__CF_Inst_n5), .ZN(S_1_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_1_G_Inst_3__CF_Inst_U1 ( .A(S_1_Rq1[3]), .ZN(
        S_1_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_1_G_Inst_4__CF_Inst_U1 ( .A1(S_1_Rq2[1]), .A2(S_1_Rq2[3]), .ZN(
        S_1_G_CF_Out[4]) );
  OR2_X1 S_1_G_Inst_5__CF_Inst_U1 ( .A1(S_1_Rq3[3]), .A2(S_1_Rq2[1]), .ZN(
        S_1_G_CF_Out[5]) );
  AND2_X1 S_1_G_Inst_6__CF_Inst_U1 ( .A1(S_1_Rq3[1]), .A2(S_1_Rq2[3]), .ZN(
        S_1_G_CF_Out[6]) );
  XNOR2_X1 S_1_G_Inst_7__CF_Inst_U2 ( .A(S_1_G_Inst_7__CF_Inst_n3), .B(
        S_1_Rq3[0]), .ZN(S_1_G_CF_Out[7]) );
  NAND2_X1 S_1_G_Inst_7__CF_Inst_U1 ( .A1(S_1_Rq1[1]), .A2(S_1_Rq3[3]), .ZN(
        S_1_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_1_G_Inst_8__CF_Inst_U1 ( .A1(S_1_Rq3[3]), .A2(S_1_Rq3[1]), .ZN(
        S_1_G_CF_Out[8]) );
  NOR2_X1 S_1_G_Inst_9__CF_Inst_U2 ( .A1(S_1_Rq1[3]), .A2(
        S_1_G_Inst_9__CF_Inst_n3), .ZN(S_1_G_CF_Out[9]) );
  INV_X1 S_1_G_Inst_9__CF_Inst_U1 ( .A(S_1_Rq1[2]), .ZN(
        S_1_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_1_G_Inst_10__CF_Inst_U2 ( .A1(S_1_Rq2[2]), .A2(
        S_1_G_Inst_10__CF_Inst_n3), .ZN(S_1_G_CF_Out[10]) );
  INV_X1 S_1_G_Inst_10__CF_Inst_U1 ( .A(S_1_Rq1[3]), .ZN(
        S_1_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_1_G_Inst_11__CF_Inst_U3 ( .A(S_1_Rq1[1]), .B(
        S_1_G_Inst_11__CF_Inst_n6), .ZN(S_1_G_CF_Out[11]) );
  NAND2_X1 S_1_G_Inst_11__CF_Inst_U2 ( .A1(S_1_Rq1[3]), .A2(
        S_1_G_Inst_11__CF_Inst_n5), .ZN(S_1_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_1_G_Inst_11__CF_Inst_U1 ( .A(S_1_Rq3[2]), .ZN(
        S_1_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_1_G_Inst_12__CF_Inst_U2 ( .A1(S_1_Rq2[3]), .A2(
        S_1_G_Inst_12__CF_Inst_n3), .ZN(S_1_G_CF_Out[12]) );
  INV_X1 S_1_G_Inst_12__CF_Inst_U1 ( .A(S_1_Rq1[2]), .ZN(
        S_1_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_1_G_Inst_13__CF_Inst_U1 ( .A1(S_1_Rq2[2]), .A2(S_1_Rq2[3]), .ZN(
        S_1_G_CF_Out[13]) );
  XNOR2_X1 S_1_G_Inst_14__CF_Inst_U3 ( .A(S_1_Rq2[1]), .B(
        S_1_G_Inst_14__CF_Inst_n6), .ZN(S_1_G_CF_Out[14]) );
  NAND2_X1 S_1_G_Inst_14__CF_Inst_U2 ( .A1(S_1_Rq3[2]), .A2(
        S_1_G_Inst_14__CF_Inst_n5), .ZN(S_1_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_1_G_Inst_14__CF_Inst_U1 ( .A(S_1_Rq2[3]), .ZN(
        S_1_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_1_G_Inst_15__CF_Inst_U2 ( .A(S_1_G_Inst_15__CF_Inst_n3), .B(
        S_1_Rq3[1]), .ZN(S_1_G_CF_Out[15]) );
  NAND2_X1 S_1_G_Inst_15__CF_Inst_U1 ( .A1(S_1_Rq1[2]), .A2(S_1_Rq3[3]), .ZN(
        S_1_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_1_G_Inst_16__CF_Inst_U1 ( .A1(S_1_Rq2[2]), .A2(S_1_Rq3[3]), .ZN(
        S_1_G_CF_Out[16]) );
  NOR2_X1 S_1_G_Inst_17__CF_Inst_U2 ( .A1(S_1_Rq3[3]), .A2(
        S_1_G_Inst_17__CF_Inst_n3), .ZN(S_1_G_CF_Out[17]) );
  INV_X1 S_1_G_Inst_17__CF_Inst_U1 ( .A(S_1_Rq3[2]), .ZN(
        S_1_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_1_G_InstXOR_0__Compression1_U2 ( .A(
        S_1_G_InstXOR_0__Compression1_n3), .B(S_1_G_CF_Reg[2]), .ZN(
        S_1_G_out1[0]) );
  XNOR2_X1 S_1_G_InstXOR_0__Compression1_U1 ( .A(S_1_G_CF_Reg[0]), .B(
        S_1_G_CF_Reg[1]), .ZN(S_1_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_1_G_InstXOR_0__Compression2_U2 ( .A(
        S_1_G_InstXOR_0__Compression2_n3), .B(S_1_G_CF_Reg[5]), .ZN(
        RF2_SHIFTROWS[9]) );
  XNOR2_X1 S_1_G_InstXOR_0__Compression2_U1 ( .A(S_1_G_CF_Reg[3]), .B(
        S_1_G_CF_Reg[4]), .ZN(S_1_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_1_G_InstXOR_0__Compression3_U2 ( .A(
        S_1_G_InstXOR_0__Compression3_n3), .B(S_1_G_CF_Reg[8]), .ZN(
        RF3_SHIFTROWS[9]) );
  XNOR2_X1 S_1_G_InstXOR_0__Compression3_U1 ( .A(S_1_G_CF_Reg[6]), .B(
        S_1_G_CF_Reg[7]), .ZN(S_1_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_1_G_InstXOR_1__Compression1_U2 ( .A(
        S_1_G_InstXOR_1__Compression1_n3), .B(S_1_G_CF_Reg[11]), .ZN(
        S_1_G_out1[1]) );
  XNOR2_X1 S_1_G_InstXOR_1__Compression1_U1 ( .A(S_1_G_CF_Reg[9]), .B(
        S_1_G_CF_Reg[10]), .ZN(S_1_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_1_G_InstXOR_1__Compression2_U2 ( .A(
        S_1_G_InstXOR_1__Compression2_n3), .B(S_1_G_CF_Reg[14]), .ZN(
        RF2_SHIFTROWS[8]) );
  XNOR2_X1 S_1_G_InstXOR_1__Compression2_U1 ( .A(S_1_G_CF_Reg[12]), .B(
        S_1_G_CF_Reg[13]), .ZN(S_1_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_1_G_InstXOR_1__Compression3_U2 ( .A(
        S_1_G_InstXOR_1__Compression3_n3), .B(S_1_G_CF_Reg[17]), .ZN(
        RF3_SHIFTROWS[8]) );
  XNOR2_X1 S_1_G_InstXOR_1__Compression3_U1 ( .A(S_1_G_CF_Reg[15]), .B(
        S_1_G_CF_Reg[16]), .ZN(S_1_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_1_OutputAffine_U4 ( .A(S_1_G_out1[3]), .ZN(RF1_SHIFTROWS[11]) );
  INV_X1 S_1_OutputAffine_U3 ( .A(S_1_G_out1[2]), .ZN(RF1_SHIFTROWS[10]) );
  INV_X1 S_1_OutputAffine_U2 ( .A(S_1_G_out1[1]), .ZN(RF1_SHIFTROWS[8]) );
  INV_X1 S_1_OutputAffine_U1 ( .A(S_1_G_out1[0]), .ZN(RF1_SHIFTROWS[9]) );
  DFF_X1 S_2_Rq3_reg_0_ ( .D(S_2_q3[0]), .CK(CLK), .Q(S_2_Rq3[0]), .QN() );
  DFF_X1 S_2_Rq3_reg_1_ ( .D(S_2_q3[1]), .CK(CLK), .Q(S_2_Rq3[1]), .QN() );
  DFF_X1 S_2_Rq3_reg_2_ ( .D(S_2_q3[2]), .CK(CLK), .Q(S_2_Rq3[2]), .QN() );
  DFF_X1 S_2_Rq3_reg_3_ ( .D(S_2_q3[3]), .CK(CLK), .Q(S_2_Rq3[3]), .QN() );
  DFF_X1 S_2_Rq2_reg_0_ ( .D(S_2_q2[0]), .CK(CLK), .Q(S_2_Rq2[0]), .QN() );
  DFF_X1 S_2_Rq2_reg_1_ ( .D(S_2_q2[1]), .CK(CLK), .Q(S_2_Rq2[1]), .QN() );
  DFF_X1 S_2_Rq2_reg_2_ ( .D(S_2_q2[2]), .CK(CLK), .Q(S_2_Rq2[2]), .QN() );
  DFF_X1 S_2_Rq2_reg_3_ ( .D(S_2_q2[3]), .CK(CLK), .Q(S_2_Rq2[3]), .QN() );
  DFF_X1 S_2_Rq1_reg_0_ ( .D(S_2_q1[0]), .CK(CLK), .Q(S_2_Rq1[0]), .QN() );
  DFF_X1 S_2_Rq1_reg_1_ ( .D(S_2_q1[1]), .CK(CLK), .Q(S_2_Rq1[1]), .QN() );
  DFF_X1 S_2_Rq1_reg_2_ ( .D(S_2_q1[2]), .CK(CLK), .Q(S_2_Rq1[2]), .QN() );
  DFF_X1 S_2_Rq1_reg_3_ ( .D(S_2_q1[3]), .CK(CLK), .Q(S_2_Rq1[3]), .QN() );
  INV_X1 S_2_InputAffine_U4 ( .A(SUB_IN1[8]), .ZN(S_2_F_in1[0]) );
  INV_X1 S_2_InputAffine_U3 ( .A(SUB_IN1[10]), .ZN(S_2_F_in1[3]) );
  INV_X1 S_2_InputAffine_U2 ( .A(SUB_IN1[11]), .ZN(S_2_F_in1[1]) );
  INV_X1 S_2_InputAffine_U1 ( .A(SUB_IN1[9]), .ZN(S_2_F_in1[2]) );
  XNOR2_X1 S_2_F_U18 ( .A(S_2_F_n12), .B(FRESH[19]), .ZN(S_2_q3[3]) );
  XNOR2_X1 S_2_F_U17 ( .A(FRESH[18]), .B(S_2_F_q3[3]), .ZN(S_2_F_n12) );
  XNOR2_X1 S_2_F_U16 ( .A(S_2_F_n11), .B(FRESH[17]), .ZN(S_2_q3[2]) );
  XNOR2_X1 S_2_F_U15 ( .A(FRESH[16]), .B(S_2_F_q3[2]), .ZN(S_2_F_n11) );
  XOR2_X1 S_2_F_U14 ( .A(FRESH[19]), .B(S_2_F_q2[3]), .Z(S_2_q2[3]) );
  XOR2_X1 S_2_F_U13 ( .A(FRESH[17]), .B(S_2_F_q2[2]), .Z(S_2_q2[2]) );
  XOR2_X1 S_2_F_U12 ( .A(FRESH[18]), .B(S_2_F_q1[3]), .Z(S_2_q1[3]) );
  XOR2_X1 S_2_F_U11 ( .A(FRESH[16]), .B(S_2_F_q1[2]), .Z(S_2_q1[2]) );
  XNOR2_X1 S_2_F_U10 ( .A(S_2_F_n10), .B(FRESH[21]), .ZN(S_2_F_N5) );
  XNOR2_X1 S_2_F_U9 ( .A(S_2_F_in3[3]), .B(FRESH[20]), .ZN(S_2_F_n10) );
  XOR2_X1 S_2_F_U8 ( .A(FRESH[21]), .B(S_2_F_in2[3]), .Z(S_2_F_N4) );
  XOR2_X1 S_2_F_U7 ( .A(FRESH[20]), .B(S_2_F_in1[3]), .Z(S_2_F_N3) );
  XNOR2_X1 S_2_F_U6 ( .A(S_2_F_n9), .B(FRESH[23]), .ZN(S_2_F_N2) );
  XNOR2_X1 S_2_F_U5 ( .A(S_2_F_in3[2]), .B(FRESH[22]), .ZN(S_2_F_n9) );
  XOR2_X1 S_2_F_U4 ( .A(FRESH[23]), .B(S_2_F_in2[2]), .Z(S_2_F_N1) );
  XOR2_X1 S_2_F_U3 ( .A(FRESH[22]), .B(S_2_F_in1[2]), .Z(S_2_F_N0) );
  DFF_X1 S_2_F_CF_Reg_reg_0_ ( .D(S_2_F_CF_Out[0]), .CK(CLK), .Q(
        S_2_F_CF_Reg[0]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_1_ ( .D(S_2_F_CF_Out[1]), .CK(CLK), .Q(
        S_2_F_CF_Reg[1]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_2_ ( .D(S_2_F_CF_Out[2]), .CK(CLK), .Q(
        S_2_F_CF_Reg[2]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_3_ ( .D(S_2_F_CF_Out[3]), .CK(CLK), .Q(
        S_2_F_CF_Reg[3]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_4_ ( .D(S_2_F_CF_Out[4]), .CK(CLK), .Q(
        S_2_F_CF_Reg[4]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_5_ ( .D(S_2_F_CF_Out[5]), .CK(CLK), .Q(
        S_2_F_CF_Reg[5]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_6_ ( .D(S_2_F_CF_Out[6]), .CK(CLK), .Q(
        S_2_F_CF_Reg[6]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_7_ ( .D(S_2_F_CF_Out[7]), .CK(CLK), .Q(
        S_2_F_CF_Reg[7]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_8_ ( .D(S_2_F_CF_Out[8]), .CK(CLK), .Q(
        S_2_F_CF_Reg[8]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_9_ ( .D(S_2_F_CF_Out[9]), .CK(CLK), .Q(
        S_2_F_CF_Reg[9]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_10_ ( .D(S_2_F_CF_Out[10]), .CK(CLK), .Q(
        S_2_F_CF_Reg[10]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_11_ ( .D(S_2_F_CF_Out[11]), .CK(CLK), .Q(
        S_2_F_CF_Reg[11]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_12_ ( .D(S_2_F_CF_Out[12]), .CK(CLK), .Q(
        S_2_F_CF_Reg[12]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_13_ ( .D(S_2_F_CF_Out[13]), .CK(CLK), .Q(
        S_2_F_CF_Reg[13]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_14_ ( .D(S_2_F_CF_Out[14]), .CK(CLK), .Q(
        S_2_F_CF_Reg[14]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_15_ ( .D(S_2_F_CF_Out[15]), .CK(CLK), .Q(
        S_2_F_CF_Reg[15]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_16_ ( .D(S_2_F_CF_Out[16]), .CK(CLK), .Q(
        S_2_F_CF_Reg[16]), .QN() );
  DFF_X1 S_2_F_CF_Reg_reg_17_ ( .D(S_2_F_CF_Out[17]), .CK(CLK), .Q(
        S_2_F_CF_Reg[17]), .QN() );
  DFF_X1 S_2_F_out2_reg_0_ ( .D(S_2_F_N4), .CK(CLK), .Q(S_2_q2[0]), .QN() );
  DFF_X1 S_2_F_out2_reg_1_ ( .D(S_2_F_N1), .CK(CLK), .Q(S_2_q2[1]), .QN() );
  DFF_X1 S_2_F_out3_reg_0_ ( .D(S_2_F_N5), .CK(CLK), .Q(S_2_q3[0]), .QN() );
  DFF_X1 S_2_F_out3_reg_1_ ( .D(S_2_F_N2), .CK(CLK), .Q(S_2_q3[1]), .QN() );
  DFF_X1 S_2_F_out1_reg_0_ ( .D(S_2_F_N3), .CK(CLK), .Q(S_2_q1[0]), .QN() );
  DFF_X1 S_2_F_out1_reg_1_ ( .D(S_2_F_N0), .CK(CLK), .Q(S_2_q1[1]), .QN() );
  NOR2_X1 S_2_F_Inst_0__CF_Inst_U2 ( .A1(S_2_F_in1[2]), .A2(
        S_2_F_Inst_0__CF_Inst_n3), .ZN(S_2_F_CF_Out[0]) );
  INV_X1 S_2_F_Inst_0__CF_Inst_U1 ( .A(S_2_F_in1[3]), .ZN(
        S_2_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_2_F_Inst_1__CF_Inst_U2 ( .A(S_2_F_Inst_1__CF_Inst_n3), .B(
        S_2_F_in1[1]), .ZN(S_2_F_CF_Out[1]) );
  NAND2_X1 S_2_F_Inst_1__CF_Inst_U1 ( .A1(S_2_F_in2[2]), .A2(S_2_F_in1[3]), 
        .ZN(S_2_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_2_F_Inst_2__CF_Inst_U1 ( .A1(S_2_F_in1[3]), .A2(S_2_F_in3[2]), .ZN(
        S_2_F_CF_Out[2]) );
  NOR2_X1 S_2_F_Inst_3__CF_Inst_U2 ( .A1(S_2_F_in2[3]), .A2(
        S_2_F_Inst_3__CF_Inst_n3), .ZN(S_2_F_CF_Out[3]) );
  INV_X1 S_2_F_Inst_3__CF_Inst_U1 ( .A(S_2_F_in1[2]), .ZN(
        S_2_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_2_F_Inst_4__CF_Inst_U2 ( .A(S_2_F_Inst_4__CF_Inst_n3), .B(
        S_2_F_in2[1]), .ZN(S_2_F_CF_Out[4]) );
  NAND2_X1 S_2_F_Inst_4__CF_Inst_U1 ( .A1(S_2_F_in2[2]), .A2(S_2_F_in2[3]), 
        .ZN(S_2_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_2_F_Inst_5__CF_Inst_U1 ( .A1(S_2_F_in3[2]), .A2(S_2_F_in2[3]), 
        .ZN(S_2_F_CF_Out[5]) );
  XNOR2_X1 S_2_F_Inst_6__CF_Inst_U2 ( .A(S_2_F_Inst_6__CF_Inst_n7), .B(
        S_2_F_in3[1]), .ZN(S_2_F_CF_Out[6]) );
  NOR2_X1 S_2_F_Inst_6__CF_Inst_U1 ( .A1(S_2_F_in1[2]), .A2(S_2_F_in3[3]), 
        .ZN(S_2_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_2_F_Inst_7__CF_Inst_U1 ( .A1(S_2_F_in2[2]), .A2(S_2_F_in3[3]), 
        .ZN(S_2_F_CF_Out[7]) );
  OR2_X1 S_2_F_Inst_8__CF_Inst_U1 ( .A1(S_2_F_in3[3]), .A2(S_2_F_in3[2]), .ZN(
        S_2_F_CF_Out[8]) );
  NOR2_X1 S_2_F_Inst_9__CF_Inst_U2 ( .A1(S_2_F_in1[3]), .A2(
        S_2_F_Inst_9__CF_Inst_n3), .ZN(S_2_F_CF_Out[9]) );
  INV_X1 S_2_F_Inst_9__CF_Inst_U1 ( .A(S_2_F_in1[1]), .ZN(
        S_2_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_2_F_Inst_10__CF_Inst_U1 ( .A1(S_2_F_in2[1]), .A2(S_2_F_in1[3]), 
        .ZN(S_2_F_CF_Out[10]) );
  XNOR2_X1 S_2_F_Inst_11__CF_Inst_U2 ( .A(S_2_F_Inst_11__CF_Inst_n3), .B(
        S_2_F_in1[0]), .ZN(S_2_F_CF_Out[11]) );
  NAND2_X1 S_2_F_Inst_11__CF_Inst_U1 ( .A1(S_2_F_in3[1]), .A2(S_2_F_in1[3]), 
        .ZN(S_2_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_2_F_Inst_12__CF_Inst_U2 ( .A(S_2_F_Inst_12__CF_Inst_n3), .B(
        S_2_F_in2[0]), .ZN(S_2_F_CF_Out[12]) );
  NAND2_X1 S_2_F_Inst_12__CF_Inst_U1 ( .A1(S_2_F_in1[1]), .A2(S_2_F_in2[3]), 
        .ZN(S_2_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_2_F_Inst_13__CF_Inst_U2 ( .A1(S_2_F_in2[3]), .A2(
        S_2_F_Inst_13__CF_Inst_n3), .ZN(S_2_F_CF_Out[13]) );
  INV_X1 S_2_F_Inst_13__CF_Inst_U1 ( .A(S_2_F_in2[1]), .ZN(
        S_2_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_2_F_Inst_14__CF_Inst_U1 ( .A1(S_2_F_in3[1]), .A2(S_2_F_in2[3]), 
        .ZN(S_2_F_CF_Out[14]) );
  XNOR2_X1 S_2_F_Inst_15__CF_Inst_U2 ( .A(S_2_F_Inst_15__CF_Inst_n7), .B(
        S_2_F_in3[0]), .ZN(S_2_F_CF_Out[15]) );
  NOR2_X1 S_2_F_Inst_15__CF_Inst_U1 ( .A1(S_2_F_in1[1]), .A2(S_2_F_in3[3]), 
        .ZN(S_2_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_2_F_Inst_16__CF_Inst_U2 ( .A1(S_2_F_in3[3]), .A2(
        S_2_F_Inst_16__CF_Inst_n3), .ZN(S_2_F_CF_Out[16]) );
  INV_X1 S_2_F_Inst_16__CF_Inst_U1 ( .A(S_2_F_in2[1]), .ZN(
        S_2_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_2_F_Inst_17__CF_Inst_U2 ( .A1(S_2_F_in3[1]), .A2(
        S_2_F_Inst_17__CF_Inst_n3), .ZN(S_2_F_CF_Out[17]) );
  INV_X1 S_2_F_Inst_17__CF_Inst_U1 ( .A(S_2_F_in3[3]), .ZN(
        S_2_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_2_F_InstXOR_0__Compression1_U2 ( .A(
        S_2_F_InstXOR_0__Compression1_n3), .B(S_2_F_CF_Reg[2]), .ZN(
        S_2_F_q1[2]) );
  XNOR2_X1 S_2_F_InstXOR_0__Compression1_U1 ( .A(S_2_F_CF_Reg[0]), .B(
        S_2_F_CF_Reg[1]), .ZN(S_2_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_2_F_InstXOR_0__Compression2_U2 ( .A(
        S_2_F_InstXOR_0__Compression2_n3), .B(S_2_F_CF_Reg[5]), .ZN(
        S_2_F_q2[2]) );
  XNOR2_X1 S_2_F_InstXOR_0__Compression2_U1 ( .A(S_2_F_CF_Reg[3]), .B(
        S_2_F_CF_Reg[4]), .ZN(S_2_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_2_F_InstXOR_0__Compression3_U2 ( .A(
        S_2_F_InstXOR_0__Compression3_n3), .B(S_2_F_CF_Reg[8]), .ZN(
        S_2_F_q3[2]) );
  XNOR2_X1 S_2_F_InstXOR_0__Compression3_U1 ( .A(S_2_F_CF_Reg[6]), .B(
        S_2_F_CF_Reg[7]), .ZN(S_2_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_2_F_InstXOR_1__Compression1_U2 ( .A(
        S_2_F_InstXOR_1__Compression1_n3), .B(S_2_F_CF_Reg[11]), .ZN(
        S_2_F_q1[3]) );
  XNOR2_X1 S_2_F_InstXOR_1__Compression1_U1 ( .A(S_2_F_CF_Reg[9]), .B(
        S_2_F_CF_Reg[10]), .ZN(S_2_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_2_F_InstXOR_1__Compression2_U2 ( .A(
        S_2_F_InstXOR_1__Compression2_n3), .B(S_2_F_CF_Reg[14]), .ZN(
        S_2_F_q2[3]) );
  XNOR2_X1 S_2_F_InstXOR_1__Compression2_U1 ( .A(S_2_F_CF_Reg[12]), .B(
        S_2_F_CF_Reg[13]), .ZN(S_2_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_2_F_InstXOR_1__Compression3_U2 ( .A(
        S_2_F_InstXOR_1__Compression3_n3), .B(S_2_F_CF_Reg[17]), .ZN(
        S_2_F_q3[3]) );
  XNOR2_X1 S_2_F_InstXOR_1__Compression3_U1 ( .A(S_2_F_CF_Reg[15]), .B(
        S_2_F_CF_Reg[16]), .ZN(S_2_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_2_G_CF_Reg_reg_0_ ( .D(S_2_G_CF_Out[0]), .CK(CLK), .Q(
        S_2_G_CF_Reg[0]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_1_ ( .D(S_2_G_CF_Out[1]), .CK(CLK), .Q(
        S_2_G_CF_Reg[1]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_2_ ( .D(S_2_G_CF_Out[2]), .CK(CLK), .Q(
        S_2_G_CF_Reg[2]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_3_ ( .D(S_2_G_CF_Out[3]), .CK(CLK), .Q(
        S_2_G_CF_Reg[3]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_4_ ( .D(S_2_G_CF_Out[4]), .CK(CLK), .Q(
        S_2_G_CF_Reg[4]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_5_ ( .D(S_2_G_CF_Out[5]), .CK(CLK), .Q(
        S_2_G_CF_Reg[5]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_6_ ( .D(S_2_G_CF_Out[6]), .CK(CLK), .Q(
        S_2_G_CF_Reg[6]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_7_ ( .D(S_2_G_CF_Out[7]), .CK(CLK), .Q(
        S_2_G_CF_Reg[7]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_8_ ( .D(S_2_G_CF_Out[8]), .CK(CLK), .Q(
        S_2_G_CF_Reg[8]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_9_ ( .D(S_2_G_CF_Out[9]), .CK(CLK), .Q(
        S_2_G_CF_Reg[9]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_10_ ( .D(S_2_G_CF_Out[10]), .CK(CLK), .Q(
        S_2_G_CF_Reg[10]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_11_ ( .D(S_2_G_CF_Out[11]), .CK(CLK), .Q(
        S_2_G_CF_Reg[11]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_12_ ( .D(S_2_G_CF_Out[12]), .CK(CLK), .Q(
        S_2_G_CF_Reg[12]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_13_ ( .D(S_2_G_CF_Out[13]), .CK(CLK), .Q(
        S_2_G_CF_Reg[13]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_14_ ( .D(S_2_G_CF_Out[14]), .CK(CLK), .Q(
        S_2_G_CF_Reg[14]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_15_ ( .D(S_2_G_CF_Out[15]), .CK(CLK), .Q(
        S_2_G_CF_Reg[15]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_16_ ( .D(S_2_G_CF_Out[16]), .CK(CLK), .Q(
        S_2_G_CF_Reg[16]), .QN() );
  DFF_X1 S_2_G_CF_Reg_reg_17_ ( .D(S_2_G_CF_Out[17]), .CK(CLK), .Q(
        S_2_G_CF_Reg[17]), .QN() );
  DFF_X1 S_2_G_out1_reg_2_ ( .D(S_2_Rq1[2]), .CK(CLK), .Q(S_2_G_out1[2]), 
        .QN() );
  DFF_X1 S_2_G_out1_reg_3_ ( .D(S_2_Rq1[3]), .CK(CLK), .Q(S_2_G_out1[3]), 
        .QN() );
  DFF_X1 S_2_G_out2_reg_2_ ( .D(S_2_Rq2[2]), .CK(CLK), .Q(RF2_SHIFTROWS[14]), 
        .QN() );
  DFF_X1 S_2_G_out2_reg_3_ ( .D(S_2_Rq2[3]), .CK(CLK), .Q(RF2_SHIFTROWS[15]), 
        .QN() );
  DFF_X1 S_2_G_out3_reg_2_ ( .D(S_2_Rq3[2]), .CK(CLK), .Q(RF3_SHIFTROWS[14]), 
        .QN() );
  DFF_X1 S_2_G_out3_reg_3_ ( .D(S_2_Rq3[3]), .CK(CLK), .Q(RF3_SHIFTROWS[15]), 
        .QN() );
  AND2_X1 S_2_G_Inst_0__CF_Inst_U1 ( .A1(S_2_Rq1[1]), .A2(S_2_Rq1[3]), .ZN(
        S_2_G_CF_Out[0]) );
  NOR2_X1 S_2_G_Inst_1__CF_Inst_U2 ( .A1(S_2_Rq1[3]), .A2(
        S_2_G_Inst_1__CF_Inst_n3), .ZN(S_2_G_CF_Out[1]) );
  INV_X1 S_2_G_Inst_1__CF_Inst_U1 ( .A(S_2_Rq2[1]), .ZN(
        S_2_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_2_G_Inst_2__CF_Inst_U2 ( .A(S_2_G_Inst_2__CF_Inst_n3), .B(
        S_2_Rq2[0]), .ZN(S_2_G_CF_Out[2]) );
  NAND2_X1 S_2_G_Inst_2__CF_Inst_U1 ( .A1(S_2_Rq1[1]), .A2(S_2_Rq2[3]), .ZN(
        S_2_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_2_G_Inst_3__CF_Inst_U3 ( .A(S_2_Rq1[0]), .B(
        S_2_G_Inst_3__CF_Inst_n6), .ZN(S_2_G_CF_Out[3]) );
  NAND2_X1 S_2_G_Inst_3__CF_Inst_U2 ( .A1(S_2_Rq3[1]), .A2(
        S_2_G_Inst_3__CF_Inst_n5), .ZN(S_2_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_2_G_Inst_3__CF_Inst_U1 ( .A(S_2_Rq1[3]), .ZN(
        S_2_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_2_G_Inst_4__CF_Inst_U1 ( .A1(S_2_Rq2[1]), .A2(S_2_Rq2[3]), .ZN(
        S_2_G_CF_Out[4]) );
  OR2_X1 S_2_G_Inst_5__CF_Inst_U1 ( .A1(S_2_Rq3[3]), .A2(S_2_Rq2[1]), .ZN(
        S_2_G_CF_Out[5]) );
  AND2_X1 S_2_G_Inst_6__CF_Inst_U1 ( .A1(S_2_Rq3[1]), .A2(S_2_Rq2[3]), .ZN(
        S_2_G_CF_Out[6]) );
  XNOR2_X1 S_2_G_Inst_7__CF_Inst_U2 ( .A(S_2_G_Inst_7__CF_Inst_n3), .B(
        S_2_Rq3[0]), .ZN(S_2_G_CF_Out[7]) );
  NAND2_X1 S_2_G_Inst_7__CF_Inst_U1 ( .A1(S_2_Rq1[1]), .A2(S_2_Rq3[3]), .ZN(
        S_2_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_2_G_Inst_8__CF_Inst_U1 ( .A1(S_2_Rq3[3]), .A2(S_2_Rq3[1]), .ZN(
        S_2_G_CF_Out[8]) );
  NOR2_X1 S_2_G_Inst_9__CF_Inst_U2 ( .A1(S_2_Rq1[3]), .A2(
        S_2_G_Inst_9__CF_Inst_n3), .ZN(S_2_G_CF_Out[9]) );
  INV_X1 S_2_G_Inst_9__CF_Inst_U1 ( .A(S_2_Rq1[2]), .ZN(
        S_2_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_2_G_Inst_10__CF_Inst_U2 ( .A1(S_2_Rq2[2]), .A2(
        S_2_G_Inst_10__CF_Inst_n3), .ZN(S_2_G_CF_Out[10]) );
  INV_X1 S_2_G_Inst_10__CF_Inst_U1 ( .A(S_2_Rq1[3]), .ZN(
        S_2_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_2_G_Inst_11__CF_Inst_U3 ( .A(S_2_Rq1[1]), .B(
        S_2_G_Inst_11__CF_Inst_n6), .ZN(S_2_G_CF_Out[11]) );
  NAND2_X1 S_2_G_Inst_11__CF_Inst_U2 ( .A1(S_2_Rq1[3]), .A2(
        S_2_G_Inst_11__CF_Inst_n5), .ZN(S_2_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_2_G_Inst_11__CF_Inst_U1 ( .A(S_2_Rq3[2]), .ZN(
        S_2_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_2_G_Inst_12__CF_Inst_U2 ( .A1(S_2_Rq2[3]), .A2(
        S_2_G_Inst_12__CF_Inst_n3), .ZN(S_2_G_CF_Out[12]) );
  INV_X1 S_2_G_Inst_12__CF_Inst_U1 ( .A(S_2_Rq1[2]), .ZN(
        S_2_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_2_G_Inst_13__CF_Inst_U1 ( .A1(S_2_Rq2[2]), .A2(S_2_Rq2[3]), .ZN(
        S_2_G_CF_Out[13]) );
  XNOR2_X1 S_2_G_Inst_14__CF_Inst_U3 ( .A(S_2_Rq2[1]), .B(
        S_2_G_Inst_14__CF_Inst_n6), .ZN(S_2_G_CF_Out[14]) );
  NAND2_X1 S_2_G_Inst_14__CF_Inst_U2 ( .A1(S_2_Rq3[2]), .A2(
        S_2_G_Inst_14__CF_Inst_n5), .ZN(S_2_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_2_G_Inst_14__CF_Inst_U1 ( .A(S_2_Rq2[3]), .ZN(
        S_2_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_2_G_Inst_15__CF_Inst_U2 ( .A(S_2_G_Inst_15__CF_Inst_n3), .B(
        S_2_Rq3[1]), .ZN(S_2_G_CF_Out[15]) );
  NAND2_X1 S_2_G_Inst_15__CF_Inst_U1 ( .A1(S_2_Rq1[2]), .A2(S_2_Rq3[3]), .ZN(
        S_2_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_2_G_Inst_16__CF_Inst_U1 ( .A1(S_2_Rq2[2]), .A2(S_2_Rq3[3]), .ZN(
        S_2_G_CF_Out[16]) );
  NOR2_X1 S_2_G_Inst_17__CF_Inst_U2 ( .A1(S_2_Rq3[3]), .A2(
        S_2_G_Inst_17__CF_Inst_n3), .ZN(S_2_G_CF_Out[17]) );
  INV_X1 S_2_G_Inst_17__CF_Inst_U1 ( .A(S_2_Rq3[2]), .ZN(
        S_2_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_2_G_InstXOR_0__Compression1_U2 ( .A(
        S_2_G_InstXOR_0__Compression1_n3), .B(S_2_G_CF_Reg[2]), .ZN(
        S_2_G_out1[0]) );
  XNOR2_X1 S_2_G_InstXOR_0__Compression1_U1 ( .A(S_2_G_CF_Reg[0]), .B(
        S_2_G_CF_Reg[1]), .ZN(S_2_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_2_G_InstXOR_0__Compression2_U2 ( .A(
        S_2_G_InstXOR_0__Compression2_n3), .B(S_2_G_CF_Reg[5]), .ZN(
        RF2_SHIFTROWS[13]) );
  XNOR2_X1 S_2_G_InstXOR_0__Compression2_U1 ( .A(S_2_G_CF_Reg[3]), .B(
        S_2_G_CF_Reg[4]), .ZN(S_2_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_2_G_InstXOR_0__Compression3_U2 ( .A(
        S_2_G_InstXOR_0__Compression3_n3), .B(S_2_G_CF_Reg[8]), .ZN(
        RF3_SHIFTROWS[13]) );
  XNOR2_X1 S_2_G_InstXOR_0__Compression3_U1 ( .A(S_2_G_CF_Reg[6]), .B(
        S_2_G_CF_Reg[7]), .ZN(S_2_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_2_G_InstXOR_1__Compression1_U2 ( .A(
        S_2_G_InstXOR_1__Compression1_n3), .B(S_2_G_CF_Reg[11]), .ZN(
        S_2_G_out1[1]) );
  XNOR2_X1 S_2_G_InstXOR_1__Compression1_U1 ( .A(S_2_G_CF_Reg[9]), .B(
        S_2_G_CF_Reg[10]), .ZN(S_2_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_2_G_InstXOR_1__Compression2_U2 ( .A(
        S_2_G_InstXOR_1__Compression2_n3), .B(S_2_G_CF_Reg[14]), .ZN(
        RF2_SHIFTROWS[12]) );
  XNOR2_X1 S_2_G_InstXOR_1__Compression2_U1 ( .A(S_2_G_CF_Reg[12]), .B(
        S_2_G_CF_Reg[13]), .ZN(S_2_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_2_G_InstXOR_1__Compression3_U2 ( .A(
        S_2_G_InstXOR_1__Compression3_n3), .B(S_2_G_CF_Reg[17]), .ZN(
        RF3_SHIFTROWS[12]) );
  XNOR2_X1 S_2_G_InstXOR_1__Compression3_U1 ( .A(S_2_G_CF_Reg[15]), .B(
        S_2_G_CF_Reg[16]), .ZN(S_2_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_2_OutputAffine_U4 ( .A(S_2_G_out1[3]), .ZN(RF1_SHIFTROWS[15]) );
  INV_X1 S_2_OutputAffine_U3 ( .A(S_2_G_out1[2]), .ZN(RF1_SHIFTROWS[14]) );
  INV_X1 S_2_OutputAffine_U2 ( .A(S_2_G_out1[1]), .ZN(RF1_SHIFTROWS[12]) );
  INV_X1 S_2_OutputAffine_U1 ( .A(S_2_G_out1[0]), .ZN(RF1_SHIFTROWS[13]) );
  DFF_X1 S_3_Rq3_reg_0_ ( .D(S_3_q3[0]), .CK(CLK), .Q(S_3_Rq3[0]), .QN() );
  DFF_X1 S_3_Rq3_reg_1_ ( .D(S_3_q3[1]), .CK(CLK), .Q(S_3_Rq3[1]), .QN() );
  DFF_X1 S_3_Rq3_reg_2_ ( .D(S_3_q3[2]), .CK(CLK), .Q(S_3_Rq3[2]), .QN() );
  DFF_X1 S_3_Rq3_reg_3_ ( .D(S_3_q3[3]), .CK(CLK), .Q(S_3_Rq3[3]), .QN() );
  DFF_X1 S_3_Rq2_reg_0_ ( .D(S_3_q2[0]), .CK(CLK), .Q(S_3_Rq2[0]), .QN() );
  DFF_X1 S_3_Rq2_reg_1_ ( .D(S_3_q2[1]), .CK(CLK), .Q(S_3_Rq2[1]), .QN() );
  DFF_X1 S_3_Rq2_reg_2_ ( .D(S_3_q2[2]), .CK(CLK), .Q(S_3_Rq2[2]), .QN() );
  DFF_X1 S_3_Rq2_reg_3_ ( .D(S_3_q2[3]), .CK(CLK), .Q(S_3_Rq2[3]), .QN() );
  DFF_X1 S_3_Rq1_reg_0_ ( .D(S_3_q1[0]), .CK(CLK), .Q(S_3_Rq1[0]), .QN() );
  DFF_X1 S_3_Rq1_reg_1_ ( .D(S_3_q1[1]), .CK(CLK), .Q(S_3_Rq1[1]), .QN() );
  DFF_X1 S_3_Rq1_reg_2_ ( .D(S_3_q1[2]), .CK(CLK), .Q(S_3_Rq1[2]), .QN() );
  DFF_X1 S_3_Rq1_reg_3_ ( .D(S_3_q1[3]), .CK(CLK), .Q(S_3_Rq1[3]), .QN() );
  INV_X1 S_3_InputAffine_U4 ( .A(SUB_IN1[12]), .ZN(S_3_F_in1[0]) );
  INV_X1 S_3_InputAffine_U3 ( .A(SUB_IN1[14]), .ZN(S_3_F_in1[3]) );
  INV_X1 S_3_InputAffine_U2 ( .A(SUB_IN1[15]), .ZN(S_3_F_in1[1]) );
  INV_X1 S_3_InputAffine_U1 ( .A(SUB_IN1[13]), .ZN(S_3_F_in1[2]) );
  XNOR2_X1 S_3_F_U18 ( .A(S_3_F_n12), .B(FRESH[27]), .ZN(S_3_q3[3]) );
  XNOR2_X1 S_3_F_U17 ( .A(FRESH[26]), .B(S_3_F_q3[3]), .ZN(S_3_F_n12) );
  XNOR2_X1 S_3_F_U16 ( .A(S_3_F_n11), .B(FRESH[25]), .ZN(S_3_q3[2]) );
  XNOR2_X1 S_3_F_U15 ( .A(FRESH[24]), .B(S_3_F_q3[2]), .ZN(S_3_F_n11) );
  XOR2_X1 S_3_F_U14 ( .A(FRESH[27]), .B(S_3_F_q2[3]), .Z(S_3_q2[3]) );
  XOR2_X1 S_3_F_U13 ( .A(FRESH[25]), .B(S_3_F_q2[2]), .Z(S_3_q2[2]) );
  XOR2_X1 S_3_F_U12 ( .A(FRESH[26]), .B(S_3_F_q1[3]), .Z(S_3_q1[3]) );
  XOR2_X1 S_3_F_U11 ( .A(FRESH[24]), .B(S_3_F_q1[2]), .Z(S_3_q1[2]) );
  XNOR2_X1 S_3_F_U10 ( .A(S_3_F_n10), .B(FRESH[29]), .ZN(S_3_F_N5) );
  XNOR2_X1 S_3_F_U9 ( .A(S_3_F_in3[3]), .B(FRESH[28]), .ZN(S_3_F_n10) );
  XOR2_X1 S_3_F_U8 ( .A(FRESH[29]), .B(S_3_F_in2[3]), .Z(S_3_F_N4) );
  XOR2_X1 S_3_F_U7 ( .A(FRESH[28]), .B(S_3_F_in1[3]), .Z(S_3_F_N3) );
  XNOR2_X1 S_3_F_U6 ( .A(S_3_F_n9), .B(FRESH[31]), .ZN(S_3_F_N2) );
  XNOR2_X1 S_3_F_U5 ( .A(S_3_F_in3[2]), .B(FRESH[30]), .ZN(S_3_F_n9) );
  XOR2_X1 S_3_F_U4 ( .A(FRESH[31]), .B(S_3_F_in2[2]), .Z(S_3_F_N1) );
  XOR2_X1 S_3_F_U3 ( .A(FRESH[30]), .B(S_3_F_in1[2]), .Z(S_3_F_N0) );
  DFF_X1 S_3_F_CF_Reg_reg_0_ ( .D(S_3_F_CF_Out[0]), .CK(CLK), .Q(
        S_3_F_CF_Reg[0]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_1_ ( .D(S_3_F_CF_Out[1]), .CK(CLK), .Q(
        S_3_F_CF_Reg[1]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_2_ ( .D(S_3_F_CF_Out[2]), .CK(CLK), .Q(
        S_3_F_CF_Reg[2]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_3_ ( .D(S_3_F_CF_Out[3]), .CK(CLK), .Q(
        S_3_F_CF_Reg[3]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_4_ ( .D(S_3_F_CF_Out[4]), .CK(CLK), .Q(
        S_3_F_CF_Reg[4]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_5_ ( .D(S_3_F_CF_Out[5]), .CK(CLK), .Q(
        S_3_F_CF_Reg[5]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_6_ ( .D(S_3_F_CF_Out[6]), .CK(CLK), .Q(
        S_3_F_CF_Reg[6]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_7_ ( .D(S_3_F_CF_Out[7]), .CK(CLK), .Q(
        S_3_F_CF_Reg[7]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_8_ ( .D(S_3_F_CF_Out[8]), .CK(CLK), .Q(
        S_3_F_CF_Reg[8]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_9_ ( .D(S_3_F_CF_Out[9]), .CK(CLK), .Q(
        S_3_F_CF_Reg[9]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_10_ ( .D(S_3_F_CF_Out[10]), .CK(CLK), .Q(
        S_3_F_CF_Reg[10]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_11_ ( .D(S_3_F_CF_Out[11]), .CK(CLK), .Q(
        S_3_F_CF_Reg[11]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_12_ ( .D(S_3_F_CF_Out[12]), .CK(CLK), .Q(
        S_3_F_CF_Reg[12]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_13_ ( .D(S_3_F_CF_Out[13]), .CK(CLK), .Q(
        S_3_F_CF_Reg[13]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_14_ ( .D(S_3_F_CF_Out[14]), .CK(CLK), .Q(
        S_3_F_CF_Reg[14]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_15_ ( .D(S_3_F_CF_Out[15]), .CK(CLK), .Q(
        S_3_F_CF_Reg[15]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_16_ ( .D(S_3_F_CF_Out[16]), .CK(CLK), .Q(
        S_3_F_CF_Reg[16]), .QN() );
  DFF_X1 S_3_F_CF_Reg_reg_17_ ( .D(S_3_F_CF_Out[17]), .CK(CLK), .Q(
        S_3_F_CF_Reg[17]), .QN() );
  DFF_X1 S_3_F_out2_reg_0_ ( .D(S_3_F_N4), .CK(CLK), .Q(S_3_q2[0]), .QN() );
  DFF_X1 S_3_F_out2_reg_1_ ( .D(S_3_F_N1), .CK(CLK), .Q(S_3_q2[1]), .QN() );
  DFF_X1 S_3_F_out3_reg_0_ ( .D(S_3_F_N5), .CK(CLK), .Q(S_3_q3[0]), .QN() );
  DFF_X1 S_3_F_out3_reg_1_ ( .D(S_3_F_N2), .CK(CLK), .Q(S_3_q3[1]), .QN() );
  DFF_X1 S_3_F_out1_reg_0_ ( .D(S_3_F_N3), .CK(CLK), .Q(S_3_q1[0]), .QN() );
  DFF_X1 S_3_F_out1_reg_1_ ( .D(S_3_F_N0), .CK(CLK), .Q(S_3_q1[1]), .QN() );
  NOR2_X1 S_3_F_Inst_0__CF_Inst_U2 ( .A1(S_3_F_in1[2]), .A2(
        S_3_F_Inst_0__CF_Inst_n3), .ZN(S_3_F_CF_Out[0]) );
  INV_X1 S_3_F_Inst_0__CF_Inst_U1 ( .A(S_3_F_in1[3]), .ZN(
        S_3_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_3_F_Inst_1__CF_Inst_U2 ( .A(S_3_F_Inst_1__CF_Inst_n3), .B(
        S_3_F_in1[1]), .ZN(S_3_F_CF_Out[1]) );
  NAND2_X1 S_3_F_Inst_1__CF_Inst_U1 ( .A1(S_3_F_in2[2]), .A2(S_3_F_in1[3]), 
        .ZN(S_3_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_3_F_Inst_2__CF_Inst_U1 ( .A1(S_3_F_in1[3]), .A2(S_3_F_in3[2]), .ZN(
        S_3_F_CF_Out[2]) );
  NOR2_X1 S_3_F_Inst_3__CF_Inst_U2 ( .A1(S_3_F_in2[3]), .A2(
        S_3_F_Inst_3__CF_Inst_n3), .ZN(S_3_F_CF_Out[3]) );
  INV_X1 S_3_F_Inst_3__CF_Inst_U1 ( .A(S_3_F_in1[2]), .ZN(
        S_3_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_3_F_Inst_4__CF_Inst_U2 ( .A(S_3_F_Inst_4__CF_Inst_n3), .B(
        S_3_F_in2[1]), .ZN(S_3_F_CF_Out[4]) );
  NAND2_X1 S_3_F_Inst_4__CF_Inst_U1 ( .A1(S_3_F_in2[2]), .A2(S_3_F_in2[3]), 
        .ZN(S_3_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_3_F_Inst_5__CF_Inst_U1 ( .A1(S_3_F_in3[2]), .A2(S_3_F_in2[3]), 
        .ZN(S_3_F_CF_Out[5]) );
  XNOR2_X1 S_3_F_Inst_6__CF_Inst_U2 ( .A(S_3_F_Inst_6__CF_Inst_n7), .B(
        S_3_F_in3[1]), .ZN(S_3_F_CF_Out[6]) );
  NOR2_X1 S_3_F_Inst_6__CF_Inst_U1 ( .A1(S_3_F_in1[2]), .A2(S_3_F_in3[3]), 
        .ZN(S_3_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_3_F_Inst_7__CF_Inst_U1 ( .A1(S_3_F_in2[2]), .A2(S_3_F_in3[3]), 
        .ZN(S_3_F_CF_Out[7]) );
  OR2_X1 S_3_F_Inst_8__CF_Inst_U1 ( .A1(S_3_F_in3[3]), .A2(S_3_F_in3[2]), .ZN(
        S_3_F_CF_Out[8]) );
  NOR2_X1 S_3_F_Inst_9__CF_Inst_U2 ( .A1(S_3_F_in1[3]), .A2(
        S_3_F_Inst_9__CF_Inst_n3), .ZN(S_3_F_CF_Out[9]) );
  INV_X1 S_3_F_Inst_9__CF_Inst_U1 ( .A(S_3_F_in1[1]), .ZN(
        S_3_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_3_F_Inst_10__CF_Inst_U1 ( .A1(S_3_F_in2[1]), .A2(S_3_F_in1[3]), 
        .ZN(S_3_F_CF_Out[10]) );
  XNOR2_X1 S_3_F_Inst_11__CF_Inst_U2 ( .A(S_3_F_Inst_11__CF_Inst_n3), .B(
        S_3_F_in1[0]), .ZN(S_3_F_CF_Out[11]) );
  NAND2_X1 S_3_F_Inst_11__CF_Inst_U1 ( .A1(S_3_F_in3[1]), .A2(S_3_F_in1[3]), 
        .ZN(S_3_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_3_F_Inst_12__CF_Inst_U2 ( .A(S_3_F_Inst_12__CF_Inst_n3), .B(
        S_3_F_in2[0]), .ZN(S_3_F_CF_Out[12]) );
  NAND2_X1 S_3_F_Inst_12__CF_Inst_U1 ( .A1(S_3_F_in1[1]), .A2(S_3_F_in2[3]), 
        .ZN(S_3_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_3_F_Inst_13__CF_Inst_U2 ( .A1(S_3_F_in2[3]), .A2(
        S_3_F_Inst_13__CF_Inst_n3), .ZN(S_3_F_CF_Out[13]) );
  INV_X1 S_3_F_Inst_13__CF_Inst_U1 ( .A(S_3_F_in2[1]), .ZN(
        S_3_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_3_F_Inst_14__CF_Inst_U1 ( .A1(S_3_F_in3[1]), .A2(S_3_F_in2[3]), 
        .ZN(S_3_F_CF_Out[14]) );
  XNOR2_X1 S_3_F_Inst_15__CF_Inst_U2 ( .A(S_3_F_Inst_15__CF_Inst_n7), .B(
        S_3_F_in3[0]), .ZN(S_3_F_CF_Out[15]) );
  NOR2_X1 S_3_F_Inst_15__CF_Inst_U1 ( .A1(S_3_F_in1[1]), .A2(S_3_F_in3[3]), 
        .ZN(S_3_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_3_F_Inst_16__CF_Inst_U2 ( .A1(S_3_F_in3[3]), .A2(
        S_3_F_Inst_16__CF_Inst_n3), .ZN(S_3_F_CF_Out[16]) );
  INV_X1 S_3_F_Inst_16__CF_Inst_U1 ( .A(S_3_F_in2[1]), .ZN(
        S_3_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_3_F_Inst_17__CF_Inst_U2 ( .A1(S_3_F_in3[1]), .A2(
        S_3_F_Inst_17__CF_Inst_n3), .ZN(S_3_F_CF_Out[17]) );
  INV_X1 S_3_F_Inst_17__CF_Inst_U1 ( .A(S_3_F_in3[3]), .ZN(
        S_3_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_3_F_InstXOR_0__Compression1_U2 ( .A(
        S_3_F_InstXOR_0__Compression1_n3), .B(S_3_F_CF_Reg[2]), .ZN(
        S_3_F_q1[2]) );
  XNOR2_X1 S_3_F_InstXOR_0__Compression1_U1 ( .A(S_3_F_CF_Reg[0]), .B(
        S_3_F_CF_Reg[1]), .ZN(S_3_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_3_F_InstXOR_0__Compression2_U2 ( .A(
        S_3_F_InstXOR_0__Compression2_n3), .B(S_3_F_CF_Reg[5]), .ZN(
        S_3_F_q2[2]) );
  XNOR2_X1 S_3_F_InstXOR_0__Compression2_U1 ( .A(S_3_F_CF_Reg[3]), .B(
        S_3_F_CF_Reg[4]), .ZN(S_3_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_3_F_InstXOR_0__Compression3_U2 ( .A(
        S_3_F_InstXOR_0__Compression3_n3), .B(S_3_F_CF_Reg[8]), .ZN(
        S_3_F_q3[2]) );
  XNOR2_X1 S_3_F_InstXOR_0__Compression3_U1 ( .A(S_3_F_CF_Reg[6]), .B(
        S_3_F_CF_Reg[7]), .ZN(S_3_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_3_F_InstXOR_1__Compression1_U2 ( .A(
        S_3_F_InstXOR_1__Compression1_n3), .B(S_3_F_CF_Reg[11]), .ZN(
        S_3_F_q1[3]) );
  XNOR2_X1 S_3_F_InstXOR_1__Compression1_U1 ( .A(S_3_F_CF_Reg[9]), .B(
        S_3_F_CF_Reg[10]), .ZN(S_3_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_3_F_InstXOR_1__Compression2_U2 ( .A(
        S_3_F_InstXOR_1__Compression2_n3), .B(S_3_F_CF_Reg[14]), .ZN(
        S_3_F_q2[3]) );
  XNOR2_X1 S_3_F_InstXOR_1__Compression2_U1 ( .A(S_3_F_CF_Reg[12]), .B(
        S_3_F_CF_Reg[13]), .ZN(S_3_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_3_F_InstXOR_1__Compression3_U2 ( .A(
        S_3_F_InstXOR_1__Compression3_n3), .B(S_3_F_CF_Reg[17]), .ZN(
        S_3_F_q3[3]) );
  XNOR2_X1 S_3_F_InstXOR_1__Compression3_U1 ( .A(S_3_F_CF_Reg[15]), .B(
        S_3_F_CF_Reg[16]), .ZN(S_3_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_3_G_CF_Reg_reg_0_ ( .D(S_3_G_CF_Out[0]), .CK(CLK), .Q(
        S_3_G_CF_Reg[0]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_1_ ( .D(S_3_G_CF_Out[1]), .CK(CLK), .Q(
        S_3_G_CF_Reg[1]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_2_ ( .D(S_3_G_CF_Out[2]), .CK(CLK), .Q(
        S_3_G_CF_Reg[2]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_3_ ( .D(S_3_G_CF_Out[3]), .CK(CLK), .Q(
        S_3_G_CF_Reg[3]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_4_ ( .D(S_3_G_CF_Out[4]), .CK(CLK), .Q(
        S_3_G_CF_Reg[4]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_5_ ( .D(S_3_G_CF_Out[5]), .CK(CLK), .Q(
        S_3_G_CF_Reg[5]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_6_ ( .D(S_3_G_CF_Out[6]), .CK(CLK), .Q(
        S_3_G_CF_Reg[6]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_7_ ( .D(S_3_G_CF_Out[7]), .CK(CLK), .Q(
        S_3_G_CF_Reg[7]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_8_ ( .D(S_3_G_CF_Out[8]), .CK(CLK), .Q(
        S_3_G_CF_Reg[8]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_9_ ( .D(S_3_G_CF_Out[9]), .CK(CLK), .Q(
        S_3_G_CF_Reg[9]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_10_ ( .D(S_3_G_CF_Out[10]), .CK(CLK), .Q(
        S_3_G_CF_Reg[10]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_11_ ( .D(S_3_G_CF_Out[11]), .CK(CLK), .Q(
        S_3_G_CF_Reg[11]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_12_ ( .D(S_3_G_CF_Out[12]), .CK(CLK), .Q(
        S_3_G_CF_Reg[12]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_13_ ( .D(S_3_G_CF_Out[13]), .CK(CLK), .Q(
        S_3_G_CF_Reg[13]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_14_ ( .D(S_3_G_CF_Out[14]), .CK(CLK), .Q(
        S_3_G_CF_Reg[14]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_15_ ( .D(S_3_G_CF_Out[15]), .CK(CLK), .Q(
        S_3_G_CF_Reg[15]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_16_ ( .D(S_3_G_CF_Out[16]), .CK(CLK), .Q(
        S_3_G_CF_Reg[16]), .QN() );
  DFF_X1 S_3_G_CF_Reg_reg_17_ ( .D(S_3_G_CF_Out[17]), .CK(CLK), .Q(
        S_3_G_CF_Reg[17]), .QN() );
  DFF_X1 S_3_G_out1_reg_2_ ( .D(S_3_Rq1[2]), .CK(CLK), .Q(S_3_G_out1[2]), 
        .QN() );
  DFF_X1 S_3_G_out1_reg_3_ ( .D(S_3_Rq1[3]), .CK(CLK), .Q(S_3_G_out1[3]), 
        .QN() );
  DFF_X1 S_3_G_out2_reg_2_ ( .D(S_3_Rq2[2]), .CK(CLK), .Q(RF2_SHIFTROWS[2]), 
        .QN() );
  DFF_X1 S_3_G_out2_reg_3_ ( .D(S_3_Rq2[3]), .CK(CLK), .Q(RF2_SHIFTROWS[3]), 
        .QN() );
  DFF_X1 S_3_G_out3_reg_2_ ( .D(S_3_Rq3[2]), .CK(CLK), .Q(RF3_SHIFTROWS[2]), 
        .QN() );
  DFF_X1 S_3_G_out3_reg_3_ ( .D(S_3_Rq3[3]), .CK(CLK), .Q(RF3_SHIFTROWS[3]), 
        .QN() );
  AND2_X1 S_3_G_Inst_0__CF_Inst_U1 ( .A1(S_3_Rq1[1]), .A2(S_3_Rq1[3]), .ZN(
        S_3_G_CF_Out[0]) );
  NOR2_X1 S_3_G_Inst_1__CF_Inst_U2 ( .A1(S_3_Rq1[3]), .A2(
        S_3_G_Inst_1__CF_Inst_n3), .ZN(S_3_G_CF_Out[1]) );
  INV_X1 S_3_G_Inst_1__CF_Inst_U1 ( .A(S_3_Rq2[1]), .ZN(
        S_3_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_3_G_Inst_2__CF_Inst_U2 ( .A(S_3_G_Inst_2__CF_Inst_n3), .B(
        S_3_Rq2[0]), .ZN(S_3_G_CF_Out[2]) );
  NAND2_X1 S_3_G_Inst_2__CF_Inst_U1 ( .A1(S_3_Rq1[1]), .A2(S_3_Rq2[3]), .ZN(
        S_3_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_3_G_Inst_3__CF_Inst_U3 ( .A(S_3_Rq1[0]), .B(
        S_3_G_Inst_3__CF_Inst_n6), .ZN(S_3_G_CF_Out[3]) );
  NAND2_X1 S_3_G_Inst_3__CF_Inst_U2 ( .A1(S_3_Rq3[1]), .A2(
        S_3_G_Inst_3__CF_Inst_n5), .ZN(S_3_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_3_G_Inst_3__CF_Inst_U1 ( .A(S_3_Rq1[3]), .ZN(
        S_3_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_3_G_Inst_4__CF_Inst_U1 ( .A1(S_3_Rq2[1]), .A2(S_3_Rq2[3]), .ZN(
        S_3_G_CF_Out[4]) );
  OR2_X1 S_3_G_Inst_5__CF_Inst_U1 ( .A1(S_3_Rq3[3]), .A2(S_3_Rq2[1]), .ZN(
        S_3_G_CF_Out[5]) );
  AND2_X1 S_3_G_Inst_6__CF_Inst_U1 ( .A1(S_3_Rq3[1]), .A2(S_3_Rq2[3]), .ZN(
        S_3_G_CF_Out[6]) );
  XNOR2_X1 S_3_G_Inst_7__CF_Inst_U2 ( .A(S_3_G_Inst_7__CF_Inst_n3), .B(
        S_3_Rq3[0]), .ZN(S_3_G_CF_Out[7]) );
  NAND2_X1 S_3_G_Inst_7__CF_Inst_U1 ( .A1(S_3_Rq1[1]), .A2(S_3_Rq3[3]), .ZN(
        S_3_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_3_G_Inst_8__CF_Inst_U1 ( .A1(S_3_Rq3[3]), .A2(S_3_Rq3[1]), .ZN(
        S_3_G_CF_Out[8]) );
  NOR2_X1 S_3_G_Inst_9__CF_Inst_U2 ( .A1(S_3_Rq1[3]), .A2(
        S_3_G_Inst_9__CF_Inst_n3), .ZN(S_3_G_CF_Out[9]) );
  INV_X1 S_3_G_Inst_9__CF_Inst_U1 ( .A(S_3_Rq1[2]), .ZN(
        S_3_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_3_G_Inst_10__CF_Inst_U2 ( .A1(S_3_Rq2[2]), .A2(
        S_3_G_Inst_10__CF_Inst_n3), .ZN(S_3_G_CF_Out[10]) );
  INV_X1 S_3_G_Inst_10__CF_Inst_U1 ( .A(S_3_Rq1[3]), .ZN(
        S_3_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_3_G_Inst_11__CF_Inst_U3 ( .A(S_3_Rq1[1]), .B(
        S_3_G_Inst_11__CF_Inst_n6), .ZN(S_3_G_CF_Out[11]) );
  NAND2_X1 S_3_G_Inst_11__CF_Inst_U2 ( .A1(S_3_Rq1[3]), .A2(
        S_3_G_Inst_11__CF_Inst_n5), .ZN(S_3_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_3_G_Inst_11__CF_Inst_U1 ( .A(S_3_Rq3[2]), .ZN(
        S_3_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_3_G_Inst_12__CF_Inst_U2 ( .A1(S_3_Rq2[3]), .A2(
        S_3_G_Inst_12__CF_Inst_n3), .ZN(S_3_G_CF_Out[12]) );
  INV_X1 S_3_G_Inst_12__CF_Inst_U1 ( .A(S_3_Rq1[2]), .ZN(
        S_3_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_3_G_Inst_13__CF_Inst_U1 ( .A1(S_3_Rq2[2]), .A2(S_3_Rq2[3]), .ZN(
        S_3_G_CF_Out[13]) );
  XNOR2_X1 S_3_G_Inst_14__CF_Inst_U3 ( .A(S_3_Rq2[1]), .B(
        S_3_G_Inst_14__CF_Inst_n6), .ZN(S_3_G_CF_Out[14]) );
  NAND2_X1 S_3_G_Inst_14__CF_Inst_U2 ( .A1(S_3_Rq3[2]), .A2(
        S_3_G_Inst_14__CF_Inst_n5), .ZN(S_3_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_3_G_Inst_14__CF_Inst_U1 ( .A(S_3_Rq2[3]), .ZN(
        S_3_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_3_G_Inst_15__CF_Inst_U2 ( .A(S_3_G_Inst_15__CF_Inst_n3), .B(
        S_3_Rq3[1]), .ZN(S_3_G_CF_Out[15]) );
  NAND2_X1 S_3_G_Inst_15__CF_Inst_U1 ( .A1(S_3_Rq1[2]), .A2(S_3_Rq3[3]), .ZN(
        S_3_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_3_G_Inst_16__CF_Inst_U1 ( .A1(S_3_Rq2[2]), .A2(S_3_Rq3[3]), .ZN(
        S_3_G_CF_Out[16]) );
  NOR2_X1 S_3_G_Inst_17__CF_Inst_U2 ( .A1(S_3_Rq3[3]), .A2(
        S_3_G_Inst_17__CF_Inst_n3), .ZN(S_3_G_CF_Out[17]) );
  INV_X1 S_3_G_Inst_17__CF_Inst_U1 ( .A(S_3_Rq3[2]), .ZN(
        S_3_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_3_G_InstXOR_0__Compression1_U2 ( .A(
        S_3_G_InstXOR_0__Compression1_n3), .B(S_3_G_CF_Reg[2]), .ZN(
        S_3_G_out1[0]) );
  XNOR2_X1 S_3_G_InstXOR_0__Compression1_U1 ( .A(S_3_G_CF_Reg[0]), .B(
        S_3_G_CF_Reg[1]), .ZN(S_3_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_3_G_InstXOR_0__Compression2_U2 ( .A(
        S_3_G_InstXOR_0__Compression2_n3), .B(S_3_G_CF_Reg[5]), .ZN(
        RF2_SHIFTROWS[1]) );
  XNOR2_X1 S_3_G_InstXOR_0__Compression2_U1 ( .A(S_3_G_CF_Reg[3]), .B(
        S_3_G_CF_Reg[4]), .ZN(S_3_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_3_G_InstXOR_0__Compression3_U2 ( .A(
        S_3_G_InstXOR_0__Compression3_n3), .B(S_3_G_CF_Reg[8]), .ZN(
        RF3_SHIFTROWS[1]) );
  XNOR2_X1 S_3_G_InstXOR_0__Compression3_U1 ( .A(S_3_G_CF_Reg[6]), .B(
        S_3_G_CF_Reg[7]), .ZN(S_3_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_3_G_InstXOR_1__Compression1_U2 ( .A(
        S_3_G_InstXOR_1__Compression1_n3), .B(S_3_G_CF_Reg[11]), .ZN(
        S_3_G_out1[1]) );
  XNOR2_X1 S_3_G_InstXOR_1__Compression1_U1 ( .A(S_3_G_CF_Reg[9]), .B(
        S_3_G_CF_Reg[10]), .ZN(S_3_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_3_G_InstXOR_1__Compression2_U2 ( .A(
        S_3_G_InstXOR_1__Compression2_n3), .B(S_3_G_CF_Reg[14]), .ZN(
        RF2_SHIFTROWS[0]) );
  XNOR2_X1 S_3_G_InstXOR_1__Compression2_U1 ( .A(S_3_G_CF_Reg[12]), .B(
        S_3_G_CF_Reg[13]), .ZN(S_3_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_3_G_InstXOR_1__Compression3_U2 ( .A(
        S_3_G_InstXOR_1__Compression3_n3), .B(S_3_G_CF_Reg[17]), .ZN(
        RF3_SHIFTROWS[0]) );
  XNOR2_X1 S_3_G_InstXOR_1__Compression3_U1 ( .A(S_3_G_CF_Reg[15]), .B(
        S_3_G_CF_Reg[16]), .ZN(S_3_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_3_OutputAffine_U4 ( .A(S_3_G_out1[3]), .ZN(RF1_SHIFTROWS[3]) );
  INV_X1 S_3_OutputAffine_U3 ( .A(S_3_G_out1[2]), .ZN(RF1_SHIFTROWS[2]) );
  INV_X1 S_3_OutputAffine_U2 ( .A(S_3_G_out1[1]), .ZN(RF1_SHIFTROWS[0]) );
  INV_X1 S_3_OutputAffine_U1 ( .A(S_3_G_out1[0]), .ZN(RF1_SHIFTROWS[1]) );
  DFF_X1 S_4_Rq3_reg_0_ ( .D(S_4_q3[0]), .CK(CLK), .Q(S_4_Rq3[0]), .QN() );
  DFF_X1 S_4_Rq3_reg_1_ ( .D(S_4_q3[1]), .CK(CLK), .Q(S_4_Rq3[1]), .QN() );
  DFF_X1 S_4_Rq3_reg_2_ ( .D(S_4_q3[2]), .CK(CLK), .Q(S_4_Rq3[2]), .QN() );
  DFF_X1 S_4_Rq3_reg_3_ ( .D(S_4_q3[3]), .CK(CLK), .Q(S_4_Rq3[3]), .QN() );
  DFF_X1 S_4_Rq2_reg_0_ ( .D(S_4_q2[0]), .CK(CLK), .Q(S_4_Rq2[0]), .QN() );
  DFF_X1 S_4_Rq2_reg_1_ ( .D(S_4_q2[1]), .CK(CLK), .Q(S_4_Rq2[1]), .QN() );
  DFF_X1 S_4_Rq2_reg_2_ ( .D(S_4_q2[2]), .CK(CLK), .Q(S_4_Rq2[2]), .QN() );
  DFF_X1 S_4_Rq2_reg_3_ ( .D(S_4_q2[3]), .CK(CLK), .Q(S_4_Rq2[3]), .QN() );
  DFF_X1 S_4_Rq1_reg_0_ ( .D(S_4_q1[0]), .CK(CLK), .Q(S_4_Rq1[0]), .QN() );
  DFF_X1 S_4_Rq1_reg_1_ ( .D(S_4_q1[1]), .CK(CLK), .Q(S_4_Rq1[1]), .QN() );
  DFF_X1 S_4_Rq1_reg_2_ ( .D(S_4_q1[2]), .CK(CLK), .Q(S_4_Rq1[2]), .QN() );
  DFF_X1 S_4_Rq1_reg_3_ ( .D(S_4_q1[3]), .CK(CLK), .Q(S_4_Rq1[3]), .QN() );
  INV_X1 S_4_InputAffine_U4 ( .A(SUB_IN1[16]), .ZN(S_4_F_in1[0]) );
  INV_X1 S_4_InputAffine_U3 ( .A(SUB_IN1[18]), .ZN(S_4_F_in1[3]) );
  INV_X1 S_4_InputAffine_U2 ( .A(SUB_IN1[19]), .ZN(S_4_F_in1[1]) );
  INV_X1 S_4_InputAffine_U1 ( .A(SUB_IN1[17]), .ZN(S_4_F_in1[2]) );
  XNOR2_X1 S_4_F_U18 ( .A(S_4_F_n12), .B(FRESH[35]), .ZN(S_4_q3[3]) );
  XNOR2_X1 S_4_F_U17 ( .A(FRESH[34]), .B(S_4_F_q3[3]), .ZN(S_4_F_n12) );
  XNOR2_X1 S_4_F_U16 ( .A(S_4_F_n11), .B(FRESH[33]), .ZN(S_4_q3[2]) );
  XNOR2_X1 S_4_F_U15 ( .A(FRESH[32]), .B(S_4_F_q3[2]), .ZN(S_4_F_n11) );
  XOR2_X1 S_4_F_U14 ( .A(FRESH[35]), .B(S_4_F_q2[3]), .Z(S_4_q2[3]) );
  XOR2_X1 S_4_F_U13 ( .A(FRESH[33]), .B(S_4_F_q2[2]), .Z(S_4_q2[2]) );
  XOR2_X1 S_4_F_U12 ( .A(FRESH[34]), .B(S_4_F_q1[3]), .Z(S_4_q1[3]) );
  XOR2_X1 S_4_F_U11 ( .A(FRESH[32]), .B(S_4_F_q1[2]), .Z(S_4_q1[2]) );
  XNOR2_X1 S_4_F_U10 ( .A(S_4_F_n10), .B(FRESH[37]), .ZN(S_4_F_N5) );
  XNOR2_X1 S_4_F_U9 ( .A(S_4_F_in3[3]), .B(FRESH[36]), .ZN(S_4_F_n10) );
  XOR2_X1 S_4_F_U8 ( .A(FRESH[37]), .B(S_4_F_in2[3]), .Z(S_4_F_N4) );
  XOR2_X1 S_4_F_U7 ( .A(FRESH[36]), .B(S_4_F_in1[3]), .Z(S_4_F_N3) );
  XNOR2_X1 S_4_F_U6 ( .A(S_4_F_n9), .B(FRESH[39]), .ZN(S_4_F_N2) );
  XNOR2_X1 S_4_F_U5 ( .A(S_4_F_in3[2]), .B(FRESH[38]), .ZN(S_4_F_n9) );
  XOR2_X1 S_4_F_U4 ( .A(FRESH[39]), .B(S_4_F_in2[2]), .Z(S_4_F_N1) );
  XOR2_X1 S_4_F_U3 ( .A(FRESH[38]), .B(S_4_F_in1[2]), .Z(S_4_F_N0) );
  DFF_X1 S_4_F_CF_Reg_reg_0_ ( .D(S_4_F_CF_Out[0]), .CK(CLK), .Q(
        S_4_F_CF_Reg[0]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_1_ ( .D(S_4_F_CF_Out[1]), .CK(CLK), .Q(
        S_4_F_CF_Reg[1]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_2_ ( .D(S_4_F_CF_Out[2]), .CK(CLK), .Q(
        S_4_F_CF_Reg[2]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_3_ ( .D(S_4_F_CF_Out[3]), .CK(CLK), .Q(
        S_4_F_CF_Reg[3]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_4_ ( .D(S_4_F_CF_Out[4]), .CK(CLK), .Q(
        S_4_F_CF_Reg[4]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_5_ ( .D(S_4_F_CF_Out[5]), .CK(CLK), .Q(
        S_4_F_CF_Reg[5]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_6_ ( .D(S_4_F_CF_Out[6]), .CK(CLK), .Q(
        S_4_F_CF_Reg[6]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_7_ ( .D(S_4_F_CF_Out[7]), .CK(CLK), .Q(
        S_4_F_CF_Reg[7]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_8_ ( .D(S_4_F_CF_Out[8]), .CK(CLK), .Q(
        S_4_F_CF_Reg[8]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_9_ ( .D(S_4_F_CF_Out[9]), .CK(CLK), .Q(
        S_4_F_CF_Reg[9]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_10_ ( .D(S_4_F_CF_Out[10]), .CK(CLK), .Q(
        S_4_F_CF_Reg[10]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_11_ ( .D(S_4_F_CF_Out[11]), .CK(CLK), .Q(
        S_4_F_CF_Reg[11]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_12_ ( .D(S_4_F_CF_Out[12]), .CK(CLK), .Q(
        S_4_F_CF_Reg[12]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_13_ ( .D(S_4_F_CF_Out[13]), .CK(CLK), .Q(
        S_4_F_CF_Reg[13]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_14_ ( .D(S_4_F_CF_Out[14]), .CK(CLK), .Q(
        S_4_F_CF_Reg[14]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_15_ ( .D(S_4_F_CF_Out[15]), .CK(CLK), .Q(
        S_4_F_CF_Reg[15]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_16_ ( .D(S_4_F_CF_Out[16]), .CK(CLK), .Q(
        S_4_F_CF_Reg[16]), .QN() );
  DFF_X1 S_4_F_CF_Reg_reg_17_ ( .D(S_4_F_CF_Out[17]), .CK(CLK), .Q(
        S_4_F_CF_Reg[17]), .QN() );
  DFF_X1 S_4_F_out2_reg_0_ ( .D(S_4_F_N4), .CK(CLK), .Q(S_4_q2[0]), .QN() );
  DFF_X1 S_4_F_out2_reg_1_ ( .D(S_4_F_N1), .CK(CLK), .Q(S_4_q2[1]), .QN() );
  DFF_X1 S_4_F_out3_reg_0_ ( .D(S_4_F_N5), .CK(CLK), .Q(S_4_q3[0]), .QN() );
  DFF_X1 S_4_F_out3_reg_1_ ( .D(S_4_F_N2), .CK(CLK), .Q(S_4_q3[1]), .QN() );
  DFF_X1 S_4_F_out1_reg_0_ ( .D(S_4_F_N3), .CK(CLK), .Q(S_4_q1[0]), .QN() );
  DFF_X1 S_4_F_out1_reg_1_ ( .D(S_4_F_N0), .CK(CLK), .Q(S_4_q1[1]), .QN() );
  NOR2_X1 S_4_F_Inst_0__CF_Inst_U2 ( .A1(S_4_F_in1[2]), .A2(
        S_4_F_Inst_0__CF_Inst_n3), .ZN(S_4_F_CF_Out[0]) );
  INV_X1 S_4_F_Inst_0__CF_Inst_U1 ( .A(S_4_F_in1[3]), .ZN(
        S_4_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_4_F_Inst_1__CF_Inst_U2 ( .A(S_4_F_Inst_1__CF_Inst_n3), .B(
        S_4_F_in1[1]), .ZN(S_4_F_CF_Out[1]) );
  NAND2_X1 S_4_F_Inst_1__CF_Inst_U1 ( .A1(S_4_F_in2[2]), .A2(S_4_F_in1[3]), 
        .ZN(S_4_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_4_F_Inst_2__CF_Inst_U1 ( .A1(S_4_F_in1[3]), .A2(S_4_F_in3[2]), .ZN(
        S_4_F_CF_Out[2]) );
  NOR2_X1 S_4_F_Inst_3__CF_Inst_U2 ( .A1(S_4_F_in2[3]), .A2(
        S_4_F_Inst_3__CF_Inst_n3), .ZN(S_4_F_CF_Out[3]) );
  INV_X1 S_4_F_Inst_3__CF_Inst_U1 ( .A(S_4_F_in1[2]), .ZN(
        S_4_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_4_F_Inst_4__CF_Inst_U2 ( .A(S_4_F_Inst_4__CF_Inst_n3), .B(
        S_4_F_in2[1]), .ZN(S_4_F_CF_Out[4]) );
  NAND2_X1 S_4_F_Inst_4__CF_Inst_U1 ( .A1(S_4_F_in2[2]), .A2(S_4_F_in2[3]), 
        .ZN(S_4_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_4_F_Inst_5__CF_Inst_U1 ( .A1(S_4_F_in3[2]), .A2(S_4_F_in2[3]), 
        .ZN(S_4_F_CF_Out[5]) );
  XNOR2_X1 S_4_F_Inst_6__CF_Inst_U2 ( .A(S_4_F_Inst_6__CF_Inst_n7), .B(
        S_4_F_in3[1]), .ZN(S_4_F_CF_Out[6]) );
  NOR2_X1 S_4_F_Inst_6__CF_Inst_U1 ( .A1(S_4_F_in1[2]), .A2(S_4_F_in3[3]), 
        .ZN(S_4_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_4_F_Inst_7__CF_Inst_U1 ( .A1(S_4_F_in2[2]), .A2(S_4_F_in3[3]), 
        .ZN(S_4_F_CF_Out[7]) );
  OR2_X1 S_4_F_Inst_8__CF_Inst_U1 ( .A1(S_4_F_in3[3]), .A2(S_4_F_in3[2]), .ZN(
        S_4_F_CF_Out[8]) );
  NOR2_X1 S_4_F_Inst_9__CF_Inst_U2 ( .A1(S_4_F_in1[3]), .A2(
        S_4_F_Inst_9__CF_Inst_n3), .ZN(S_4_F_CF_Out[9]) );
  INV_X1 S_4_F_Inst_9__CF_Inst_U1 ( .A(S_4_F_in1[1]), .ZN(
        S_4_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_4_F_Inst_10__CF_Inst_U1 ( .A1(S_4_F_in2[1]), .A2(S_4_F_in1[3]), 
        .ZN(S_4_F_CF_Out[10]) );
  XNOR2_X1 S_4_F_Inst_11__CF_Inst_U2 ( .A(S_4_F_Inst_11__CF_Inst_n3), .B(
        S_4_F_in1[0]), .ZN(S_4_F_CF_Out[11]) );
  NAND2_X1 S_4_F_Inst_11__CF_Inst_U1 ( .A1(S_4_F_in3[1]), .A2(S_4_F_in1[3]), 
        .ZN(S_4_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_4_F_Inst_12__CF_Inst_U2 ( .A(S_4_F_Inst_12__CF_Inst_n3), .B(
        S_4_F_in2[0]), .ZN(S_4_F_CF_Out[12]) );
  NAND2_X1 S_4_F_Inst_12__CF_Inst_U1 ( .A1(S_4_F_in1[1]), .A2(S_4_F_in2[3]), 
        .ZN(S_4_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_4_F_Inst_13__CF_Inst_U2 ( .A1(S_4_F_in2[3]), .A2(
        S_4_F_Inst_13__CF_Inst_n3), .ZN(S_4_F_CF_Out[13]) );
  INV_X1 S_4_F_Inst_13__CF_Inst_U1 ( .A(S_4_F_in2[1]), .ZN(
        S_4_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_4_F_Inst_14__CF_Inst_U1 ( .A1(S_4_F_in3[1]), .A2(S_4_F_in2[3]), 
        .ZN(S_4_F_CF_Out[14]) );
  XNOR2_X1 S_4_F_Inst_15__CF_Inst_U2 ( .A(S_4_F_Inst_15__CF_Inst_n7), .B(
        S_4_F_in3[0]), .ZN(S_4_F_CF_Out[15]) );
  NOR2_X1 S_4_F_Inst_15__CF_Inst_U1 ( .A1(S_4_F_in1[1]), .A2(S_4_F_in3[3]), 
        .ZN(S_4_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_4_F_Inst_16__CF_Inst_U2 ( .A1(S_4_F_in3[3]), .A2(
        S_4_F_Inst_16__CF_Inst_n3), .ZN(S_4_F_CF_Out[16]) );
  INV_X1 S_4_F_Inst_16__CF_Inst_U1 ( .A(S_4_F_in2[1]), .ZN(
        S_4_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_4_F_Inst_17__CF_Inst_U2 ( .A1(S_4_F_in3[1]), .A2(
        S_4_F_Inst_17__CF_Inst_n3), .ZN(S_4_F_CF_Out[17]) );
  INV_X1 S_4_F_Inst_17__CF_Inst_U1 ( .A(S_4_F_in3[3]), .ZN(
        S_4_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_4_F_InstXOR_0__Compression1_U2 ( .A(
        S_4_F_InstXOR_0__Compression1_n3), .B(S_4_F_CF_Reg[2]), .ZN(
        S_4_F_q1[2]) );
  XNOR2_X1 S_4_F_InstXOR_0__Compression1_U1 ( .A(S_4_F_CF_Reg[0]), .B(
        S_4_F_CF_Reg[1]), .ZN(S_4_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_4_F_InstXOR_0__Compression2_U2 ( .A(
        S_4_F_InstXOR_0__Compression2_n3), .B(S_4_F_CF_Reg[5]), .ZN(
        S_4_F_q2[2]) );
  XNOR2_X1 S_4_F_InstXOR_0__Compression2_U1 ( .A(S_4_F_CF_Reg[3]), .B(
        S_4_F_CF_Reg[4]), .ZN(S_4_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_4_F_InstXOR_0__Compression3_U2 ( .A(
        S_4_F_InstXOR_0__Compression3_n3), .B(S_4_F_CF_Reg[8]), .ZN(
        S_4_F_q3[2]) );
  XNOR2_X1 S_4_F_InstXOR_0__Compression3_U1 ( .A(S_4_F_CF_Reg[6]), .B(
        S_4_F_CF_Reg[7]), .ZN(S_4_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_4_F_InstXOR_1__Compression1_U2 ( .A(
        S_4_F_InstXOR_1__Compression1_n3), .B(S_4_F_CF_Reg[11]), .ZN(
        S_4_F_q1[3]) );
  XNOR2_X1 S_4_F_InstXOR_1__Compression1_U1 ( .A(S_4_F_CF_Reg[9]), .B(
        S_4_F_CF_Reg[10]), .ZN(S_4_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_4_F_InstXOR_1__Compression2_U2 ( .A(
        S_4_F_InstXOR_1__Compression2_n3), .B(S_4_F_CF_Reg[14]), .ZN(
        S_4_F_q2[3]) );
  XNOR2_X1 S_4_F_InstXOR_1__Compression2_U1 ( .A(S_4_F_CF_Reg[12]), .B(
        S_4_F_CF_Reg[13]), .ZN(S_4_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_4_F_InstXOR_1__Compression3_U2 ( .A(
        S_4_F_InstXOR_1__Compression3_n3), .B(S_4_F_CF_Reg[17]), .ZN(
        S_4_F_q3[3]) );
  XNOR2_X1 S_4_F_InstXOR_1__Compression3_U1 ( .A(S_4_F_CF_Reg[15]), .B(
        S_4_F_CF_Reg[16]), .ZN(S_4_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_4_G_CF_Reg_reg_0_ ( .D(S_4_G_CF_Out[0]), .CK(CLK), .Q(
        S_4_G_CF_Reg[0]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_1_ ( .D(S_4_G_CF_Out[1]), .CK(CLK), .Q(
        S_4_G_CF_Reg[1]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_2_ ( .D(S_4_G_CF_Out[2]), .CK(CLK), .Q(
        S_4_G_CF_Reg[2]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_3_ ( .D(S_4_G_CF_Out[3]), .CK(CLK), .Q(
        S_4_G_CF_Reg[3]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_4_ ( .D(S_4_G_CF_Out[4]), .CK(CLK), .Q(
        S_4_G_CF_Reg[4]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_5_ ( .D(S_4_G_CF_Out[5]), .CK(CLK), .Q(
        S_4_G_CF_Reg[5]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_6_ ( .D(S_4_G_CF_Out[6]), .CK(CLK), .Q(
        S_4_G_CF_Reg[6]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_7_ ( .D(S_4_G_CF_Out[7]), .CK(CLK), .Q(
        S_4_G_CF_Reg[7]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_8_ ( .D(S_4_G_CF_Out[8]), .CK(CLK), .Q(
        S_4_G_CF_Reg[8]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_9_ ( .D(S_4_G_CF_Out[9]), .CK(CLK), .Q(
        S_4_G_CF_Reg[9]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_10_ ( .D(S_4_G_CF_Out[10]), .CK(CLK), .Q(
        S_4_G_CF_Reg[10]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_11_ ( .D(S_4_G_CF_Out[11]), .CK(CLK), .Q(
        S_4_G_CF_Reg[11]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_12_ ( .D(S_4_G_CF_Out[12]), .CK(CLK), .Q(
        S_4_G_CF_Reg[12]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_13_ ( .D(S_4_G_CF_Out[13]), .CK(CLK), .Q(
        S_4_G_CF_Reg[13]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_14_ ( .D(S_4_G_CF_Out[14]), .CK(CLK), .Q(
        S_4_G_CF_Reg[14]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_15_ ( .D(S_4_G_CF_Out[15]), .CK(CLK), .Q(
        S_4_G_CF_Reg[15]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_16_ ( .D(S_4_G_CF_Out[16]), .CK(CLK), .Q(
        S_4_G_CF_Reg[16]), .QN() );
  DFF_X1 S_4_G_CF_Reg_reg_17_ ( .D(S_4_G_CF_Out[17]), .CK(CLK), .Q(
        S_4_G_CF_Reg[17]), .QN() );
  DFF_X1 S_4_G_out1_reg_2_ ( .D(S_4_Rq1[2]), .CK(CLK), .Q(S_4_G_out1[2]), 
        .QN() );
  DFF_X1 S_4_G_out1_reg_3_ ( .D(S_4_Rq1[3]), .CK(CLK), .Q(S_4_G_out1[3]), 
        .QN() );
  DFF_X1 S_4_G_out2_reg_2_ ( .D(S_4_Rq2[2]), .CK(CLK), .Q(RF2_SHIFTROWS[26]), 
        .QN() );
  DFF_X1 S_4_G_out2_reg_3_ ( .D(S_4_Rq2[3]), .CK(CLK), .Q(RF2_SHIFTROWS[27]), 
        .QN() );
  DFF_X1 S_4_G_out3_reg_2_ ( .D(S_4_Rq3[2]), .CK(CLK), .Q(RF3_SHIFTROWS[26]), 
        .QN() );
  DFF_X1 S_4_G_out3_reg_3_ ( .D(S_4_Rq3[3]), .CK(CLK), .Q(RF3_SHIFTROWS[27]), 
        .QN() );
  AND2_X1 S_4_G_Inst_0__CF_Inst_U1 ( .A1(S_4_Rq1[1]), .A2(S_4_Rq1[3]), .ZN(
        S_4_G_CF_Out[0]) );
  NOR2_X1 S_4_G_Inst_1__CF_Inst_U2 ( .A1(S_4_Rq1[3]), .A2(
        S_4_G_Inst_1__CF_Inst_n3), .ZN(S_4_G_CF_Out[1]) );
  INV_X1 S_4_G_Inst_1__CF_Inst_U1 ( .A(S_4_Rq2[1]), .ZN(
        S_4_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_4_G_Inst_2__CF_Inst_U2 ( .A(S_4_G_Inst_2__CF_Inst_n3), .B(
        S_4_Rq2[0]), .ZN(S_4_G_CF_Out[2]) );
  NAND2_X1 S_4_G_Inst_2__CF_Inst_U1 ( .A1(S_4_Rq1[1]), .A2(S_4_Rq2[3]), .ZN(
        S_4_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_4_G_Inst_3__CF_Inst_U3 ( .A(S_4_Rq1[0]), .B(
        S_4_G_Inst_3__CF_Inst_n6), .ZN(S_4_G_CF_Out[3]) );
  NAND2_X1 S_4_G_Inst_3__CF_Inst_U2 ( .A1(S_4_Rq3[1]), .A2(
        S_4_G_Inst_3__CF_Inst_n5), .ZN(S_4_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_4_G_Inst_3__CF_Inst_U1 ( .A(S_4_Rq1[3]), .ZN(
        S_4_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_4_G_Inst_4__CF_Inst_U1 ( .A1(S_4_Rq2[1]), .A2(S_4_Rq2[3]), .ZN(
        S_4_G_CF_Out[4]) );
  OR2_X1 S_4_G_Inst_5__CF_Inst_U1 ( .A1(S_4_Rq3[3]), .A2(S_4_Rq2[1]), .ZN(
        S_4_G_CF_Out[5]) );
  AND2_X1 S_4_G_Inst_6__CF_Inst_U1 ( .A1(S_4_Rq3[1]), .A2(S_4_Rq2[3]), .ZN(
        S_4_G_CF_Out[6]) );
  XNOR2_X1 S_4_G_Inst_7__CF_Inst_U2 ( .A(S_4_G_Inst_7__CF_Inst_n3), .B(
        S_4_Rq3[0]), .ZN(S_4_G_CF_Out[7]) );
  NAND2_X1 S_4_G_Inst_7__CF_Inst_U1 ( .A1(S_4_Rq1[1]), .A2(S_4_Rq3[3]), .ZN(
        S_4_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_4_G_Inst_8__CF_Inst_U1 ( .A1(S_4_Rq3[3]), .A2(S_4_Rq3[1]), .ZN(
        S_4_G_CF_Out[8]) );
  NOR2_X1 S_4_G_Inst_9__CF_Inst_U2 ( .A1(S_4_Rq1[3]), .A2(
        S_4_G_Inst_9__CF_Inst_n3), .ZN(S_4_G_CF_Out[9]) );
  INV_X1 S_4_G_Inst_9__CF_Inst_U1 ( .A(S_4_Rq1[2]), .ZN(
        S_4_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_4_G_Inst_10__CF_Inst_U2 ( .A1(S_4_Rq2[2]), .A2(
        S_4_G_Inst_10__CF_Inst_n3), .ZN(S_4_G_CF_Out[10]) );
  INV_X1 S_4_G_Inst_10__CF_Inst_U1 ( .A(S_4_Rq1[3]), .ZN(
        S_4_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_4_G_Inst_11__CF_Inst_U3 ( .A(S_4_Rq1[1]), .B(
        S_4_G_Inst_11__CF_Inst_n6), .ZN(S_4_G_CF_Out[11]) );
  NAND2_X1 S_4_G_Inst_11__CF_Inst_U2 ( .A1(S_4_Rq1[3]), .A2(
        S_4_G_Inst_11__CF_Inst_n5), .ZN(S_4_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_4_G_Inst_11__CF_Inst_U1 ( .A(S_4_Rq3[2]), .ZN(
        S_4_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_4_G_Inst_12__CF_Inst_U2 ( .A1(S_4_Rq2[3]), .A2(
        S_4_G_Inst_12__CF_Inst_n3), .ZN(S_4_G_CF_Out[12]) );
  INV_X1 S_4_G_Inst_12__CF_Inst_U1 ( .A(S_4_Rq1[2]), .ZN(
        S_4_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_4_G_Inst_13__CF_Inst_U1 ( .A1(S_4_Rq2[2]), .A2(S_4_Rq2[3]), .ZN(
        S_4_G_CF_Out[13]) );
  XNOR2_X1 S_4_G_Inst_14__CF_Inst_U3 ( .A(S_4_Rq2[1]), .B(
        S_4_G_Inst_14__CF_Inst_n6), .ZN(S_4_G_CF_Out[14]) );
  NAND2_X1 S_4_G_Inst_14__CF_Inst_U2 ( .A1(S_4_Rq3[2]), .A2(
        S_4_G_Inst_14__CF_Inst_n5), .ZN(S_4_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_4_G_Inst_14__CF_Inst_U1 ( .A(S_4_Rq2[3]), .ZN(
        S_4_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_4_G_Inst_15__CF_Inst_U2 ( .A(S_4_G_Inst_15__CF_Inst_n3), .B(
        S_4_Rq3[1]), .ZN(S_4_G_CF_Out[15]) );
  NAND2_X1 S_4_G_Inst_15__CF_Inst_U1 ( .A1(S_4_Rq1[2]), .A2(S_4_Rq3[3]), .ZN(
        S_4_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_4_G_Inst_16__CF_Inst_U1 ( .A1(S_4_Rq2[2]), .A2(S_4_Rq3[3]), .ZN(
        S_4_G_CF_Out[16]) );
  NOR2_X1 S_4_G_Inst_17__CF_Inst_U2 ( .A1(S_4_Rq3[3]), .A2(
        S_4_G_Inst_17__CF_Inst_n3), .ZN(S_4_G_CF_Out[17]) );
  INV_X1 S_4_G_Inst_17__CF_Inst_U1 ( .A(S_4_Rq3[2]), .ZN(
        S_4_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_4_G_InstXOR_0__Compression1_U2 ( .A(
        S_4_G_InstXOR_0__Compression1_n3), .B(S_4_G_CF_Reg[2]), .ZN(
        S_4_G_out1[0]) );
  XNOR2_X1 S_4_G_InstXOR_0__Compression1_U1 ( .A(S_4_G_CF_Reg[0]), .B(
        S_4_G_CF_Reg[1]), .ZN(S_4_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_4_G_InstXOR_0__Compression2_U2 ( .A(
        S_4_G_InstXOR_0__Compression2_n3), .B(S_4_G_CF_Reg[5]), .ZN(
        RF2_SHIFTROWS[25]) );
  XNOR2_X1 S_4_G_InstXOR_0__Compression2_U1 ( .A(S_4_G_CF_Reg[3]), .B(
        S_4_G_CF_Reg[4]), .ZN(S_4_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_4_G_InstXOR_0__Compression3_U2 ( .A(
        S_4_G_InstXOR_0__Compression3_n3), .B(S_4_G_CF_Reg[8]), .ZN(
        RF3_SHIFTROWS[25]) );
  XNOR2_X1 S_4_G_InstXOR_0__Compression3_U1 ( .A(S_4_G_CF_Reg[6]), .B(
        S_4_G_CF_Reg[7]), .ZN(S_4_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_4_G_InstXOR_1__Compression1_U2 ( .A(
        S_4_G_InstXOR_1__Compression1_n3), .B(S_4_G_CF_Reg[11]), .ZN(
        S_4_G_out1[1]) );
  XNOR2_X1 S_4_G_InstXOR_1__Compression1_U1 ( .A(S_4_G_CF_Reg[9]), .B(
        S_4_G_CF_Reg[10]), .ZN(S_4_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_4_G_InstXOR_1__Compression2_U2 ( .A(
        S_4_G_InstXOR_1__Compression2_n3), .B(S_4_G_CF_Reg[14]), .ZN(
        RF2_SHIFTROWS[24]) );
  XNOR2_X1 S_4_G_InstXOR_1__Compression2_U1 ( .A(S_4_G_CF_Reg[12]), .B(
        S_4_G_CF_Reg[13]), .ZN(S_4_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_4_G_InstXOR_1__Compression3_U2 ( .A(
        S_4_G_InstXOR_1__Compression3_n3), .B(S_4_G_CF_Reg[17]), .ZN(
        RF3_SHIFTROWS[24]) );
  XNOR2_X1 S_4_G_InstXOR_1__Compression3_U1 ( .A(S_4_G_CF_Reg[15]), .B(
        S_4_G_CF_Reg[16]), .ZN(S_4_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_4_OutputAffine_U4 ( .A(S_4_G_out1[3]), .ZN(RF1_SHIFTROWS[27]) );
  INV_X1 S_4_OutputAffine_U3 ( .A(S_4_G_out1[2]), .ZN(RF1_SHIFTROWS[26]) );
  INV_X1 S_4_OutputAffine_U2 ( .A(S_4_G_out1[1]), .ZN(RF1_SHIFTROWS[24]) );
  INV_X1 S_4_OutputAffine_U1 ( .A(S_4_G_out1[0]), .ZN(RF1_SHIFTROWS[25]) );
  DFF_X1 S_5_Rq3_reg_0_ ( .D(S_5_q3[0]), .CK(CLK), .Q(S_5_Rq3[0]), .QN() );
  DFF_X1 S_5_Rq3_reg_1_ ( .D(S_5_q3[1]), .CK(CLK), .Q(S_5_Rq3[1]), .QN() );
  DFF_X1 S_5_Rq3_reg_2_ ( .D(S_5_q3[2]), .CK(CLK), .Q(S_5_Rq3[2]), .QN() );
  DFF_X1 S_5_Rq3_reg_3_ ( .D(S_5_q3[3]), .CK(CLK), .Q(S_5_Rq3[3]), .QN() );
  DFF_X1 S_5_Rq2_reg_0_ ( .D(S_5_q2[0]), .CK(CLK), .Q(S_5_Rq2[0]), .QN() );
  DFF_X1 S_5_Rq2_reg_1_ ( .D(S_5_q2[1]), .CK(CLK), .Q(S_5_Rq2[1]), .QN() );
  DFF_X1 S_5_Rq2_reg_2_ ( .D(S_5_q2[2]), .CK(CLK), .Q(S_5_Rq2[2]), .QN() );
  DFF_X1 S_5_Rq2_reg_3_ ( .D(S_5_q2[3]), .CK(CLK), .Q(S_5_Rq2[3]), .QN() );
  DFF_X1 S_5_Rq1_reg_0_ ( .D(S_5_q1[0]), .CK(CLK), .Q(S_5_Rq1[0]), .QN() );
  DFF_X1 S_5_Rq1_reg_1_ ( .D(S_5_q1[1]), .CK(CLK), .Q(S_5_Rq1[1]), .QN() );
  DFF_X1 S_5_Rq1_reg_2_ ( .D(S_5_q1[2]), .CK(CLK), .Q(S_5_Rq1[2]), .QN() );
  DFF_X1 S_5_Rq1_reg_3_ ( .D(S_5_q1[3]), .CK(CLK), .Q(S_5_Rq1[3]), .QN() );
  INV_X1 S_5_InputAffine_U4 ( .A(SUB_IN1[20]), .ZN(S_5_F_in1[0]) );
  INV_X1 S_5_InputAffine_U3 ( .A(SUB_IN1[22]), .ZN(S_5_F_in1[3]) );
  INV_X1 S_5_InputAffine_U2 ( .A(SUB_IN1[23]), .ZN(S_5_F_in1[1]) );
  INV_X1 S_5_InputAffine_U1 ( .A(SUB_IN1[21]), .ZN(S_5_F_in1[2]) );
  XNOR2_X1 S_5_F_U18 ( .A(S_5_F_n12), .B(FRESH[43]), .ZN(S_5_q3[3]) );
  XNOR2_X1 S_5_F_U17 ( .A(FRESH[42]), .B(S_5_F_q3[3]), .ZN(S_5_F_n12) );
  XNOR2_X1 S_5_F_U16 ( .A(S_5_F_n11), .B(FRESH[41]), .ZN(S_5_q3[2]) );
  XNOR2_X1 S_5_F_U15 ( .A(FRESH[40]), .B(S_5_F_q3[2]), .ZN(S_5_F_n11) );
  XOR2_X1 S_5_F_U14 ( .A(FRESH[43]), .B(S_5_F_q2[3]), .Z(S_5_q2[3]) );
  XOR2_X1 S_5_F_U13 ( .A(FRESH[41]), .B(S_5_F_q2[2]), .Z(S_5_q2[2]) );
  XOR2_X1 S_5_F_U12 ( .A(FRESH[42]), .B(S_5_F_q1[3]), .Z(S_5_q1[3]) );
  XOR2_X1 S_5_F_U11 ( .A(FRESH[40]), .B(S_5_F_q1[2]), .Z(S_5_q1[2]) );
  XNOR2_X1 S_5_F_U10 ( .A(S_5_F_n10), .B(FRESH[45]), .ZN(S_5_F_N5) );
  XNOR2_X1 S_5_F_U9 ( .A(S_5_F_in3[3]), .B(FRESH[44]), .ZN(S_5_F_n10) );
  XOR2_X1 S_5_F_U8 ( .A(FRESH[45]), .B(S_5_F_in2[3]), .Z(S_5_F_N4) );
  XOR2_X1 S_5_F_U7 ( .A(FRESH[44]), .B(S_5_F_in1[3]), .Z(S_5_F_N3) );
  XNOR2_X1 S_5_F_U6 ( .A(S_5_F_n9), .B(FRESH[47]), .ZN(S_5_F_N2) );
  XNOR2_X1 S_5_F_U5 ( .A(S_5_F_in3[2]), .B(FRESH[46]), .ZN(S_5_F_n9) );
  XOR2_X1 S_5_F_U4 ( .A(FRESH[47]), .B(S_5_F_in2[2]), .Z(S_5_F_N1) );
  XOR2_X1 S_5_F_U3 ( .A(FRESH[46]), .B(S_5_F_in1[2]), .Z(S_5_F_N0) );
  DFF_X1 S_5_F_CF_Reg_reg_0_ ( .D(S_5_F_CF_Out[0]), .CK(CLK), .Q(
        S_5_F_CF_Reg[0]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_1_ ( .D(S_5_F_CF_Out[1]), .CK(CLK), .Q(
        S_5_F_CF_Reg[1]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_2_ ( .D(S_5_F_CF_Out[2]), .CK(CLK), .Q(
        S_5_F_CF_Reg[2]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_3_ ( .D(S_5_F_CF_Out[3]), .CK(CLK), .Q(
        S_5_F_CF_Reg[3]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_4_ ( .D(S_5_F_CF_Out[4]), .CK(CLK), .Q(
        S_5_F_CF_Reg[4]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_5_ ( .D(S_5_F_CF_Out[5]), .CK(CLK), .Q(
        S_5_F_CF_Reg[5]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_6_ ( .D(S_5_F_CF_Out[6]), .CK(CLK), .Q(
        S_5_F_CF_Reg[6]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_7_ ( .D(S_5_F_CF_Out[7]), .CK(CLK), .Q(
        S_5_F_CF_Reg[7]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_8_ ( .D(S_5_F_CF_Out[8]), .CK(CLK), .Q(
        S_5_F_CF_Reg[8]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_9_ ( .D(S_5_F_CF_Out[9]), .CK(CLK), .Q(
        S_5_F_CF_Reg[9]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_10_ ( .D(S_5_F_CF_Out[10]), .CK(CLK), .Q(
        S_5_F_CF_Reg[10]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_11_ ( .D(S_5_F_CF_Out[11]), .CK(CLK), .Q(
        S_5_F_CF_Reg[11]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_12_ ( .D(S_5_F_CF_Out[12]), .CK(CLK), .Q(
        S_5_F_CF_Reg[12]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_13_ ( .D(S_5_F_CF_Out[13]), .CK(CLK), .Q(
        S_5_F_CF_Reg[13]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_14_ ( .D(S_5_F_CF_Out[14]), .CK(CLK), .Q(
        S_5_F_CF_Reg[14]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_15_ ( .D(S_5_F_CF_Out[15]), .CK(CLK), .Q(
        S_5_F_CF_Reg[15]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_16_ ( .D(S_5_F_CF_Out[16]), .CK(CLK), .Q(
        S_5_F_CF_Reg[16]), .QN() );
  DFF_X1 S_5_F_CF_Reg_reg_17_ ( .D(S_5_F_CF_Out[17]), .CK(CLK), .Q(
        S_5_F_CF_Reg[17]), .QN() );
  DFF_X1 S_5_F_out2_reg_0_ ( .D(S_5_F_N4), .CK(CLK), .Q(S_5_q2[0]), .QN() );
  DFF_X1 S_5_F_out2_reg_1_ ( .D(S_5_F_N1), .CK(CLK), .Q(S_5_q2[1]), .QN() );
  DFF_X1 S_5_F_out3_reg_0_ ( .D(S_5_F_N5), .CK(CLK), .Q(S_5_q3[0]), .QN() );
  DFF_X1 S_5_F_out3_reg_1_ ( .D(S_5_F_N2), .CK(CLK), .Q(S_5_q3[1]), .QN() );
  DFF_X1 S_5_F_out1_reg_0_ ( .D(S_5_F_N3), .CK(CLK), .Q(S_5_q1[0]), .QN() );
  DFF_X1 S_5_F_out1_reg_1_ ( .D(S_5_F_N0), .CK(CLK), .Q(S_5_q1[1]), .QN() );
  NOR2_X1 S_5_F_Inst_0__CF_Inst_U2 ( .A1(S_5_F_in1[2]), .A2(
        S_5_F_Inst_0__CF_Inst_n3), .ZN(S_5_F_CF_Out[0]) );
  INV_X1 S_5_F_Inst_0__CF_Inst_U1 ( .A(S_5_F_in1[3]), .ZN(
        S_5_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_5_F_Inst_1__CF_Inst_U2 ( .A(S_5_F_Inst_1__CF_Inst_n3), .B(
        S_5_F_in1[1]), .ZN(S_5_F_CF_Out[1]) );
  NAND2_X1 S_5_F_Inst_1__CF_Inst_U1 ( .A1(S_5_F_in2[2]), .A2(S_5_F_in1[3]), 
        .ZN(S_5_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_5_F_Inst_2__CF_Inst_U1 ( .A1(S_5_F_in1[3]), .A2(S_5_F_in3[2]), .ZN(
        S_5_F_CF_Out[2]) );
  NOR2_X1 S_5_F_Inst_3__CF_Inst_U2 ( .A1(S_5_F_in2[3]), .A2(
        S_5_F_Inst_3__CF_Inst_n3), .ZN(S_5_F_CF_Out[3]) );
  INV_X1 S_5_F_Inst_3__CF_Inst_U1 ( .A(S_5_F_in1[2]), .ZN(
        S_5_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_5_F_Inst_4__CF_Inst_U2 ( .A(S_5_F_Inst_4__CF_Inst_n3), .B(
        S_5_F_in2[1]), .ZN(S_5_F_CF_Out[4]) );
  NAND2_X1 S_5_F_Inst_4__CF_Inst_U1 ( .A1(S_5_F_in2[2]), .A2(S_5_F_in2[3]), 
        .ZN(S_5_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_5_F_Inst_5__CF_Inst_U1 ( .A1(S_5_F_in3[2]), .A2(S_5_F_in2[3]), 
        .ZN(S_5_F_CF_Out[5]) );
  XNOR2_X1 S_5_F_Inst_6__CF_Inst_U2 ( .A(S_5_F_Inst_6__CF_Inst_n7), .B(
        S_5_F_in3[1]), .ZN(S_5_F_CF_Out[6]) );
  NOR2_X1 S_5_F_Inst_6__CF_Inst_U1 ( .A1(S_5_F_in1[2]), .A2(S_5_F_in3[3]), 
        .ZN(S_5_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_5_F_Inst_7__CF_Inst_U1 ( .A1(S_5_F_in2[2]), .A2(S_5_F_in3[3]), 
        .ZN(S_5_F_CF_Out[7]) );
  OR2_X1 S_5_F_Inst_8__CF_Inst_U1 ( .A1(S_5_F_in3[3]), .A2(S_5_F_in3[2]), .ZN(
        S_5_F_CF_Out[8]) );
  NOR2_X1 S_5_F_Inst_9__CF_Inst_U2 ( .A1(S_5_F_in1[3]), .A2(
        S_5_F_Inst_9__CF_Inst_n3), .ZN(S_5_F_CF_Out[9]) );
  INV_X1 S_5_F_Inst_9__CF_Inst_U1 ( .A(S_5_F_in1[1]), .ZN(
        S_5_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_5_F_Inst_10__CF_Inst_U1 ( .A1(S_5_F_in2[1]), .A2(S_5_F_in1[3]), 
        .ZN(S_5_F_CF_Out[10]) );
  XNOR2_X1 S_5_F_Inst_11__CF_Inst_U2 ( .A(S_5_F_Inst_11__CF_Inst_n3), .B(
        S_5_F_in1[0]), .ZN(S_5_F_CF_Out[11]) );
  NAND2_X1 S_5_F_Inst_11__CF_Inst_U1 ( .A1(S_5_F_in3[1]), .A2(S_5_F_in1[3]), 
        .ZN(S_5_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_5_F_Inst_12__CF_Inst_U2 ( .A(S_5_F_Inst_12__CF_Inst_n3), .B(
        S_5_F_in2[0]), .ZN(S_5_F_CF_Out[12]) );
  NAND2_X1 S_5_F_Inst_12__CF_Inst_U1 ( .A1(S_5_F_in1[1]), .A2(S_5_F_in2[3]), 
        .ZN(S_5_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_5_F_Inst_13__CF_Inst_U2 ( .A1(S_5_F_in2[3]), .A2(
        S_5_F_Inst_13__CF_Inst_n3), .ZN(S_5_F_CF_Out[13]) );
  INV_X1 S_5_F_Inst_13__CF_Inst_U1 ( .A(S_5_F_in2[1]), .ZN(
        S_5_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_5_F_Inst_14__CF_Inst_U1 ( .A1(S_5_F_in3[1]), .A2(S_5_F_in2[3]), 
        .ZN(S_5_F_CF_Out[14]) );
  XNOR2_X1 S_5_F_Inst_15__CF_Inst_U2 ( .A(S_5_F_Inst_15__CF_Inst_n7), .B(
        S_5_F_in3[0]), .ZN(S_5_F_CF_Out[15]) );
  NOR2_X1 S_5_F_Inst_15__CF_Inst_U1 ( .A1(S_5_F_in1[1]), .A2(S_5_F_in3[3]), 
        .ZN(S_5_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_5_F_Inst_16__CF_Inst_U2 ( .A1(S_5_F_in3[3]), .A2(
        S_5_F_Inst_16__CF_Inst_n3), .ZN(S_5_F_CF_Out[16]) );
  INV_X1 S_5_F_Inst_16__CF_Inst_U1 ( .A(S_5_F_in2[1]), .ZN(
        S_5_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_5_F_Inst_17__CF_Inst_U2 ( .A1(S_5_F_in3[1]), .A2(
        S_5_F_Inst_17__CF_Inst_n3), .ZN(S_5_F_CF_Out[17]) );
  INV_X1 S_5_F_Inst_17__CF_Inst_U1 ( .A(S_5_F_in3[3]), .ZN(
        S_5_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_5_F_InstXOR_0__Compression1_U2 ( .A(
        S_5_F_InstXOR_0__Compression1_n3), .B(S_5_F_CF_Reg[2]), .ZN(
        S_5_F_q1[2]) );
  XNOR2_X1 S_5_F_InstXOR_0__Compression1_U1 ( .A(S_5_F_CF_Reg[0]), .B(
        S_5_F_CF_Reg[1]), .ZN(S_5_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_5_F_InstXOR_0__Compression2_U2 ( .A(
        S_5_F_InstXOR_0__Compression2_n3), .B(S_5_F_CF_Reg[5]), .ZN(
        S_5_F_q2[2]) );
  XNOR2_X1 S_5_F_InstXOR_0__Compression2_U1 ( .A(S_5_F_CF_Reg[3]), .B(
        S_5_F_CF_Reg[4]), .ZN(S_5_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_5_F_InstXOR_0__Compression3_U2 ( .A(
        S_5_F_InstXOR_0__Compression3_n3), .B(S_5_F_CF_Reg[8]), .ZN(
        S_5_F_q3[2]) );
  XNOR2_X1 S_5_F_InstXOR_0__Compression3_U1 ( .A(S_5_F_CF_Reg[6]), .B(
        S_5_F_CF_Reg[7]), .ZN(S_5_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_5_F_InstXOR_1__Compression1_U2 ( .A(
        S_5_F_InstXOR_1__Compression1_n3), .B(S_5_F_CF_Reg[11]), .ZN(
        S_5_F_q1[3]) );
  XNOR2_X1 S_5_F_InstXOR_1__Compression1_U1 ( .A(S_5_F_CF_Reg[9]), .B(
        S_5_F_CF_Reg[10]), .ZN(S_5_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_5_F_InstXOR_1__Compression2_U2 ( .A(
        S_5_F_InstXOR_1__Compression2_n3), .B(S_5_F_CF_Reg[14]), .ZN(
        S_5_F_q2[3]) );
  XNOR2_X1 S_5_F_InstXOR_1__Compression2_U1 ( .A(S_5_F_CF_Reg[12]), .B(
        S_5_F_CF_Reg[13]), .ZN(S_5_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_5_F_InstXOR_1__Compression3_U2 ( .A(
        S_5_F_InstXOR_1__Compression3_n3), .B(S_5_F_CF_Reg[17]), .ZN(
        S_5_F_q3[3]) );
  XNOR2_X1 S_5_F_InstXOR_1__Compression3_U1 ( .A(S_5_F_CF_Reg[15]), .B(
        S_5_F_CF_Reg[16]), .ZN(S_5_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_5_G_CF_Reg_reg_0_ ( .D(S_5_G_CF_Out[0]), .CK(CLK), .Q(
        S_5_G_CF_Reg[0]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_1_ ( .D(S_5_G_CF_Out[1]), .CK(CLK), .Q(
        S_5_G_CF_Reg[1]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_2_ ( .D(S_5_G_CF_Out[2]), .CK(CLK), .Q(
        S_5_G_CF_Reg[2]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_3_ ( .D(S_5_G_CF_Out[3]), .CK(CLK), .Q(
        S_5_G_CF_Reg[3]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_4_ ( .D(S_5_G_CF_Out[4]), .CK(CLK), .Q(
        S_5_G_CF_Reg[4]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_5_ ( .D(S_5_G_CF_Out[5]), .CK(CLK), .Q(
        S_5_G_CF_Reg[5]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_6_ ( .D(S_5_G_CF_Out[6]), .CK(CLK), .Q(
        S_5_G_CF_Reg[6]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_7_ ( .D(S_5_G_CF_Out[7]), .CK(CLK), .Q(
        S_5_G_CF_Reg[7]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_8_ ( .D(S_5_G_CF_Out[8]), .CK(CLK), .Q(
        S_5_G_CF_Reg[8]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_9_ ( .D(S_5_G_CF_Out[9]), .CK(CLK), .Q(
        S_5_G_CF_Reg[9]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_10_ ( .D(S_5_G_CF_Out[10]), .CK(CLK), .Q(
        S_5_G_CF_Reg[10]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_11_ ( .D(S_5_G_CF_Out[11]), .CK(CLK), .Q(
        S_5_G_CF_Reg[11]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_12_ ( .D(S_5_G_CF_Out[12]), .CK(CLK), .Q(
        S_5_G_CF_Reg[12]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_13_ ( .D(S_5_G_CF_Out[13]), .CK(CLK), .Q(
        S_5_G_CF_Reg[13]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_14_ ( .D(S_5_G_CF_Out[14]), .CK(CLK), .Q(
        S_5_G_CF_Reg[14]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_15_ ( .D(S_5_G_CF_Out[15]), .CK(CLK), .Q(
        S_5_G_CF_Reg[15]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_16_ ( .D(S_5_G_CF_Out[16]), .CK(CLK), .Q(
        S_5_G_CF_Reg[16]), .QN() );
  DFF_X1 S_5_G_CF_Reg_reg_17_ ( .D(S_5_G_CF_Out[17]), .CK(CLK), .Q(
        S_5_G_CF_Reg[17]), .QN() );
  DFF_X1 S_5_G_out1_reg_2_ ( .D(S_5_Rq1[2]), .CK(CLK), .Q(S_5_G_out1[2]), 
        .QN() );
  DFF_X1 S_5_G_out1_reg_3_ ( .D(S_5_Rq1[3]), .CK(CLK), .Q(S_5_G_out1[3]), 
        .QN() );
  DFF_X1 S_5_G_out2_reg_2_ ( .D(S_5_Rq2[2]), .CK(CLK), .Q(RF2_SHIFTROWS[30]), 
        .QN() );
  DFF_X1 S_5_G_out2_reg_3_ ( .D(S_5_Rq2[3]), .CK(CLK), .Q(RF2_SHIFTROWS[31]), 
        .QN() );
  DFF_X1 S_5_G_out3_reg_2_ ( .D(S_5_Rq3[2]), .CK(CLK), .Q(RF3_SHIFTROWS[30]), 
        .QN() );
  DFF_X1 S_5_G_out3_reg_3_ ( .D(S_5_Rq3[3]), .CK(CLK), .Q(RF3_SHIFTROWS[31]), 
        .QN() );
  AND2_X1 S_5_G_Inst_0__CF_Inst_U1 ( .A1(S_5_Rq1[1]), .A2(S_5_Rq1[3]), .ZN(
        S_5_G_CF_Out[0]) );
  NOR2_X1 S_5_G_Inst_1__CF_Inst_U2 ( .A1(S_5_Rq1[3]), .A2(
        S_5_G_Inst_1__CF_Inst_n3), .ZN(S_5_G_CF_Out[1]) );
  INV_X1 S_5_G_Inst_1__CF_Inst_U1 ( .A(S_5_Rq2[1]), .ZN(
        S_5_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_5_G_Inst_2__CF_Inst_U2 ( .A(S_5_G_Inst_2__CF_Inst_n3), .B(
        S_5_Rq2[0]), .ZN(S_5_G_CF_Out[2]) );
  NAND2_X1 S_5_G_Inst_2__CF_Inst_U1 ( .A1(S_5_Rq1[1]), .A2(S_5_Rq2[3]), .ZN(
        S_5_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_5_G_Inst_3__CF_Inst_U3 ( .A(S_5_Rq1[0]), .B(
        S_5_G_Inst_3__CF_Inst_n6), .ZN(S_5_G_CF_Out[3]) );
  NAND2_X1 S_5_G_Inst_3__CF_Inst_U2 ( .A1(S_5_Rq3[1]), .A2(
        S_5_G_Inst_3__CF_Inst_n5), .ZN(S_5_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_5_G_Inst_3__CF_Inst_U1 ( .A(S_5_Rq1[3]), .ZN(
        S_5_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_5_G_Inst_4__CF_Inst_U1 ( .A1(S_5_Rq2[1]), .A2(S_5_Rq2[3]), .ZN(
        S_5_G_CF_Out[4]) );
  OR2_X1 S_5_G_Inst_5__CF_Inst_U1 ( .A1(S_5_Rq3[3]), .A2(S_5_Rq2[1]), .ZN(
        S_5_G_CF_Out[5]) );
  AND2_X1 S_5_G_Inst_6__CF_Inst_U1 ( .A1(S_5_Rq3[1]), .A2(S_5_Rq2[3]), .ZN(
        S_5_G_CF_Out[6]) );
  XNOR2_X1 S_5_G_Inst_7__CF_Inst_U2 ( .A(S_5_G_Inst_7__CF_Inst_n3), .B(
        S_5_Rq3[0]), .ZN(S_5_G_CF_Out[7]) );
  NAND2_X1 S_5_G_Inst_7__CF_Inst_U1 ( .A1(S_5_Rq1[1]), .A2(S_5_Rq3[3]), .ZN(
        S_5_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_5_G_Inst_8__CF_Inst_U1 ( .A1(S_5_Rq3[3]), .A2(S_5_Rq3[1]), .ZN(
        S_5_G_CF_Out[8]) );
  NOR2_X1 S_5_G_Inst_9__CF_Inst_U2 ( .A1(S_5_Rq1[3]), .A2(
        S_5_G_Inst_9__CF_Inst_n3), .ZN(S_5_G_CF_Out[9]) );
  INV_X1 S_5_G_Inst_9__CF_Inst_U1 ( .A(S_5_Rq1[2]), .ZN(
        S_5_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_5_G_Inst_10__CF_Inst_U2 ( .A1(S_5_Rq2[2]), .A2(
        S_5_G_Inst_10__CF_Inst_n3), .ZN(S_5_G_CF_Out[10]) );
  INV_X1 S_5_G_Inst_10__CF_Inst_U1 ( .A(S_5_Rq1[3]), .ZN(
        S_5_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_5_G_Inst_11__CF_Inst_U3 ( .A(S_5_Rq1[1]), .B(
        S_5_G_Inst_11__CF_Inst_n6), .ZN(S_5_G_CF_Out[11]) );
  NAND2_X1 S_5_G_Inst_11__CF_Inst_U2 ( .A1(S_5_Rq1[3]), .A2(
        S_5_G_Inst_11__CF_Inst_n5), .ZN(S_5_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_5_G_Inst_11__CF_Inst_U1 ( .A(S_5_Rq3[2]), .ZN(
        S_5_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_5_G_Inst_12__CF_Inst_U2 ( .A1(S_5_Rq2[3]), .A2(
        S_5_G_Inst_12__CF_Inst_n3), .ZN(S_5_G_CF_Out[12]) );
  INV_X1 S_5_G_Inst_12__CF_Inst_U1 ( .A(S_5_Rq1[2]), .ZN(
        S_5_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_5_G_Inst_13__CF_Inst_U1 ( .A1(S_5_Rq2[2]), .A2(S_5_Rq2[3]), .ZN(
        S_5_G_CF_Out[13]) );
  XNOR2_X1 S_5_G_Inst_14__CF_Inst_U3 ( .A(S_5_Rq2[1]), .B(
        S_5_G_Inst_14__CF_Inst_n6), .ZN(S_5_G_CF_Out[14]) );
  NAND2_X1 S_5_G_Inst_14__CF_Inst_U2 ( .A1(S_5_Rq3[2]), .A2(
        S_5_G_Inst_14__CF_Inst_n5), .ZN(S_5_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_5_G_Inst_14__CF_Inst_U1 ( .A(S_5_Rq2[3]), .ZN(
        S_5_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_5_G_Inst_15__CF_Inst_U2 ( .A(S_5_G_Inst_15__CF_Inst_n3), .B(
        S_5_Rq3[1]), .ZN(S_5_G_CF_Out[15]) );
  NAND2_X1 S_5_G_Inst_15__CF_Inst_U1 ( .A1(S_5_Rq1[2]), .A2(S_5_Rq3[3]), .ZN(
        S_5_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_5_G_Inst_16__CF_Inst_U1 ( .A1(S_5_Rq2[2]), .A2(S_5_Rq3[3]), .ZN(
        S_5_G_CF_Out[16]) );
  NOR2_X1 S_5_G_Inst_17__CF_Inst_U2 ( .A1(S_5_Rq3[3]), .A2(
        S_5_G_Inst_17__CF_Inst_n3), .ZN(S_5_G_CF_Out[17]) );
  INV_X1 S_5_G_Inst_17__CF_Inst_U1 ( .A(S_5_Rq3[2]), .ZN(
        S_5_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_5_G_InstXOR_0__Compression1_U2 ( .A(
        S_5_G_InstXOR_0__Compression1_n3), .B(S_5_G_CF_Reg[2]), .ZN(
        S_5_G_out1[0]) );
  XNOR2_X1 S_5_G_InstXOR_0__Compression1_U1 ( .A(S_5_G_CF_Reg[0]), .B(
        S_5_G_CF_Reg[1]), .ZN(S_5_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_5_G_InstXOR_0__Compression2_U2 ( .A(
        S_5_G_InstXOR_0__Compression2_n3), .B(S_5_G_CF_Reg[5]), .ZN(
        RF2_SHIFTROWS[29]) );
  XNOR2_X1 S_5_G_InstXOR_0__Compression2_U1 ( .A(S_5_G_CF_Reg[3]), .B(
        S_5_G_CF_Reg[4]), .ZN(S_5_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_5_G_InstXOR_0__Compression3_U2 ( .A(
        S_5_G_InstXOR_0__Compression3_n3), .B(S_5_G_CF_Reg[8]), .ZN(
        RF3_SHIFTROWS[29]) );
  XNOR2_X1 S_5_G_InstXOR_0__Compression3_U1 ( .A(S_5_G_CF_Reg[6]), .B(
        S_5_G_CF_Reg[7]), .ZN(S_5_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_5_G_InstXOR_1__Compression1_U2 ( .A(
        S_5_G_InstXOR_1__Compression1_n3), .B(S_5_G_CF_Reg[11]), .ZN(
        S_5_G_out1[1]) );
  XNOR2_X1 S_5_G_InstXOR_1__Compression1_U1 ( .A(S_5_G_CF_Reg[9]), .B(
        S_5_G_CF_Reg[10]), .ZN(S_5_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_5_G_InstXOR_1__Compression2_U2 ( .A(
        S_5_G_InstXOR_1__Compression2_n3), .B(S_5_G_CF_Reg[14]), .ZN(
        RF2_SHIFTROWS[28]) );
  XNOR2_X1 S_5_G_InstXOR_1__Compression2_U1 ( .A(S_5_G_CF_Reg[12]), .B(
        S_5_G_CF_Reg[13]), .ZN(S_5_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_5_G_InstXOR_1__Compression3_U2 ( .A(
        S_5_G_InstXOR_1__Compression3_n3), .B(S_5_G_CF_Reg[17]), .ZN(
        RF3_SHIFTROWS[28]) );
  XNOR2_X1 S_5_G_InstXOR_1__Compression3_U1 ( .A(S_5_G_CF_Reg[15]), .B(
        S_5_G_CF_Reg[16]), .ZN(S_5_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_5_OutputAffine_U4 ( .A(S_5_G_out1[3]), .ZN(RF1_SHIFTROWS[31]) );
  INV_X1 S_5_OutputAffine_U3 ( .A(S_5_G_out1[2]), .ZN(RF1_SHIFTROWS[30]) );
  INV_X1 S_5_OutputAffine_U2 ( .A(S_5_G_out1[1]), .ZN(RF1_SHIFTROWS[28]) );
  INV_X1 S_5_OutputAffine_U1 ( .A(S_5_G_out1[0]), .ZN(RF1_SHIFTROWS[29]) );
  DFF_X1 S_6_Rq3_reg_0_ ( .D(S_6_q3[0]), .CK(CLK), .Q(S_6_Rq3[0]), .QN() );
  DFF_X1 S_6_Rq3_reg_1_ ( .D(S_6_q3[1]), .CK(CLK), .Q(S_6_Rq3[1]), .QN() );
  DFF_X1 S_6_Rq3_reg_2_ ( .D(S_6_q3[2]), .CK(CLK), .Q(S_6_Rq3[2]), .QN() );
  DFF_X1 S_6_Rq3_reg_3_ ( .D(S_6_q3[3]), .CK(CLK), .Q(S_6_Rq3[3]), .QN() );
  DFF_X1 S_6_Rq2_reg_0_ ( .D(S_6_q2[0]), .CK(CLK), .Q(S_6_Rq2[0]), .QN() );
  DFF_X1 S_6_Rq2_reg_1_ ( .D(S_6_q2[1]), .CK(CLK), .Q(S_6_Rq2[1]), .QN() );
  DFF_X1 S_6_Rq2_reg_2_ ( .D(S_6_q2[2]), .CK(CLK), .Q(S_6_Rq2[2]), .QN() );
  DFF_X1 S_6_Rq2_reg_3_ ( .D(S_6_q2[3]), .CK(CLK), .Q(S_6_Rq2[3]), .QN() );
  DFF_X1 S_6_Rq1_reg_0_ ( .D(S_6_q1[0]), .CK(CLK), .Q(S_6_Rq1[0]), .QN() );
  DFF_X1 S_6_Rq1_reg_1_ ( .D(S_6_q1[1]), .CK(CLK), .Q(S_6_Rq1[1]), .QN() );
  DFF_X1 S_6_Rq1_reg_2_ ( .D(S_6_q1[2]), .CK(CLK), .Q(S_6_Rq1[2]), .QN() );
  DFF_X1 S_6_Rq1_reg_3_ ( .D(S_6_q1[3]), .CK(CLK), .Q(S_6_Rq1[3]), .QN() );
  INV_X1 S_6_InputAffine_U4 ( .A(SUB_IN1[24]), .ZN(S_6_F_in1[0]) );
  INV_X1 S_6_InputAffine_U3 ( .A(SUB_IN1[26]), .ZN(S_6_F_in1[3]) );
  INV_X1 S_6_InputAffine_U2 ( .A(SUB_IN1[27]), .ZN(S_6_F_in1[1]) );
  INV_X1 S_6_InputAffine_U1 ( .A(SUB_IN1[25]), .ZN(S_6_F_in1[2]) );
  XNOR2_X1 S_6_F_U18 ( .A(S_6_F_n12), .B(FRESH[51]), .ZN(S_6_q3[3]) );
  XNOR2_X1 S_6_F_U17 ( .A(FRESH[50]), .B(S_6_F_q3[3]), .ZN(S_6_F_n12) );
  XNOR2_X1 S_6_F_U16 ( .A(S_6_F_n11), .B(FRESH[49]), .ZN(S_6_q3[2]) );
  XNOR2_X1 S_6_F_U15 ( .A(FRESH[48]), .B(S_6_F_q3[2]), .ZN(S_6_F_n11) );
  XOR2_X1 S_6_F_U14 ( .A(FRESH[51]), .B(S_6_F_q2[3]), .Z(S_6_q2[3]) );
  XOR2_X1 S_6_F_U13 ( .A(FRESH[49]), .B(S_6_F_q2[2]), .Z(S_6_q2[2]) );
  XOR2_X1 S_6_F_U12 ( .A(FRESH[50]), .B(S_6_F_q1[3]), .Z(S_6_q1[3]) );
  XOR2_X1 S_6_F_U11 ( .A(FRESH[48]), .B(S_6_F_q1[2]), .Z(S_6_q1[2]) );
  XNOR2_X1 S_6_F_U10 ( .A(S_6_F_n10), .B(FRESH[53]), .ZN(S_6_F_N5) );
  XNOR2_X1 S_6_F_U9 ( .A(S_6_F_in3[3]), .B(FRESH[52]), .ZN(S_6_F_n10) );
  XOR2_X1 S_6_F_U8 ( .A(FRESH[53]), .B(S_6_F_in2[3]), .Z(S_6_F_N4) );
  XOR2_X1 S_6_F_U7 ( .A(FRESH[52]), .B(S_6_F_in1[3]), .Z(S_6_F_N3) );
  XNOR2_X1 S_6_F_U6 ( .A(S_6_F_n9), .B(FRESH[55]), .ZN(S_6_F_N2) );
  XNOR2_X1 S_6_F_U5 ( .A(S_6_F_in3[2]), .B(FRESH[54]), .ZN(S_6_F_n9) );
  XOR2_X1 S_6_F_U4 ( .A(FRESH[55]), .B(S_6_F_in2[2]), .Z(S_6_F_N1) );
  XOR2_X1 S_6_F_U3 ( .A(FRESH[54]), .B(S_6_F_in1[2]), .Z(S_6_F_N0) );
  DFF_X1 S_6_F_CF_Reg_reg_0_ ( .D(S_6_F_CF_Out[0]), .CK(CLK), .Q(
        S_6_F_CF_Reg[0]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_1_ ( .D(S_6_F_CF_Out[1]), .CK(CLK), .Q(
        S_6_F_CF_Reg[1]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_2_ ( .D(S_6_F_CF_Out[2]), .CK(CLK), .Q(
        S_6_F_CF_Reg[2]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_3_ ( .D(S_6_F_CF_Out[3]), .CK(CLK), .Q(
        S_6_F_CF_Reg[3]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_4_ ( .D(S_6_F_CF_Out[4]), .CK(CLK), .Q(
        S_6_F_CF_Reg[4]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_5_ ( .D(S_6_F_CF_Out[5]), .CK(CLK), .Q(
        S_6_F_CF_Reg[5]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_6_ ( .D(S_6_F_CF_Out[6]), .CK(CLK), .Q(
        S_6_F_CF_Reg[6]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_7_ ( .D(S_6_F_CF_Out[7]), .CK(CLK), .Q(
        S_6_F_CF_Reg[7]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_8_ ( .D(S_6_F_CF_Out[8]), .CK(CLK), .Q(
        S_6_F_CF_Reg[8]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_9_ ( .D(S_6_F_CF_Out[9]), .CK(CLK), .Q(
        S_6_F_CF_Reg[9]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_10_ ( .D(S_6_F_CF_Out[10]), .CK(CLK), .Q(
        S_6_F_CF_Reg[10]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_11_ ( .D(S_6_F_CF_Out[11]), .CK(CLK), .Q(
        S_6_F_CF_Reg[11]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_12_ ( .D(S_6_F_CF_Out[12]), .CK(CLK), .Q(
        S_6_F_CF_Reg[12]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_13_ ( .D(S_6_F_CF_Out[13]), .CK(CLK), .Q(
        S_6_F_CF_Reg[13]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_14_ ( .D(S_6_F_CF_Out[14]), .CK(CLK), .Q(
        S_6_F_CF_Reg[14]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_15_ ( .D(S_6_F_CF_Out[15]), .CK(CLK), .Q(
        S_6_F_CF_Reg[15]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_16_ ( .D(S_6_F_CF_Out[16]), .CK(CLK), .Q(
        S_6_F_CF_Reg[16]), .QN() );
  DFF_X1 S_6_F_CF_Reg_reg_17_ ( .D(S_6_F_CF_Out[17]), .CK(CLK), .Q(
        S_6_F_CF_Reg[17]), .QN() );
  DFF_X1 S_6_F_out2_reg_0_ ( .D(S_6_F_N4), .CK(CLK), .Q(S_6_q2[0]), .QN() );
  DFF_X1 S_6_F_out2_reg_1_ ( .D(S_6_F_N1), .CK(CLK), .Q(S_6_q2[1]), .QN() );
  DFF_X1 S_6_F_out3_reg_0_ ( .D(S_6_F_N5), .CK(CLK), .Q(S_6_q3[0]), .QN() );
  DFF_X1 S_6_F_out3_reg_1_ ( .D(S_6_F_N2), .CK(CLK), .Q(S_6_q3[1]), .QN() );
  DFF_X1 S_6_F_out1_reg_0_ ( .D(S_6_F_N3), .CK(CLK), .Q(S_6_q1[0]), .QN() );
  DFF_X1 S_6_F_out1_reg_1_ ( .D(S_6_F_N0), .CK(CLK), .Q(S_6_q1[1]), .QN() );
  NOR2_X1 S_6_F_Inst_0__CF_Inst_U2 ( .A1(S_6_F_in1[2]), .A2(
        S_6_F_Inst_0__CF_Inst_n3), .ZN(S_6_F_CF_Out[0]) );
  INV_X1 S_6_F_Inst_0__CF_Inst_U1 ( .A(S_6_F_in1[3]), .ZN(
        S_6_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_6_F_Inst_1__CF_Inst_U2 ( .A(S_6_F_Inst_1__CF_Inst_n3), .B(
        S_6_F_in1[1]), .ZN(S_6_F_CF_Out[1]) );
  NAND2_X1 S_6_F_Inst_1__CF_Inst_U1 ( .A1(S_6_F_in2[2]), .A2(S_6_F_in1[3]), 
        .ZN(S_6_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_6_F_Inst_2__CF_Inst_U1 ( .A1(S_6_F_in1[3]), .A2(S_6_F_in3[2]), .ZN(
        S_6_F_CF_Out[2]) );
  NOR2_X1 S_6_F_Inst_3__CF_Inst_U2 ( .A1(S_6_F_in2[3]), .A2(
        S_6_F_Inst_3__CF_Inst_n3), .ZN(S_6_F_CF_Out[3]) );
  INV_X1 S_6_F_Inst_3__CF_Inst_U1 ( .A(S_6_F_in1[2]), .ZN(
        S_6_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_6_F_Inst_4__CF_Inst_U2 ( .A(S_6_F_Inst_4__CF_Inst_n3), .B(
        S_6_F_in2[1]), .ZN(S_6_F_CF_Out[4]) );
  NAND2_X1 S_6_F_Inst_4__CF_Inst_U1 ( .A1(S_6_F_in2[2]), .A2(S_6_F_in2[3]), 
        .ZN(S_6_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_6_F_Inst_5__CF_Inst_U1 ( .A1(S_6_F_in3[2]), .A2(S_6_F_in2[3]), 
        .ZN(S_6_F_CF_Out[5]) );
  XNOR2_X1 S_6_F_Inst_6__CF_Inst_U2 ( .A(S_6_F_Inst_6__CF_Inst_n7), .B(
        S_6_F_in3[1]), .ZN(S_6_F_CF_Out[6]) );
  NOR2_X1 S_6_F_Inst_6__CF_Inst_U1 ( .A1(S_6_F_in1[2]), .A2(S_6_F_in3[3]), 
        .ZN(S_6_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_6_F_Inst_7__CF_Inst_U1 ( .A1(S_6_F_in2[2]), .A2(S_6_F_in3[3]), 
        .ZN(S_6_F_CF_Out[7]) );
  OR2_X1 S_6_F_Inst_8__CF_Inst_U1 ( .A1(S_6_F_in3[3]), .A2(S_6_F_in3[2]), .ZN(
        S_6_F_CF_Out[8]) );
  NOR2_X1 S_6_F_Inst_9__CF_Inst_U2 ( .A1(S_6_F_in1[3]), .A2(
        S_6_F_Inst_9__CF_Inst_n3), .ZN(S_6_F_CF_Out[9]) );
  INV_X1 S_6_F_Inst_9__CF_Inst_U1 ( .A(S_6_F_in1[1]), .ZN(
        S_6_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_6_F_Inst_10__CF_Inst_U1 ( .A1(S_6_F_in2[1]), .A2(S_6_F_in1[3]), 
        .ZN(S_6_F_CF_Out[10]) );
  XNOR2_X1 S_6_F_Inst_11__CF_Inst_U2 ( .A(S_6_F_Inst_11__CF_Inst_n3), .B(
        S_6_F_in1[0]), .ZN(S_6_F_CF_Out[11]) );
  NAND2_X1 S_6_F_Inst_11__CF_Inst_U1 ( .A1(S_6_F_in3[1]), .A2(S_6_F_in1[3]), 
        .ZN(S_6_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_6_F_Inst_12__CF_Inst_U2 ( .A(S_6_F_Inst_12__CF_Inst_n3), .B(
        S_6_F_in2[0]), .ZN(S_6_F_CF_Out[12]) );
  NAND2_X1 S_6_F_Inst_12__CF_Inst_U1 ( .A1(S_6_F_in1[1]), .A2(S_6_F_in2[3]), 
        .ZN(S_6_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_6_F_Inst_13__CF_Inst_U2 ( .A1(S_6_F_in2[3]), .A2(
        S_6_F_Inst_13__CF_Inst_n3), .ZN(S_6_F_CF_Out[13]) );
  INV_X1 S_6_F_Inst_13__CF_Inst_U1 ( .A(S_6_F_in2[1]), .ZN(
        S_6_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_6_F_Inst_14__CF_Inst_U1 ( .A1(S_6_F_in3[1]), .A2(S_6_F_in2[3]), 
        .ZN(S_6_F_CF_Out[14]) );
  XNOR2_X1 S_6_F_Inst_15__CF_Inst_U2 ( .A(S_6_F_Inst_15__CF_Inst_n7), .B(
        S_6_F_in3[0]), .ZN(S_6_F_CF_Out[15]) );
  NOR2_X1 S_6_F_Inst_15__CF_Inst_U1 ( .A1(S_6_F_in1[1]), .A2(S_6_F_in3[3]), 
        .ZN(S_6_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_6_F_Inst_16__CF_Inst_U2 ( .A1(S_6_F_in3[3]), .A2(
        S_6_F_Inst_16__CF_Inst_n3), .ZN(S_6_F_CF_Out[16]) );
  INV_X1 S_6_F_Inst_16__CF_Inst_U1 ( .A(S_6_F_in2[1]), .ZN(
        S_6_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_6_F_Inst_17__CF_Inst_U2 ( .A1(S_6_F_in3[1]), .A2(
        S_6_F_Inst_17__CF_Inst_n3), .ZN(S_6_F_CF_Out[17]) );
  INV_X1 S_6_F_Inst_17__CF_Inst_U1 ( .A(S_6_F_in3[3]), .ZN(
        S_6_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_6_F_InstXOR_0__Compression1_U2 ( .A(
        S_6_F_InstXOR_0__Compression1_n3), .B(S_6_F_CF_Reg[2]), .ZN(
        S_6_F_q1[2]) );
  XNOR2_X1 S_6_F_InstXOR_0__Compression1_U1 ( .A(S_6_F_CF_Reg[0]), .B(
        S_6_F_CF_Reg[1]), .ZN(S_6_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_6_F_InstXOR_0__Compression2_U2 ( .A(
        S_6_F_InstXOR_0__Compression2_n3), .B(S_6_F_CF_Reg[5]), .ZN(
        S_6_F_q2[2]) );
  XNOR2_X1 S_6_F_InstXOR_0__Compression2_U1 ( .A(S_6_F_CF_Reg[3]), .B(
        S_6_F_CF_Reg[4]), .ZN(S_6_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_6_F_InstXOR_0__Compression3_U2 ( .A(
        S_6_F_InstXOR_0__Compression3_n3), .B(S_6_F_CF_Reg[8]), .ZN(
        S_6_F_q3[2]) );
  XNOR2_X1 S_6_F_InstXOR_0__Compression3_U1 ( .A(S_6_F_CF_Reg[6]), .B(
        S_6_F_CF_Reg[7]), .ZN(S_6_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_6_F_InstXOR_1__Compression1_U2 ( .A(
        S_6_F_InstXOR_1__Compression1_n3), .B(S_6_F_CF_Reg[11]), .ZN(
        S_6_F_q1[3]) );
  XNOR2_X1 S_6_F_InstXOR_1__Compression1_U1 ( .A(S_6_F_CF_Reg[9]), .B(
        S_6_F_CF_Reg[10]), .ZN(S_6_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_6_F_InstXOR_1__Compression2_U2 ( .A(
        S_6_F_InstXOR_1__Compression2_n3), .B(S_6_F_CF_Reg[14]), .ZN(
        S_6_F_q2[3]) );
  XNOR2_X1 S_6_F_InstXOR_1__Compression2_U1 ( .A(S_6_F_CF_Reg[12]), .B(
        S_6_F_CF_Reg[13]), .ZN(S_6_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_6_F_InstXOR_1__Compression3_U2 ( .A(
        S_6_F_InstXOR_1__Compression3_n3), .B(S_6_F_CF_Reg[17]), .ZN(
        S_6_F_q3[3]) );
  XNOR2_X1 S_6_F_InstXOR_1__Compression3_U1 ( .A(S_6_F_CF_Reg[15]), .B(
        S_6_F_CF_Reg[16]), .ZN(S_6_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_6_G_CF_Reg_reg_0_ ( .D(S_6_G_CF_Out[0]), .CK(CLK), .Q(
        S_6_G_CF_Reg[0]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_1_ ( .D(S_6_G_CF_Out[1]), .CK(CLK), .Q(
        S_6_G_CF_Reg[1]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_2_ ( .D(S_6_G_CF_Out[2]), .CK(CLK), .Q(
        S_6_G_CF_Reg[2]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_3_ ( .D(S_6_G_CF_Out[3]), .CK(CLK), .Q(
        S_6_G_CF_Reg[3]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_4_ ( .D(S_6_G_CF_Out[4]), .CK(CLK), .Q(
        S_6_G_CF_Reg[4]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_5_ ( .D(S_6_G_CF_Out[5]), .CK(CLK), .Q(
        S_6_G_CF_Reg[5]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_6_ ( .D(S_6_G_CF_Out[6]), .CK(CLK), .Q(
        S_6_G_CF_Reg[6]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_7_ ( .D(S_6_G_CF_Out[7]), .CK(CLK), .Q(
        S_6_G_CF_Reg[7]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_8_ ( .D(S_6_G_CF_Out[8]), .CK(CLK), .Q(
        S_6_G_CF_Reg[8]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_9_ ( .D(S_6_G_CF_Out[9]), .CK(CLK), .Q(
        S_6_G_CF_Reg[9]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_10_ ( .D(S_6_G_CF_Out[10]), .CK(CLK), .Q(
        S_6_G_CF_Reg[10]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_11_ ( .D(S_6_G_CF_Out[11]), .CK(CLK), .Q(
        S_6_G_CF_Reg[11]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_12_ ( .D(S_6_G_CF_Out[12]), .CK(CLK), .Q(
        S_6_G_CF_Reg[12]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_13_ ( .D(S_6_G_CF_Out[13]), .CK(CLK), .Q(
        S_6_G_CF_Reg[13]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_14_ ( .D(S_6_G_CF_Out[14]), .CK(CLK), .Q(
        S_6_G_CF_Reg[14]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_15_ ( .D(S_6_G_CF_Out[15]), .CK(CLK), .Q(
        S_6_G_CF_Reg[15]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_16_ ( .D(S_6_G_CF_Out[16]), .CK(CLK), .Q(
        S_6_G_CF_Reg[16]), .QN() );
  DFF_X1 S_6_G_CF_Reg_reg_17_ ( .D(S_6_G_CF_Out[17]), .CK(CLK), .Q(
        S_6_G_CF_Reg[17]), .QN() );
  DFF_X1 S_6_G_out1_reg_2_ ( .D(S_6_Rq1[2]), .CK(CLK), .Q(S_6_G_out1[2]), 
        .QN() );
  DFF_X1 S_6_G_out1_reg_3_ ( .D(S_6_Rq1[3]), .CK(CLK), .Q(S_6_G_out1[3]), 
        .QN() );
  DFF_X1 S_6_G_out2_reg_2_ ( .D(S_6_Rq2[2]), .CK(CLK), .Q(RF2_SHIFTROWS[18]), 
        .QN() );
  DFF_X1 S_6_G_out2_reg_3_ ( .D(S_6_Rq2[3]), .CK(CLK), .Q(RF2_SHIFTROWS[19]), 
        .QN() );
  DFF_X1 S_6_G_out3_reg_2_ ( .D(S_6_Rq3[2]), .CK(CLK), .Q(RF3_SHIFTROWS[18]), 
        .QN() );
  DFF_X1 S_6_G_out3_reg_3_ ( .D(S_6_Rq3[3]), .CK(CLK), .Q(RF3_SHIFTROWS[19]), 
        .QN() );
  AND2_X1 S_6_G_Inst_0__CF_Inst_U1 ( .A1(S_6_Rq1[1]), .A2(S_6_Rq1[3]), .ZN(
        S_6_G_CF_Out[0]) );
  NOR2_X1 S_6_G_Inst_1__CF_Inst_U2 ( .A1(S_6_Rq1[3]), .A2(
        S_6_G_Inst_1__CF_Inst_n3), .ZN(S_6_G_CF_Out[1]) );
  INV_X1 S_6_G_Inst_1__CF_Inst_U1 ( .A(S_6_Rq2[1]), .ZN(
        S_6_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_6_G_Inst_2__CF_Inst_U2 ( .A(S_6_G_Inst_2__CF_Inst_n3), .B(
        S_6_Rq2[0]), .ZN(S_6_G_CF_Out[2]) );
  NAND2_X1 S_6_G_Inst_2__CF_Inst_U1 ( .A1(S_6_Rq1[1]), .A2(S_6_Rq2[3]), .ZN(
        S_6_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_6_G_Inst_3__CF_Inst_U3 ( .A(S_6_Rq1[0]), .B(
        S_6_G_Inst_3__CF_Inst_n6), .ZN(S_6_G_CF_Out[3]) );
  NAND2_X1 S_6_G_Inst_3__CF_Inst_U2 ( .A1(S_6_Rq3[1]), .A2(
        S_6_G_Inst_3__CF_Inst_n5), .ZN(S_6_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_6_G_Inst_3__CF_Inst_U1 ( .A(S_6_Rq1[3]), .ZN(
        S_6_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_6_G_Inst_4__CF_Inst_U1 ( .A1(S_6_Rq2[1]), .A2(S_6_Rq2[3]), .ZN(
        S_6_G_CF_Out[4]) );
  OR2_X1 S_6_G_Inst_5__CF_Inst_U1 ( .A1(S_6_Rq3[3]), .A2(S_6_Rq2[1]), .ZN(
        S_6_G_CF_Out[5]) );
  AND2_X1 S_6_G_Inst_6__CF_Inst_U1 ( .A1(S_6_Rq3[1]), .A2(S_6_Rq2[3]), .ZN(
        S_6_G_CF_Out[6]) );
  XNOR2_X1 S_6_G_Inst_7__CF_Inst_U2 ( .A(S_6_G_Inst_7__CF_Inst_n3), .B(
        S_6_Rq3[0]), .ZN(S_6_G_CF_Out[7]) );
  NAND2_X1 S_6_G_Inst_7__CF_Inst_U1 ( .A1(S_6_Rq1[1]), .A2(S_6_Rq3[3]), .ZN(
        S_6_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_6_G_Inst_8__CF_Inst_U1 ( .A1(S_6_Rq3[3]), .A2(S_6_Rq3[1]), .ZN(
        S_6_G_CF_Out[8]) );
  NOR2_X1 S_6_G_Inst_9__CF_Inst_U2 ( .A1(S_6_Rq1[3]), .A2(
        S_6_G_Inst_9__CF_Inst_n3), .ZN(S_6_G_CF_Out[9]) );
  INV_X1 S_6_G_Inst_9__CF_Inst_U1 ( .A(S_6_Rq1[2]), .ZN(
        S_6_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_6_G_Inst_10__CF_Inst_U2 ( .A1(S_6_Rq2[2]), .A2(
        S_6_G_Inst_10__CF_Inst_n3), .ZN(S_6_G_CF_Out[10]) );
  INV_X1 S_6_G_Inst_10__CF_Inst_U1 ( .A(S_6_Rq1[3]), .ZN(
        S_6_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_6_G_Inst_11__CF_Inst_U3 ( .A(S_6_Rq1[1]), .B(
        S_6_G_Inst_11__CF_Inst_n6), .ZN(S_6_G_CF_Out[11]) );
  NAND2_X1 S_6_G_Inst_11__CF_Inst_U2 ( .A1(S_6_Rq1[3]), .A2(
        S_6_G_Inst_11__CF_Inst_n5), .ZN(S_6_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_6_G_Inst_11__CF_Inst_U1 ( .A(S_6_Rq3[2]), .ZN(
        S_6_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_6_G_Inst_12__CF_Inst_U2 ( .A1(S_6_Rq2[3]), .A2(
        S_6_G_Inst_12__CF_Inst_n3), .ZN(S_6_G_CF_Out[12]) );
  INV_X1 S_6_G_Inst_12__CF_Inst_U1 ( .A(S_6_Rq1[2]), .ZN(
        S_6_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_6_G_Inst_13__CF_Inst_U1 ( .A1(S_6_Rq2[2]), .A2(S_6_Rq2[3]), .ZN(
        S_6_G_CF_Out[13]) );
  XNOR2_X1 S_6_G_Inst_14__CF_Inst_U3 ( .A(S_6_Rq2[1]), .B(
        S_6_G_Inst_14__CF_Inst_n6), .ZN(S_6_G_CF_Out[14]) );
  NAND2_X1 S_6_G_Inst_14__CF_Inst_U2 ( .A1(S_6_Rq3[2]), .A2(
        S_6_G_Inst_14__CF_Inst_n5), .ZN(S_6_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_6_G_Inst_14__CF_Inst_U1 ( .A(S_6_Rq2[3]), .ZN(
        S_6_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_6_G_Inst_15__CF_Inst_U2 ( .A(S_6_G_Inst_15__CF_Inst_n3), .B(
        S_6_Rq3[1]), .ZN(S_6_G_CF_Out[15]) );
  NAND2_X1 S_6_G_Inst_15__CF_Inst_U1 ( .A1(S_6_Rq1[2]), .A2(S_6_Rq3[3]), .ZN(
        S_6_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_6_G_Inst_16__CF_Inst_U1 ( .A1(S_6_Rq2[2]), .A2(S_6_Rq3[3]), .ZN(
        S_6_G_CF_Out[16]) );
  NOR2_X1 S_6_G_Inst_17__CF_Inst_U2 ( .A1(S_6_Rq3[3]), .A2(
        S_6_G_Inst_17__CF_Inst_n3), .ZN(S_6_G_CF_Out[17]) );
  INV_X1 S_6_G_Inst_17__CF_Inst_U1 ( .A(S_6_Rq3[2]), .ZN(
        S_6_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_6_G_InstXOR_0__Compression1_U2 ( .A(
        S_6_G_InstXOR_0__Compression1_n3), .B(S_6_G_CF_Reg[2]), .ZN(
        S_6_G_out1[0]) );
  XNOR2_X1 S_6_G_InstXOR_0__Compression1_U1 ( .A(S_6_G_CF_Reg[0]), .B(
        S_6_G_CF_Reg[1]), .ZN(S_6_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_6_G_InstXOR_0__Compression2_U2 ( .A(
        S_6_G_InstXOR_0__Compression2_n3), .B(S_6_G_CF_Reg[5]), .ZN(
        RF2_SHIFTROWS[17]) );
  XNOR2_X1 S_6_G_InstXOR_0__Compression2_U1 ( .A(S_6_G_CF_Reg[3]), .B(
        S_6_G_CF_Reg[4]), .ZN(S_6_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_6_G_InstXOR_0__Compression3_U2 ( .A(
        S_6_G_InstXOR_0__Compression3_n3), .B(S_6_G_CF_Reg[8]), .ZN(
        RF3_SHIFTROWS[17]) );
  XNOR2_X1 S_6_G_InstXOR_0__Compression3_U1 ( .A(S_6_G_CF_Reg[6]), .B(
        S_6_G_CF_Reg[7]), .ZN(S_6_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_6_G_InstXOR_1__Compression1_U2 ( .A(
        S_6_G_InstXOR_1__Compression1_n3), .B(S_6_G_CF_Reg[11]), .ZN(
        S_6_G_out1[1]) );
  XNOR2_X1 S_6_G_InstXOR_1__Compression1_U1 ( .A(S_6_G_CF_Reg[9]), .B(
        S_6_G_CF_Reg[10]), .ZN(S_6_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_6_G_InstXOR_1__Compression2_U2 ( .A(
        S_6_G_InstXOR_1__Compression2_n3), .B(S_6_G_CF_Reg[14]), .ZN(
        RF2_SHIFTROWS[16]) );
  XNOR2_X1 S_6_G_InstXOR_1__Compression2_U1 ( .A(S_6_G_CF_Reg[12]), .B(
        S_6_G_CF_Reg[13]), .ZN(S_6_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_6_G_InstXOR_1__Compression3_U2 ( .A(
        S_6_G_InstXOR_1__Compression3_n3), .B(S_6_G_CF_Reg[17]), .ZN(
        RF3_SHIFTROWS[16]) );
  XNOR2_X1 S_6_G_InstXOR_1__Compression3_U1 ( .A(S_6_G_CF_Reg[15]), .B(
        S_6_G_CF_Reg[16]), .ZN(S_6_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_6_OutputAffine_U4 ( .A(S_6_G_out1[3]), .ZN(RF1_SHIFTROWS[19]) );
  INV_X1 S_6_OutputAffine_U3 ( .A(S_6_G_out1[2]), .ZN(RF1_SHIFTROWS[18]) );
  INV_X1 S_6_OutputAffine_U2 ( .A(S_6_G_out1[1]), .ZN(RF1_SHIFTROWS[16]) );
  INV_X1 S_6_OutputAffine_U1 ( .A(S_6_G_out1[0]), .ZN(RF1_SHIFTROWS[17]) );
  DFF_X1 S_7_Rq3_reg_0_ ( .D(S_7_q3[0]), .CK(CLK), .Q(S_7_Rq3[0]), .QN() );
  DFF_X1 S_7_Rq3_reg_1_ ( .D(S_7_q3[1]), .CK(CLK), .Q(S_7_Rq3[1]), .QN() );
  DFF_X1 S_7_Rq3_reg_2_ ( .D(S_7_q3[2]), .CK(CLK), .Q(S_7_Rq3[2]), .QN() );
  DFF_X1 S_7_Rq3_reg_3_ ( .D(S_7_q3[3]), .CK(CLK), .Q(S_7_Rq3[3]), .QN() );
  DFF_X1 S_7_Rq2_reg_0_ ( .D(S_7_q2[0]), .CK(CLK), .Q(S_7_Rq2[0]), .QN() );
  DFF_X1 S_7_Rq2_reg_1_ ( .D(S_7_q2[1]), .CK(CLK), .Q(S_7_Rq2[1]), .QN() );
  DFF_X1 S_7_Rq2_reg_2_ ( .D(S_7_q2[2]), .CK(CLK), .Q(S_7_Rq2[2]), .QN() );
  DFF_X1 S_7_Rq2_reg_3_ ( .D(S_7_q2[3]), .CK(CLK), .Q(S_7_Rq2[3]), .QN() );
  DFF_X1 S_7_Rq1_reg_0_ ( .D(S_7_q1[0]), .CK(CLK), .Q(S_7_Rq1[0]), .QN() );
  DFF_X1 S_7_Rq1_reg_1_ ( .D(S_7_q1[1]), .CK(CLK), .Q(S_7_Rq1[1]), .QN() );
  DFF_X1 S_7_Rq1_reg_2_ ( .D(S_7_q1[2]), .CK(CLK), .Q(S_7_Rq1[2]), .QN() );
  DFF_X1 S_7_Rq1_reg_3_ ( .D(S_7_q1[3]), .CK(CLK), .Q(S_7_Rq1[3]), .QN() );
  INV_X1 S_7_InputAffine_U4 ( .A(SUB_IN1[28]), .ZN(S_7_F_in1[0]) );
  INV_X1 S_7_InputAffine_U3 ( .A(SUB_IN1[30]), .ZN(S_7_F_in1[3]) );
  INV_X1 S_7_InputAffine_U2 ( .A(SUB_IN1[31]), .ZN(S_7_F_in1[1]) );
  INV_X1 S_7_InputAffine_U1 ( .A(SUB_IN1[29]), .ZN(S_7_F_in1[2]) );
  XNOR2_X1 S_7_F_U18 ( .A(S_7_F_n12), .B(FRESH[59]), .ZN(S_7_q3[3]) );
  XNOR2_X1 S_7_F_U17 ( .A(FRESH[58]), .B(S_7_F_q3[3]), .ZN(S_7_F_n12) );
  XNOR2_X1 S_7_F_U16 ( .A(S_7_F_n11), .B(FRESH[57]), .ZN(S_7_q3[2]) );
  XNOR2_X1 S_7_F_U15 ( .A(FRESH[56]), .B(S_7_F_q3[2]), .ZN(S_7_F_n11) );
  XOR2_X1 S_7_F_U14 ( .A(FRESH[59]), .B(S_7_F_q2[3]), .Z(S_7_q2[3]) );
  XOR2_X1 S_7_F_U13 ( .A(FRESH[57]), .B(S_7_F_q2[2]), .Z(S_7_q2[2]) );
  XOR2_X1 S_7_F_U12 ( .A(FRESH[58]), .B(S_7_F_q1[3]), .Z(S_7_q1[3]) );
  XOR2_X1 S_7_F_U11 ( .A(FRESH[56]), .B(S_7_F_q1[2]), .Z(S_7_q1[2]) );
  XNOR2_X1 S_7_F_U10 ( .A(S_7_F_n10), .B(FRESH[61]), .ZN(S_7_F_N5) );
  XNOR2_X1 S_7_F_U9 ( .A(S_7_F_in3[3]), .B(FRESH[60]), .ZN(S_7_F_n10) );
  XOR2_X1 S_7_F_U8 ( .A(FRESH[61]), .B(S_7_F_in2[3]), .Z(S_7_F_N4) );
  XOR2_X1 S_7_F_U7 ( .A(FRESH[60]), .B(S_7_F_in1[3]), .Z(S_7_F_N3) );
  XNOR2_X1 S_7_F_U6 ( .A(S_7_F_n9), .B(FRESH[63]), .ZN(S_7_F_N2) );
  XNOR2_X1 S_7_F_U5 ( .A(S_7_F_in3[2]), .B(FRESH[62]), .ZN(S_7_F_n9) );
  XOR2_X1 S_7_F_U4 ( .A(FRESH[63]), .B(S_7_F_in2[2]), .Z(S_7_F_N1) );
  XOR2_X1 S_7_F_U3 ( .A(FRESH[62]), .B(S_7_F_in1[2]), .Z(S_7_F_N0) );
  DFF_X1 S_7_F_CF_Reg_reg_0_ ( .D(S_7_F_CF_Out[0]), .CK(CLK), .Q(
        S_7_F_CF_Reg[0]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_1_ ( .D(S_7_F_CF_Out[1]), .CK(CLK), .Q(
        S_7_F_CF_Reg[1]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_2_ ( .D(S_7_F_CF_Out[2]), .CK(CLK), .Q(
        S_7_F_CF_Reg[2]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_3_ ( .D(S_7_F_CF_Out[3]), .CK(CLK), .Q(
        S_7_F_CF_Reg[3]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_4_ ( .D(S_7_F_CF_Out[4]), .CK(CLK), .Q(
        S_7_F_CF_Reg[4]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_5_ ( .D(S_7_F_CF_Out[5]), .CK(CLK), .Q(
        S_7_F_CF_Reg[5]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_6_ ( .D(S_7_F_CF_Out[6]), .CK(CLK), .Q(
        S_7_F_CF_Reg[6]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_7_ ( .D(S_7_F_CF_Out[7]), .CK(CLK), .Q(
        S_7_F_CF_Reg[7]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_8_ ( .D(S_7_F_CF_Out[8]), .CK(CLK), .Q(
        S_7_F_CF_Reg[8]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_9_ ( .D(S_7_F_CF_Out[9]), .CK(CLK), .Q(
        S_7_F_CF_Reg[9]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_10_ ( .D(S_7_F_CF_Out[10]), .CK(CLK), .Q(
        S_7_F_CF_Reg[10]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_11_ ( .D(S_7_F_CF_Out[11]), .CK(CLK), .Q(
        S_7_F_CF_Reg[11]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_12_ ( .D(S_7_F_CF_Out[12]), .CK(CLK), .Q(
        S_7_F_CF_Reg[12]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_13_ ( .D(S_7_F_CF_Out[13]), .CK(CLK), .Q(
        S_7_F_CF_Reg[13]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_14_ ( .D(S_7_F_CF_Out[14]), .CK(CLK), .Q(
        S_7_F_CF_Reg[14]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_15_ ( .D(S_7_F_CF_Out[15]), .CK(CLK), .Q(
        S_7_F_CF_Reg[15]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_16_ ( .D(S_7_F_CF_Out[16]), .CK(CLK), .Q(
        S_7_F_CF_Reg[16]), .QN() );
  DFF_X1 S_7_F_CF_Reg_reg_17_ ( .D(S_7_F_CF_Out[17]), .CK(CLK), .Q(
        S_7_F_CF_Reg[17]), .QN() );
  DFF_X1 S_7_F_out2_reg_0_ ( .D(S_7_F_N4), .CK(CLK), .Q(S_7_q2[0]), .QN() );
  DFF_X1 S_7_F_out2_reg_1_ ( .D(S_7_F_N1), .CK(CLK), .Q(S_7_q2[1]), .QN() );
  DFF_X1 S_7_F_out3_reg_0_ ( .D(S_7_F_N5), .CK(CLK), .Q(S_7_q3[0]), .QN() );
  DFF_X1 S_7_F_out3_reg_1_ ( .D(S_7_F_N2), .CK(CLK), .Q(S_7_q3[1]), .QN() );
  DFF_X1 S_7_F_out1_reg_0_ ( .D(S_7_F_N3), .CK(CLK), .Q(S_7_q1[0]), .QN() );
  DFF_X1 S_7_F_out1_reg_1_ ( .D(S_7_F_N0), .CK(CLK), .Q(S_7_q1[1]), .QN() );
  NOR2_X1 S_7_F_Inst_0__CF_Inst_U2 ( .A1(S_7_F_in1[2]), .A2(
        S_7_F_Inst_0__CF_Inst_n3), .ZN(S_7_F_CF_Out[0]) );
  INV_X1 S_7_F_Inst_0__CF_Inst_U1 ( .A(S_7_F_in1[3]), .ZN(
        S_7_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_7_F_Inst_1__CF_Inst_U2 ( .A(S_7_F_Inst_1__CF_Inst_n3), .B(
        S_7_F_in1[1]), .ZN(S_7_F_CF_Out[1]) );
  NAND2_X1 S_7_F_Inst_1__CF_Inst_U1 ( .A1(S_7_F_in2[2]), .A2(S_7_F_in1[3]), 
        .ZN(S_7_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_7_F_Inst_2__CF_Inst_U1 ( .A1(S_7_F_in1[3]), .A2(S_7_F_in3[2]), .ZN(
        S_7_F_CF_Out[2]) );
  NOR2_X1 S_7_F_Inst_3__CF_Inst_U2 ( .A1(S_7_F_in2[3]), .A2(
        S_7_F_Inst_3__CF_Inst_n3), .ZN(S_7_F_CF_Out[3]) );
  INV_X1 S_7_F_Inst_3__CF_Inst_U1 ( .A(S_7_F_in1[2]), .ZN(
        S_7_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_7_F_Inst_4__CF_Inst_U2 ( .A(S_7_F_Inst_4__CF_Inst_n3), .B(
        S_7_F_in2[1]), .ZN(S_7_F_CF_Out[4]) );
  NAND2_X1 S_7_F_Inst_4__CF_Inst_U1 ( .A1(S_7_F_in2[2]), .A2(S_7_F_in2[3]), 
        .ZN(S_7_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_7_F_Inst_5__CF_Inst_U1 ( .A1(S_7_F_in3[2]), .A2(S_7_F_in2[3]), 
        .ZN(S_7_F_CF_Out[5]) );
  XNOR2_X1 S_7_F_Inst_6__CF_Inst_U2 ( .A(S_7_F_Inst_6__CF_Inst_n7), .B(
        S_7_F_in3[1]), .ZN(S_7_F_CF_Out[6]) );
  NOR2_X1 S_7_F_Inst_6__CF_Inst_U1 ( .A1(S_7_F_in1[2]), .A2(S_7_F_in3[3]), 
        .ZN(S_7_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_7_F_Inst_7__CF_Inst_U1 ( .A1(S_7_F_in2[2]), .A2(S_7_F_in3[3]), 
        .ZN(S_7_F_CF_Out[7]) );
  OR2_X1 S_7_F_Inst_8__CF_Inst_U1 ( .A1(S_7_F_in3[3]), .A2(S_7_F_in3[2]), .ZN(
        S_7_F_CF_Out[8]) );
  NOR2_X1 S_7_F_Inst_9__CF_Inst_U2 ( .A1(S_7_F_in1[3]), .A2(
        S_7_F_Inst_9__CF_Inst_n3), .ZN(S_7_F_CF_Out[9]) );
  INV_X1 S_7_F_Inst_9__CF_Inst_U1 ( .A(S_7_F_in1[1]), .ZN(
        S_7_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_7_F_Inst_10__CF_Inst_U1 ( .A1(S_7_F_in2[1]), .A2(S_7_F_in1[3]), 
        .ZN(S_7_F_CF_Out[10]) );
  XNOR2_X1 S_7_F_Inst_11__CF_Inst_U2 ( .A(S_7_F_Inst_11__CF_Inst_n3), .B(
        S_7_F_in1[0]), .ZN(S_7_F_CF_Out[11]) );
  NAND2_X1 S_7_F_Inst_11__CF_Inst_U1 ( .A1(S_7_F_in3[1]), .A2(S_7_F_in1[3]), 
        .ZN(S_7_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_7_F_Inst_12__CF_Inst_U2 ( .A(S_7_F_Inst_12__CF_Inst_n3), .B(
        S_7_F_in2[0]), .ZN(S_7_F_CF_Out[12]) );
  NAND2_X1 S_7_F_Inst_12__CF_Inst_U1 ( .A1(S_7_F_in1[1]), .A2(S_7_F_in2[3]), 
        .ZN(S_7_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_7_F_Inst_13__CF_Inst_U2 ( .A1(S_7_F_in2[3]), .A2(
        S_7_F_Inst_13__CF_Inst_n3), .ZN(S_7_F_CF_Out[13]) );
  INV_X1 S_7_F_Inst_13__CF_Inst_U1 ( .A(S_7_F_in2[1]), .ZN(
        S_7_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_7_F_Inst_14__CF_Inst_U1 ( .A1(S_7_F_in3[1]), .A2(S_7_F_in2[3]), 
        .ZN(S_7_F_CF_Out[14]) );
  XNOR2_X1 S_7_F_Inst_15__CF_Inst_U2 ( .A(S_7_F_Inst_15__CF_Inst_n7), .B(
        S_7_F_in3[0]), .ZN(S_7_F_CF_Out[15]) );
  NOR2_X1 S_7_F_Inst_15__CF_Inst_U1 ( .A1(S_7_F_in1[1]), .A2(S_7_F_in3[3]), 
        .ZN(S_7_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_7_F_Inst_16__CF_Inst_U2 ( .A1(S_7_F_in3[3]), .A2(
        S_7_F_Inst_16__CF_Inst_n3), .ZN(S_7_F_CF_Out[16]) );
  INV_X1 S_7_F_Inst_16__CF_Inst_U1 ( .A(S_7_F_in2[1]), .ZN(
        S_7_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_7_F_Inst_17__CF_Inst_U2 ( .A1(S_7_F_in3[1]), .A2(
        S_7_F_Inst_17__CF_Inst_n3), .ZN(S_7_F_CF_Out[17]) );
  INV_X1 S_7_F_Inst_17__CF_Inst_U1 ( .A(S_7_F_in3[3]), .ZN(
        S_7_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_7_F_InstXOR_0__Compression1_U2 ( .A(
        S_7_F_InstXOR_0__Compression1_n3), .B(S_7_F_CF_Reg[2]), .ZN(
        S_7_F_q1[2]) );
  XNOR2_X1 S_7_F_InstXOR_0__Compression1_U1 ( .A(S_7_F_CF_Reg[0]), .B(
        S_7_F_CF_Reg[1]), .ZN(S_7_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_7_F_InstXOR_0__Compression2_U2 ( .A(
        S_7_F_InstXOR_0__Compression2_n3), .B(S_7_F_CF_Reg[5]), .ZN(
        S_7_F_q2[2]) );
  XNOR2_X1 S_7_F_InstXOR_0__Compression2_U1 ( .A(S_7_F_CF_Reg[3]), .B(
        S_7_F_CF_Reg[4]), .ZN(S_7_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_7_F_InstXOR_0__Compression3_U2 ( .A(
        S_7_F_InstXOR_0__Compression3_n3), .B(S_7_F_CF_Reg[8]), .ZN(
        S_7_F_q3[2]) );
  XNOR2_X1 S_7_F_InstXOR_0__Compression3_U1 ( .A(S_7_F_CF_Reg[6]), .B(
        S_7_F_CF_Reg[7]), .ZN(S_7_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_7_F_InstXOR_1__Compression1_U2 ( .A(
        S_7_F_InstXOR_1__Compression1_n3), .B(S_7_F_CF_Reg[11]), .ZN(
        S_7_F_q1[3]) );
  XNOR2_X1 S_7_F_InstXOR_1__Compression1_U1 ( .A(S_7_F_CF_Reg[9]), .B(
        S_7_F_CF_Reg[10]), .ZN(S_7_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_7_F_InstXOR_1__Compression2_U2 ( .A(
        S_7_F_InstXOR_1__Compression2_n3), .B(S_7_F_CF_Reg[14]), .ZN(
        S_7_F_q2[3]) );
  XNOR2_X1 S_7_F_InstXOR_1__Compression2_U1 ( .A(S_7_F_CF_Reg[12]), .B(
        S_7_F_CF_Reg[13]), .ZN(S_7_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_7_F_InstXOR_1__Compression3_U2 ( .A(
        S_7_F_InstXOR_1__Compression3_n3), .B(S_7_F_CF_Reg[17]), .ZN(
        S_7_F_q3[3]) );
  XNOR2_X1 S_7_F_InstXOR_1__Compression3_U1 ( .A(S_7_F_CF_Reg[15]), .B(
        S_7_F_CF_Reg[16]), .ZN(S_7_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_7_G_CF_Reg_reg_0_ ( .D(S_7_G_CF_Out[0]), .CK(CLK), .Q(
        S_7_G_CF_Reg[0]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_1_ ( .D(S_7_G_CF_Out[1]), .CK(CLK), .Q(
        S_7_G_CF_Reg[1]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_2_ ( .D(S_7_G_CF_Out[2]), .CK(CLK), .Q(
        S_7_G_CF_Reg[2]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_3_ ( .D(S_7_G_CF_Out[3]), .CK(CLK), .Q(
        S_7_G_CF_Reg[3]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_4_ ( .D(S_7_G_CF_Out[4]), .CK(CLK), .Q(
        S_7_G_CF_Reg[4]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_5_ ( .D(S_7_G_CF_Out[5]), .CK(CLK), .Q(
        S_7_G_CF_Reg[5]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_6_ ( .D(S_7_G_CF_Out[6]), .CK(CLK), .Q(
        S_7_G_CF_Reg[6]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_7_ ( .D(S_7_G_CF_Out[7]), .CK(CLK), .Q(
        S_7_G_CF_Reg[7]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_8_ ( .D(S_7_G_CF_Out[8]), .CK(CLK), .Q(
        S_7_G_CF_Reg[8]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_9_ ( .D(S_7_G_CF_Out[9]), .CK(CLK), .Q(
        S_7_G_CF_Reg[9]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_10_ ( .D(S_7_G_CF_Out[10]), .CK(CLK), .Q(
        S_7_G_CF_Reg[10]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_11_ ( .D(S_7_G_CF_Out[11]), .CK(CLK), .Q(
        S_7_G_CF_Reg[11]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_12_ ( .D(S_7_G_CF_Out[12]), .CK(CLK), .Q(
        S_7_G_CF_Reg[12]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_13_ ( .D(S_7_G_CF_Out[13]), .CK(CLK), .Q(
        S_7_G_CF_Reg[13]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_14_ ( .D(S_7_G_CF_Out[14]), .CK(CLK), .Q(
        S_7_G_CF_Reg[14]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_15_ ( .D(S_7_G_CF_Out[15]), .CK(CLK), .Q(
        S_7_G_CF_Reg[15]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_16_ ( .D(S_7_G_CF_Out[16]), .CK(CLK), .Q(
        S_7_G_CF_Reg[16]), .QN() );
  DFF_X1 S_7_G_CF_Reg_reg_17_ ( .D(S_7_G_CF_Out[17]), .CK(CLK), .Q(
        S_7_G_CF_Reg[17]), .QN() );
  DFF_X1 S_7_G_out1_reg_2_ ( .D(S_7_Rq1[2]), .CK(CLK), .Q(S_7_G_out1[2]), 
        .QN() );
  DFF_X1 S_7_G_out1_reg_3_ ( .D(S_7_Rq1[3]), .CK(CLK), .Q(S_7_G_out1[3]), 
        .QN() );
  DFF_X1 S_7_G_out2_reg_2_ ( .D(S_7_Rq2[2]), .CK(CLK), .Q(RF2_SHIFTROWS[22]), 
        .QN() );
  DFF_X1 S_7_G_out2_reg_3_ ( .D(S_7_Rq2[3]), .CK(CLK), .Q(RF2_SHIFTROWS[23]), 
        .QN() );
  DFF_X1 S_7_G_out3_reg_2_ ( .D(S_7_Rq3[2]), .CK(CLK), .Q(RF3_SHIFTROWS[22]), 
        .QN() );
  DFF_X1 S_7_G_out3_reg_3_ ( .D(S_7_Rq3[3]), .CK(CLK), .Q(RF3_SHIFTROWS[23]), 
        .QN() );
  AND2_X1 S_7_G_Inst_0__CF_Inst_U1 ( .A1(S_7_Rq1[1]), .A2(S_7_Rq1[3]), .ZN(
        S_7_G_CF_Out[0]) );
  NOR2_X1 S_7_G_Inst_1__CF_Inst_U2 ( .A1(S_7_Rq1[3]), .A2(
        S_7_G_Inst_1__CF_Inst_n3), .ZN(S_7_G_CF_Out[1]) );
  INV_X1 S_7_G_Inst_1__CF_Inst_U1 ( .A(S_7_Rq2[1]), .ZN(
        S_7_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_7_G_Inst_2__CF_Inst_U2 ( .A(S_7_G_Inst_2__CF_Inst_n3), .B(
        S_7_Rq2[0]), .ZN(S_7_G_CF_Out[2]) );
  NAND2_X1 S_7_G_Inst_2__CF_Inst_U1 ( .A1(S_7_Rq1[1]), .A2(S_7_Rq2[3]), .ZN(
        S_7_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_7_G_Inst_3__CF_Inst_U3 ( .A(S_7_Rq1[0]), .B(
        S_7_G_Inst_3__CF_Inst_n6), .ZN(S_7_G_CF_Out[3]) );
  NAND2_X1 S_7_G_Inst_3__CF_Inst_U2 ( .A1(S_7_Rq3[1]), .A2(
        S_7_G_Inst_3__CF_Inst_n5), .ZN(S_7_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_7_G_Inst_3__CF_Inst_U1 ( .A(S_7_Rq1[3]), .ZN(
        S_7_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_7_G_Inst_4__CF_Inst_U1 ( .A1(S_7_Rq2[1]), .A2(S_7_Rq2[3]), .ZN(
        S_7_G_CF_Out[4]) );
  OR2_X1 S_7_G_Inst_5__CF_Inst_U1 ( .A1(S_7_Rq3[3]), .A2(S_7_Rq2[1]), .ZN(
        S_7_G_CF_Out[5]) );
  AND2_X1 S_7_G_Inst_6__CF_Inst_U1 ( .A1(S_7_Rq3[1]), .A2(S_7_Rq2[3]), .ZN(
        S_7_G_CF_Out[6]) );
  XNOR2_X1 S_7_G_Inst_7__CF_Inst_U2 ( .A(S_7_G_Inst_7__CF_Inst_n3), .B(
        S_7_Rq3[0]), .ZN(S_7_G_CF_Out[7]) );
  NAND2_X1 S_7_G_Inst_7__CF_Inst_U1 ( .A1(S_7_Rq1[1]), .A2(S_7_Rq3[3]), .ZN(
        S_7_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_7_G_Inst_8__CF_Inst_U1 ( .A1(S_7_Rq3[3]), .A2(S_7_Rq3[1]), .ZN(
        S_7_G_CF_Out[8]) );
  NOR2_X1 S_7_G_Inst_9__CF_Inst_U2 ( .A1(S_7_Rq1[3]), .A2(
        S_7_G_Inst_9__CF_Inst_n3), .ZN(S_7_G_CF_Out[9]) );
  INV_X1 S_7_G_Inst_9__CF_Inst_U1 ( .A(S_7_Rq1[2]), .ZN(
        S_7_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_7_G_Inst_10__CF_Inst_U2 ( .A1(S_7_Rq2[2]), .A2(
        S_7_G_Inst_10__CF_Inst_n3), .ZN(S_7_G_CF_Out[10]) );
  INV_X1 S_7_G_Inst_10__CF_Inst_U1 ( .A(S_7_Rq1[3]), .ZN(
        S_7_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_7_G_Inst_11__CF_Inst_U3 ( .A(S_7_Rq1[1]), .B(
        S_7_G_Inst_11__CF_Inst_n6), .ZN(S_7_G_CF_Out[11]) );
  NAND2_X1 S_7_G_Inst_11__CF_Inst_U2 ( .A1(S_7_Rq1[3]), .A2(
        S_7_G_Inst_11__CF_Inst_n5), .ZN(S_7_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_7_G_Inst_11__CF_Inst_U1 ( .A(S_7_Rq3[2]), .ZN(
        S_7_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_7_G_Inst_12__CF_Inst_U2 ( .A1(S_7_Rq2[3]), .A2(
        S_7_G_Inst_12__CF_Inst_n3), .ZN(S_7_G_CF_Out[12]) );
  INV_X1 S_7_G_Inst_12__CF_Inst_U1 ( .A(S_7_Rq1[2]), .ZN(
        S_7_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_7_G_Inst_13__CF_Inst_U1 ( .A1(S_7_Rq2[2]), .A2(S_7_Rq2[3]), .ZN(
        S_7_G_CF_Out[13]) );
  XNOR2_X1 S_7_G_Inst_14__CF_Inst_U3 ( .A(S_7_Rq2[1]), .B(
        S_7_G_Inst_14__CF_Inst_n6), .ZN(S_7_G_CF_Out[14]) );
  NAND2_X1 S_7_G_Inst_14__CF_Inst_U2 ( .A1(S_7_Rq3[2]), .A2(
        S_7_G_Inst_14__CF_Inst_n5), .ZN(S_7_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_7_G_Inst_14__CF_Inst_U1 ( .A(S_7_Rq2[3]), .ZN(
        S_7_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_7_G_Inst_15__CF_Inst_U2 ( .A(S_7_G_Inst_15__CF_Inst_n3), .B(
        S_7_Rq3[1]), .ZN(S_7_G_CF_Out[15]) );
  NAND2_X1 S_7_G_Inst_15__CF_Inst_U1 ( .A1(S_7_Rq1[2]), .A2(S_7_Rq3[3]), .ZN(
        S_7_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_7_G_Inst_16__CF_Inst_U1 ( .A1(S_7_Rq2[2]), .A2(S_7_Rq3[3]), .ZN(
        S_7_G_CF_Out[16]) );
  NOR2_X1 S_7_G_Inst_17__CF_Inst_U2 ( .A1(S_7_Rq3[3]), .A2(
        S_7_G_Inst_17__CF_Inst_n3), .ZN(S_7_G_CF_Out[17]) );
  INV_X1 S_7_G_Inst_17__CF_Inst_U1 ( .A(S_7_Rq3[2]), .ZN(
        S_7_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_7_G_InstXOR_0__Compression1_U2 ( .A(
        S_7_G_InstXOR_0__Compression1_n3), .B(S_7_G_CF_Reg[2]), .ZN(
        S_7_G_out1[0]) );
  XNOR2_X1 S_7_G_InstXOR_0__Compression1_U1 ( .A(S_7_G_CF_Reg[0]), .B(
        S_7_G_CF_Reg[1]), .ZN(S_7_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_7_G_InstXOR_0__Compression2_U2 ( .A(
        S_7_G_InstXOR_0__Compression2_n3), .B(S_7_G_CF_Reg[5]), .ZN(
        SUB_OUT2[29]) );
  XNOR2_X1 S_7_G_InstXOR_0__Compression2_U1 ( .A(S_7_G_CF_Reg[3]), .B(
        S_7_G_CF_Reg[4]), .ZN(S_7_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_7_G_InstXOR_0__Compression3_U2 ( .A(
        S_7_G_InstXOR_0__Compression3_n3), .B(S_7_G_CF_Reg[8]), .ZN(
        SUB_OUT3[29]) );
  XNOR2_X1 S_7_G_InstXOR_0__Compression3_U1 ( .A(S_7_G_CF_Reg[6]), .B(
        S_7_G_CF_Reg[7]), .ZN(S_7_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_7_G_InstXOR_1__Compression1_U2 ( .A(
        S_7_G_InstXOR_1__Compression1_n3), .B(S_7_G_CF_Reg[11]), .ZN(
        S_7_G_out1[1]) );
  XNOR2_X1 S_7_G_InstXOR_1__Compression1_U1 ( .A(S_7_G_CF_Reg[9]), .B(
        S_7_G_CF_Reg[10]), .ZN(S_7_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_7_G_InstXOR_1__Compression2_U2 ( .A(
        S_7_G_InstXOR_1__Compression2_n3), .B(S_7_G_CF_Reg[14]), .ZN(
        RF2_SHIFTROWS[20]) );
  XNOR2_X1 S_7_G_InstXOR_1__Compression2_U1 ( .A(S_7_G_CF_Reg[12]), .B(
        S_7_G_CF_Reg[13]), .ZN(S_7_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_7_G_InstXOR_1__Compression3_U2 ( .A(
        S_7_G_InstXOR_1__Compression3_n3), .B(S_7_G_CF_Reg[17]), .ZN(
        RF3_SHIFTROWS[20]) );
  XNOR2_X1 S_7_G_InstXOR_1__Compression3_U1 ( .A(S_7_G_CF_Reg[15]), .B(
        S_7_G_CF_Reg[16]), .ZN(S_7_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_7_OutputAffine_U4 ( .A(S_7_G_out1[3]), .ZN(RF1_SHIFTROWS[23]) );
  INV_X1 S_7_OutputAffine_U3 ( .A(S_7_G_out1[2]), .ZN(RF1_SHIFTROWS[22]) );
  INV_X1 S_7_OutputAffine_U2 ( .A(S_7_G_out1[1]), .ZN(RF1_SHIFTROWS[20]) );
  INV_X1 S_7_OutputAffine_U1 ( .A(S_7_G_out1[0]), .ZN(SUB_OUT1[29]) );
  DFF_X1 S_8_Rq3_reg_0_ ( .D(S_8_q3[0]), .CK(CLK), .Q(S_8_Rq3[0]), .QN() );
  DFF_X1 S_8_Rq3_reg_1_ ( .D(S_8_q3[1]), .CK(CLK), .Q(S_8_Rq3[1]), .QN() );
  DFF_X1 S_8_Rq3_reg_2_ ( .D(S_8_q3[2]), .CK(CLK), .Q(S_8_Rq3[2]), .QN() );
  DFF_X1 S_8_Rq3_reg_3_ ( .D(S_8_q3[3]), .CK(CLK), .Q(S_8_Rq3[3]), .QN() );
  DFF_X1 S_8_Rq2_reg_0_ ( .D(S_8_q2[0]), .CK(CLK), .Q(S_8_Rq2[0]), .QN() );
  DFF_X1 S_8_Rq2_reg_1_ ( .D(S_8_q2[1]), .CK(CLK), .Q(S_8_Rq2[1]), .QN() );
  DFF_X1 S_8_Rq2_reg_2_ ( .D(S_8_q2[2]), .CK(CLK), .Q(S_8_Rq2[2]), .QN() );
  DFF_X1 S_8_Rq2_reg_3_ ( .D(S_8_q2[3]), .CK(CLK), .Q(S_8_Rq2[3]), .QN() );
  DFF_X1 S_8_Rq1_reg_0_ ( .D(S_8_q1[0]), .CK(CLK), .Q(S_8_Rq1[0]), .QN() );
  DFF_X1 S_8_Rq1_reg_1_ ( .D(S_8_q1[1]), .CK(CLK), .Q(S_8_Rq1[1]), .QN() );
  DFF_X1 S_8_Rq1_reg_2_ ( .D(S_8_q1[2]), .CK(CLK), .Q(S_8_Rq1[2]), .QN() );
  DFF_X1 S_8_Rq1_reg_3_ ( .D(S_8_q1[3]), .CK(CLK), .Q(S_8_Rq1[3]), .QN() );
  INV_X1 S_8_InputAffine_U4 ( .A(SUB_IN1[32]), .ZN(S_8_F_in1[0]) );
  INV_X1 S_8_InputAffine_U3 ( .A(SUB_IN1[34]), .ZN(S_8_F_in1[3]) );
  INV_X1 S_8_InputAffine_U2 ( .A(SUB_IN1[35]), .ZN(S_8_F_in1[1]) );
  INV_X1 S_8_InputAffine_U1 ( .A(SUB_IN1[33]), .ZN(S_8_F_in1[2]) );
  XNOR2_X1 S_8_F_U18 ( .A(S_8_F_n12), .B(FRESH[67]), .ZN(S_8_q3[3]) );
  XNOR2_X1 S_8_F_U17 ( .A(FRESH[66]), .B(S_8_F_q3[3]), .ZN(S_8_F_n12) );
  XNOR2_X1 S_8_F_U16 ( .A(S_8_F_n11), .B(FRESH[65]), .ZN(S_8_q3[2]) );
  XNOR2_X1 S_8_F_U15 ( .A(FRESH[64]), .B(S_8_F_q3[2]), .ZN(S_8_F_n11) );
  XOR2_X1 S_8_F_U14 ( .A(FRESH[67]), .B(S_8_F_q2[3]), .Z(S_8_q2[3]) );
  XOR2_X1 S_8_F_U13 ( .A(FRESH[65]), .B(S_8_F_q2[2]), .Z(S_8_q2[2]) );
  XOR2_X1 S_8_F_U12 ( .A(FRESH[66]), .B(S_8_F_q1[3]), .Z(S_8_q1[3]) );
  XOR2_X1 S_8_F_U11 ( .A(FRESH[64]), .B(S_8_F_q1[2]), .Z(S_8_q1[2]) );
  XNOR2_X1 S_8_F_U10 ( .A(S_8_F_n10), .B(FRESH[69]), .ZN(S_8_F_N5) );
  XNOR2_X1 S_8_F_U9 ( .A(S_8_F_in3[3]), .B(FRESH[68]), .ZN(S_8_F_n10) );
  XOR2_X1 S_8_F_U8 ( .A(FRESH[69]), .B(S_8_F_in2[3]), .Z(S_8_F_N4) );
  XOR2_X1 S_8_F_U7 ( .A(FRESH[68]), .B(S_8_F_in1[3]), .Z(S_8_F_N3) );
  XNOR2_X1 S_8_F_U6 ( .A(S_8_F_n9), .B(FRESH[71]), .ZN(S_8_F_N2) );
  XNOR2_X1 S_8_F_U5 ( .A(S_8_F_in3[2]), .B(FRESH[70]), .ZN(S_8_F_n9) );
  XOR2_X1 S_8_F_U4 ( .A(FRESH[71]), .B(S_8_F_in2[2]), .Z(S_8_F_N1) );
  XOR2_X1 S_8_F_U3 ( .A(FRESH[70]), .B(S_8_F_in1[2]), .Z(S_8_F_N0) );
  DFF_X1 S_8_F_CF_Reg_reg_0_ ( .D(S_8_F_CF_Out[0]), .CK(CLK), .Q(
        S_8_F_CF_Reg[0]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_1_ ( .D(S_8_F_CF_Out[1]), .CK(CLK), .Q(
        S_8_F_CF_Reg[1]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_2_ ( .D(S_8_F_CF_Out[2]), .CK(CLK), .Q(
        S_8_F_CF_Reg[2]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_3_ ( .D(S_8_F_CF_Out[3]), .CK(CLK), .Q(
        S_8_F_CF_Reg[3]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_4_ ( .D(S_8_F_CF_Out[4]), .CK(CLK), .Q(
        S_8_F_CF_Reg[4]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_5_ ( .D(S_8_F_CF_Out[5]), .CK(CLK), .Q(
        S_8_F_CF_Reg[5]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_6_ ( .D(S_8_F_CF_Out[6]), .CK(CLK), .Q(
        S_8_F_CF_Reg[6]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_7_ ( .D(S_8_F_CF_Out[7]), .CK(CLK), .Q(
        S_8_F_CF_Reg[7]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_8_ ( .D(S_8_F_CF_Out[8]), .CK(CLK), .Q(
        S_8_F_CF_Reg[8]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_9_ ( .D(S_8_F_CF_Out[9]), .CK(CLK), .Q(
        S_8_F_CF_Reg[9]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_10_ ( .D(S_8_F_CF_Out[10]), .CK(CLK), .Q(
        S_8_F_CF_Reg[10]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_11_ ( .D(S_8_F_CF_Out[11]), .CK(CLK), .Q(
        S_8_F_CF_Reg[11]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_12_ ( .D(S_8_F_CF_Out[12]), .CK(CLK), .Q(
        S_8_F_CF_Reg[12]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_13_ ( .D(S_8_F_CF_Out[13]), .CK(CLK), .Q(
        S_8_F_CF_Reg[13]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_14_ ( .D(S_8_F_CF_Out[14]), .CK(CLK), .Q(
        S_8_F_CF_Reg[14]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_15_ ( .D(S_8_F_CF_Out[15]), .CK(CLK), .Q(
        S_8_F_CF_Reg[15]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_16_ ( .D(S_8_F_CF_Out[16]), .CK(CLK), .Q(
        S_8_F_CF_Reg[16]), .QN() );
  DFF_X1 S_8_F_CF_Reg_reg_17_ ( .D(S_8_F_CF_Out[17]), .CK(CLK), .Q(
        S_8_F_CF_Reg[17]), .QN() );
  DFF_X1 S_8_F_out2_reg_0_ ( .D(S_8_F_N4), .CK(CLK), .Q(S_8_q2[0]), .QN() );
  DFF_X1 S_8_F_out2_reg_1_ ( .D(S_8_F_N1), .CK(CLK), .Q(S_8_q2[1]), .QN() );
  DFF_X1 S_8_F_out3_reg_0_ ( .D(S_8_F_N5), .CK(CLK), .Q(S_8_q3[0]), .QN() );
  DFF_X1 S_8_F_out3_reg_1_ ( .D(S_8_F_N2), .CK(CLK), .Q(S_8_q3[1]), .QN() );
  DFF_X1 S_8_F_out1_reg_0_ ( .D(S_8_F_N3), .CK(CLK), .Q(S_8_q1[0]), .QN() );
  DFF_X1 S_8_F_out1_reg_1_ ( .D(S_8_F_N0), .CK(CLK), .Q(S_8_q1[1]), .QN() );
  NOR2_X1 S_8_F_Inst_0__CF_Inst_U2 ( .A1(S_8_F_in1[2]), .A2(
        S_8_F_Inst_0__CF_Inst_n3), .ZN(S_8_F_CF_Out[0]) );
  INV_X1 S_8_F_Inst_0__CF_Inst_U1 ( .A(S_8_F_in1[3]), .ZN(
        S_8_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_8_F_Inst_1__CF_Inst_U2 ( .A(S_8_F_Inst_1__CF_Inst_n3), .B(
        S_8_F_in1[1]), .ZN(S_8_F_CF_Out[1]) );
  NAND2_X1 S_8_F_Inst_1__CF_Inst_U1 ( .A1(S_8_F_in2[2]), .A2(S_8_F_in1[3]), 
        .ZN(S_8_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_8_F_Inst_2__CF_Inst_U1 ( .A1(S_8_F_in1[3]), .A2(S_8_F_in3[2]), .ZN(
        S_8_F_CF_Out[2]) );
  NOR2_X1 S_8_F_Inst_3__CF_Inst_U2 ( .A1(S_8_F_in2[3]), .A2(
        S_8_F_Inst_3__CF_Inst_n3), .ZN(S_8_F_CF_Out[3]) );
  INV_X1 S_8_F_Inst_3__CF_Inst_U1 ( .A(S_8_F_in1[2]), .ZN(
        S_8_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_8_F_Inst_4__CF_Inst_U2 ( .A(S_8_F_Inst_4__CF_Inst_n3), .B(
        S_8_F_in2[1]), .ZN(S_8_F_CF_Out[4]) );
  NAND2_X1 S_8_F_Inst_4__CF_Inst_U1 ( .A1(S_8_F_in2[2]), .A2(S_8_F_in2[3]), 
        .ZN(S_8_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_8_F_Inst_5__CF_Inst_U1 ( .A1(S_8_F_in3[2]), .A2(S_8_F_in2[3]), 
        .ZN(S_8_F_CF_Out[5]) );
  XNOR2_X1 S_8_F_Inst_6__CF_Inst_U2 ( .A(S_8_F_Inst_6__CF_Inst_n7), .B(
        S_8_F_in3[1]), .ZN(S_8_F_CF_Out[6]) );
  NOR2_X1 S_8_F_Inst_6__CF_Inst_U1 ( .A1(S_8_F_in1[2]), .A2(S_8_F_in3[3]), 
        .ZN(S_8_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_8_F_Inst_7__CF_Inst_U1 ( .A1(S_8_F_in2[2]), .A2(S_8_F_in3[3]), 
        .ZN(S_8_F_CF_Out[7]) );
  OR2_X1 S_8_F_Inst_8__CF_Inst_U1 ( .A1(S_8_F_in3[3]), .A2(S_8_F_in3[2]), .ZN(
        S_8_F_CF_Out[8]) );
  NOR2_X1 S_8_F_Inst_9__CF_Inst_U2 ( .A1(S_8_F_in1[3]), .A2(
        S_8_F_Inst_9__CF_Inst_n3), .ZN(S_8_F_CF_Out[9]) );
  INV_X1 S_8_F_Inst_9__CF_Inst_U1 ( .A(S_8_F_in1[1]), .ZN(
        S_8_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_8_F_Inst_10__CF_Inst_U1 ( .A1(S_8_F_in2[1]), .A2(S_8_F_in1[3]), 
        .ZN(S_8_F_CF_Out[10]) );
  XNOR2_X1 S_8_F_Inst_11__CF_Inst_U2 ( .A(S_8_F_Inst_11__CF_Inst_n3), .B(
        S_8_F_in1[0]), .ZN(S_8_F_CF_Out[11]) );
  NAND2_X1 S_8_F_Inst_11__CF_Inst_U1 ( .A1(S_8_F_in3[1]), .A2(S_8_F_in1[3]), 
        .ZN(S_8_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_8_F_Inst_12__CF_Inst_U2 ( .A(S_8_F_Inst_12__CF_Inst_n3), .B(
        S_8_F_in2[0]), .ZN(S_8_F_CF_Out[12]) );
  NAND2_X1 S_8_F_Inst_12__CF_Inst_U1 ( .A1(S_8_F_in1[1]), .A2(S_8_F_in2[3]), 
        .ZN(S_8_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_8_F_Inst_13__CF_Inst_U2 ( .A1(S_8_F_in2[3]), .A2(
        S_8_F_Inst_13__CF_Inst_n3), .ZN(S_8_F_CF_Out[13]) );
  INV_X1 S_8_F_Inst_13__CF_Inst_U1 ( .A(S_8_F_in2[1]), .ZN(
        S_8_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_8_F_Inst_14__CF_Inst_U1 ( .A1(S_8_F_in3[1]), .A2(S_8_F_in2[3]), 
        .ZN(S_8_F_CF_Out[14]) );
  XNOR2_X1 S_8_F_Inst_15__CF_Inst_U2 ( .A(S_8_F_Inst_15__CF_Inst_n7), .B(
        S_8_F_in3[0]), .ZN(S_8_F_CF_Out[15]) );
  NOR2_X1 S_8_F_Inst_15__CF_Inst_U1 ( .A1(S_8_F_in1[1]), .A2(S_8_F_in3[3]), 
        .ZN(S_8_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_8_F_Inst_16__CF_Inst_U2 ( .A1(S_8_F_in3[3]), .A2(
        S_8_F_Inst_16__CF_Inst_n3), .ZN(S_8_F_CF_Out[16]) );
  INV_X1 S_8_F_Inst_16__CF_Inst_U1 ( .A(S_8_F_in2[1]), .ZN(
        S_8_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_8_F_Inst_17__CF_Inst_U2 ( .A1(S_8_F_in3[1]), .A2(
        S_8_F_Inst_17__CF_Inst_n3), .ZN(S_8_F_CF_Out[17]) );
  INV_X1 S_8_F_Inst_17__CF_Inst_U1 ( .A(S_8_F_in3[3]), .ZN(
        S_8_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_8_F_InstXOR_0__Compression1_U2 ( .A(
        S_8_F_InstXOR_0__Compression1_n3), .B(S_8_F_CF_Reg[2]), .ZN(
        S_8_F_q1[2]) );
  XNOR2_X1 S_8_F_InstXOR_0__Compression1_U1 ( .A(S_8_F_CF_Reg[0]), .B(
        S_8_F_CF_Reg[1]), .ZN(S_8_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_8_F_InstXOR_0__Compression2_U2 ( .A(
        S_8_F_InstXOR_0__Compression2_n3), .B(S_8_F_CF_Reg[5]), .ZN(
        S_8_F_q2[2]) );
  XNOR2_X1 S_8_F_InstXOR_0__Compression2_U1 ( .A(S_8_F_CF_Reg[3]), .B(
        S_8_F_CF_Reg[4]), .ZN(S_8_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_8_F_InstXOR_0__Compression3_U2 ( .A(
        S_8_F_InstXOR_0__Compression3_n3), .B(S_8_F_CF_Reg[8]), .ZN(
        S_8_F_q3[2]) );
  XNOR2_X1 S_8_F_InstXOR_0__Compression3_U1 ( .A(S_8_F_CF_Reg[6]), .B(
        S_8_F_CF_Reg[7]), .ZN(S_8_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_8_F_InstXOR_1__Compression1_U2 ( .A(
        S_8_F_InstXOR_1__Compression1_n3), .B(S_8_F_CF_Reg[11]), .ZN(
        S_8_F_q1[3]) );
  XNOR2_X1 S_8_F_InstXOR_1__Compression1_U1 ( .A(S_8_F_CF_Reg[9]), .B(
        S_8_F_CF_Reg[10]), .ZN(S_8_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_8_F_InstXOR_1__Compression2_U2 ( .A(
        S_8_F_InstXOR_1__Compression2_n3), .B(S_8_F_CF_Reg[14]), .ZN(
        S_8_F_q2[3]) );
  XNOR2_X1 S_8_F_InstXOR_1__Compression2_U1 ( .A(S_8_F_CF_Reg[12]), .B(
        S_8_F_CF_Reg[13]), .ZN(S_8_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_8_F_InstXOR_1__Compression3_U2 ( .A(
        S_8_F_InstXOR_1__Compression3_n3), .B(S_8_F_CF_Reg[17]), .ZN(
        S_8_F_q3[3]) );
  XNOR2_X1 S_8_F_InstXOR_1__Compression3_U1 ( .A(S_8_F_CF_Reg[15]), .B(
        S_8_F_CF_Reg[16]), .ZN(S_8_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_8_G_CF_Reg_reg_0_ ( .D(S_8_G_CF_Out[0]), .CK(CLK), .Q(
        S_8_G_CF_Reg[0]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_1_ ( .D(S_8_G_CF_Out[1]), .CK(CLK), .Q(
        S_8_G_CF_Reg[1]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_2_ ( .D(S_8_G_CF_Out[2]), .CK(CLK), .Q(
        S_8_G_CF_Reg[2]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_3_ ( .D(S_8_G_CF_Out[3]), .CK(CLK), .Q(
        S_8_G_CF_Reg[3]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_4_ ( .D(S_8_G_CF_Out[4]), .CK(CLK), .Q(
        S_8_G_CF_Reg[4]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_5_ ( .D(S_8_G_CF_Out[5]), .CK(CLK), .Q(
        S_8_G_CF_Reg[5]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_6_ ( .D(S_8_G_CF_Out[6]), .CK(CLK), .Q(
        S_8_G_CF_Reg[6]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_7_ ( .D(S_8_G_CF_Out[7]), .CK(CLK), .Q(
        S_8_G_CF_Reg[7]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_8_ ( .D(S_8_G_CF_Out[8]), .CK(CLK), .Q(
        S_8_G_CF_Reg[8]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_9_ ( .D(S_8_G_CF_Out[9]), .CK(CLK), .Q(
        S_8_G_CF_Reg[9]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_10_ ( .D(S_8_G_CF_Out[10]), .CK(CLK), .Q(
        S_8_G_CF_Reg[10]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_11_ ( .D(S_8_G_CF_Out[11]), .CK(CLK), .Q(
        S_8_G_CF_Reg[11]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_12_ ( .D(S_8_G_CF_Out[12]), .CK(CLK), .Q(
        S_8_G_CF_Reg[12]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_13_ ( .D(S_8_G_CF_Out[13]), .CK(CLK), .Q(
        S_8_G_CF_Reg[13]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_14_ ( .D(S_8_G_CF_Out[14]), .CK(CLK), .Q(
        S_8_G_CF_Reg[14]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_15_ ( .D(S_8_G_CF_Out[15]), .CK(CLK), .Q(
        S_8_G_CF_Reg[15]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_16_ ( .D(S_8_G_CF_Out[16]), .CK(CLK), .Q(
        S_8_G_CF_Reg[16]), .QN() );
  DFF_X1 S_8_G_CF_Reg_reg_17_ ( .D(S_8_G_CF_Out[17]), .CK(CLK), .Q(
        S_8_G_CF_Reg[17]), .QN() );
  DFF_X1 S_8_G_out1_reg_2_ ( .D(S_8_Rq1[2]), .CK(CLK), .Q(S_8_G_out1[2]), 
        .QN() );
  DFF_X1 S_8_G_out1_reg_3_ ( .D(S_8_Rq1[3]), .CK(CLK), .Q(S_8_G_out1[3]), 
        .QN() );
  DFF_X1 S_8_G_out2_reg_2_ ( .D(S_8_Rq2[2]), .CK(CLK), .Q(SUB_OUT2[34]), .QN()
         );
  DFF_X1 S_8_G_out2_reg_3_ ( .D(S_8_Rq2[3]), .CK(CLK), .Q(SUB_OUT2[35]), .QN()
         );
  DFF_X1 S_8_G_out3_reg_2_ ( .D(S_8_Rq3[2]), .CK(CLK), .Q(SUB_OUT3[34]), .QN()
         );
  DFF_X1 S_8_G_out3_reg_3_ ( .D(S_8_Rq3[3]), .CK(CLK), .Q(SUB_OUT3[35]), .QN()
         );
  AND2_X1 S_8_G_Inst_0__CF_Inst_U1 ( .A1(S_8_Rq1[1]), .A2(S_8_Rq1[3]), .ZN(
        S_8_G_CF_Out[0]) );
  NOR2_X1 S_8_G_Inst_1__CF_Inst_U2 ( .A1(S_8_Rq1[3]), .A2(
        S_8_G_Inst_1__CF_Inst_n3), .ZN(S_8_G_CF_Out[1]) );
  INV_X1 S_8_G_Inst_1__CF_Inst_U1 ( .A(S_8_Rq2[1]), .ZN(
        S_8_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_8_G_Inst_2__CF_Inst_U2 ( .A(S_8_G_Inst_2__CF_Inst_n3), .B(
        S_8_Rq2[0]), .ZN(S_8_G_CF_Out[2]) );
  NAND2_X1 S_8_G_Inst_2__CF_Inst_U1 ( .A1(S_8_Rq1[1]), .A2(S_8_Rq2[3]), .ZN(
        S_8_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_8_G_Inst_3__CF_Inst_U3 ( .A(S_8_Rq1[0]), .B(
        S_8_G_Inst_3__CF_Inst_n6), .ZN(S_8_G_CF_Out[3]) );
  NAND2_X1 S_8_G_Inst_3__CF_Inst_U2 ( .A1(S_8_Rq3[1]), .A2(
        S_8_G_Inst_3__CF_Inst_n5), .ZN(S_8_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_8_G_Inst_3__CF_Inst_U1 ( .A(S_8_Rq1[3]), .ZN(
        S_8_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_8_G_Inst_4__CF_Inst_U1 ( .A1(S_8_Rq2[1]), .A2(S_8_Rq2[3]), .ZN(
        S_8_G_CF_Out[4]) );
  OR2_X1 S_8_G_Inst_5__CF_Inst_U1 ( .A1(S_8_Rq3[3]), .A2(S_8_Rq2[1]), .ZN(
        S_8_G_CF_Out[5]) );
  AND2_X1 S_8_G_Inst_6__CF_Inst_U1 ( .A1(S_8_Rq3[1]), .A2(S_8_Rq2[3]), .ZN(
        S_8_G_CF_Out[6]) );
  XNOR2_X1 S_8_G_Inst_7__CF_Inst_U2 ( .A(S_8_G_Inst_7__CF_Inst_n3), .B(
        S_8_Rq3[0]), .ZN(S_8_G_CF_Out[7]) );
  NAND2_X1 S_8_G_Inst_7__CF_Inst_U1 ( .A1(S_8_Rq1[1]), .A2(S_8_Rq3[3]), .ZN(
        S_8_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_8_G_Inst_8__CF_Inst_U1 ( .A1(S_8_Rq3[3]), .A2(S_8_Rq3[1]), .ZN(
        S_8_G_CF_Out[8]) );
  NOR2_X1 S_8_G_Inst_9__CF_Inst_U2 ( .A1(S_8_Rq1[3]), .A2(
        S_8_G_Inst_9__CF_Inst_n3), .ZN(S_8_G_CF_Out[9]) );
  INV_X1 S_8_G_Inst_9__CF_Inst_U1 ( .A(S_8_Rq1[2]), .ZN(
        S_8_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_8_G_Inst_10__CF_Inst_U2 ( .A1(S_8_Rq2[2]), .A2(
        S_8_G_Inst_10__CF_Inst_n3), .ZN(S_8_G_CF_Out[10]) );
  INV_X1 S_8_G_Inst_10__CF_Inst_U1 ( .A(S_8_Rq1[3]), .ZN(
        S_8_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_8_G_Inst_11__CF_Inst_U3 ( .A(S_8_Rq1[1]), .B(
        S_8_G_Inst_11__CF_Inst_n6), .ZN(S_8_G_CF_Out[11]) );
  NAND2_X1 S_8_G_Inst_11__CF_Inst_U2 ( .A1(S_8_Rq1[3]), .A2(
        S_8_G_Inst_11__CF_Inst_n5), .ZN(S_8_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_8_G_Inst_11__CF_Inst_U1 ( .A(S_8_Rq3[2]), .ZN(
        S_8_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_8_G_Inst_12__CF_Inst_U2 ( .A1(S_8_Rq2[3]), .A2(
        S_8_G_Inst_12__CF_Inst_n3), .ZN(S_8_G_CF_Out[12]) );
  INV_X1 S_8_G_Inst_12__CF_Inst_U1 ( .A(S_8_Rq1[2]), .ZN(
        S_8_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_8_G_Inst_13__CF_Inst_U1 ( .A1(S_8_Rq2[2]), .A2(S_8_Rq2[3]), .ZN(
        S_8_G_CF_Out[13]) );
  XNOR2_X1 S_8_G_Inst_14__CF_Inst_U3 ( .A(S_8_Rq2[1]), .B(
        S_8_G_Inst_14__CF_Inst_n6), .ZN(S_8_G_CF_Out[14]) );
  NAND2_X1 S_8_G_Inst_14__CF_Inst_U2 ( .A1(S_8_Rq3[2]), .A2(
        S_8_G_Inst_14__CF_Inst_n5), .ZN(S_8_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_8_G_Inst_14__CF_Inst_U1 ( .A(S_8_Rq2[3]), .ZN(
        S_8_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_8_G_Inst_15__CF_Inst_U2 ( .A(S_8_G_Inst_15__CF_Inst_n3), .B(
        S_8_Rq3[1]), .ZN(S_8_G_CF_Out[15]) );
  NAND2_X1 S_8_G_Inst_15__CF_Inst_U1 ( .A1(S_8_Rq1[2]), .A2(S_8_Rq3[3]), .ZN(
        S_8_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_8_G_Inst_16__CF_Inst_U1 ( .A1(S_8_Rq2[2]), .A2(S_8_Rq3[3]), .ZN(
        S_8_G_CF_Out[16]) );
  NOR2_X1 S_8_G_Inst_17__CF_Inst_U2 ( .A1(S_8_Rq3[3]), .A2(
        S_8_G_Inst_17__CF_Inst_n3), .ZN(S_8_G_CF_Out[17]) );
  INV_X1 S_8_G_Inst_17__CF_Inst_U1 ( .A(S_8_Rq3[2]), .ZN(
        S_8_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_8_G_InstXOR_0__Compression1_U2 ( .A(
        S_8_G_InstXOR_0__Compression1_n3), .B(S_8_G_CF_Reg[2]), .ZN(
        S_8_G_out1[0]) );
  XNOR2_X1 S_8_G_InstXOR_0__Compression1_U1 ( .A(S_8_G_CF_Reg[0]), .B(
        S_8_G_CF_Reg[1]), .ZN(S_8_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_8_G_InstXOR_0__Compression2_U2 ( .A(
        S_8_G_InstXOR_0__Compression2_n3), .B(S_8_G_CF_Reg[5]), .ZN(
        SUB_OUT2[33]) );
  XNOR2_X1 S_8_G_InstXOR_0__Compression2_U1 ( .A(S_8_G_CF_Reg[3]), .B(
        S_8_G_CF_Reg[4]), .ZN(S_8_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_8_G_InstXOR_0__Compression3_U2 ( .A(
        S_8_G_InstXOR_0__Compression3_n3), .B(S_8_G_CF_Reg[8]), .ZN(
        SUB_OUT3[33]) );
  XNOR2_X1 S_8_G_InstXOR_0__Compression3_U1 ( .A(S_8_G_CF_Reg[6]), .B(
        S_8_G_CF_Reg[7]), .ZN(S_8_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_8_G_InstXOR_1__Compression1_U2 ( .A(
        S_8_G_InstXOR_1__Compression1_n3), .B(S_8_G_CF_Reg[11]), .ZN(
        S_8_G_out1[1]) );
  XNOR2_X1 S_8_G_InstXOR_1__Compression1_U1 ( .A(S_8_G_CF_Reg[9]), .B(
        S_8_G_CF_Reg[10]), .ZN(S_8_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_8_G_InstXOR_1__Compression2_U2 ( .A(
        S_8_G_InstXOR_1__Compression2_n3), .B(S_8_G_CF_Reg[14]), .ZN(
        SUB_OUT2[32]) );
  XNOR2_X1 S_8_G_InstXOR_1__Compression2_U1 ( .A(S_8_G_CF_Reg[12]), .B(
        S_8_G_CF_Reg[13]), .ZN(S_8_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_8_G_InstXOR_1__Compression3_U2 ( .A(
        S_8_G_InstXOR_1__Compression3_n3), .B(S_8_G_CF_Reg[17]), .ZN(
        SUB_OUT3[32]) );
  XNOR2_X1 S_8_G_InstXOR_1__Compression3_U1 ( .A(S_8_G_CF_Reg[15]), .B(
        S_8_G_CF_Reg[16]), .ZN(S_8_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_8_OutputAffine_U4 ( .A(S_8_G_out1[3]), .ZN(SUB_OUT1[35]) );
  INV_X1 S_8_OutputAffine_U3 ( .A(S_8_G_out1[2]), .ZN(SUB_OUT1[34]) );
  INV_X1 S_8_OutputAffine_U2 ( .A(S_8_G_out1[1]), .ZN(SUB_OUT1[32]) );
  INV_X1 S_8_OutputAffine_U1 ( .A(S_8_G_out1[0]), .ZN(SUB_OUT1[33]) );
  DFF_X1 S_9_Rq3_reg_0_ ( .D(S_9_q3[0]), .CK(CLK), .Q(S_9_Rq3[0]), .QN() );
  DFF_X1 S_9_Rq3_reg_1_ ( .D(S_9_q3[1]), .CK(CLK), .Q(S_9_Rq3[1]), .QN() );
  DFF_X1 S_9_Rq3_reg_2_ ( .D(S_9_q3[2]), .CK(CLK), .Q(S_9_Rq3[2]), .QN() );
  DFF_X1 S_9_Rq3_reg_3_ ( .D(S_9_q3[3]), .CK(CLK), .Q(S_9_Rq3[3]), .QN() );
  DFF_X1 S_9_Rq2_reg_0_ ( .D(S_9_q2[0]), .CK(CLK), .Q(S_9_Rq2[0]), .QN() );
  DFF_X1 S_9_Rq2_reg_1_ ( .D(S_9_q2[1]), .CK(CLK), .Q(S_9_Rq2[1]), .QN() );
  DFF_X1 S_9_Rq2_reg_2_ ( .D(S_9_q2[2]), .CK(CLK), .Q(S_9_Rq2[2]), .QN() );
  DFF_X1 S_9_Rq2_reg_3_ ( .D(S_9_q2[3]), .CK(CLK), .Q(S_9_Rq2[3]), .QN() );
  DFF_X1 S_9_Rq1_reg_0_ ( .D(S_9_q1[0]), .CK(CLK), .Q(S_9_Rq1[0]), .QN() );
  DFF_X1 S_9_Rq1_reg_1_ ( .D(S_9_q1[1]), .CK(CLK), .Q(S_9_Rq1[1]), .QN() );
  DFF_X1 S_9_Rq1_reg_2_ ( .D(S_9_q1[2]), .CK(CLK), .Q(S_9_Rq1[2]), .QN() );
  DFF_X1 S_9_Rq1_reg_3_ ( .D(S_9_q1[3]), .CK(CLK), .Q(S_9_Rq1[3]), .QN() );
  INV_X1 S_9_InputAffine_U4 ( .A(SUB_IN1[36]), .ZN(S_9_F_in1[0]) );
  INV_X1 S_9_InputAffine_U3 ( .A(SUB_IN1[38]), .ZN(S_9_F_in1[3]) );
  INV_X1 S_9_InputAffine_U2 ( .A(SUB_IN1[39]), .ZN(S_9_F_in1[1]) );
  INV_X1 S_9_InputAffine_U1 ( .A(SUB_IN1[37]), .ZN(S_9_F_in1[2]) );
  XNOR2_X1 S_9_F_U18 ( .A(S_9_F_n12), .B(FRESH[75]), .ZN(S_9_q3[3]) );
  XNOR2_X1 S_9_F_U17 ( .A(FRESH[74]), .B(S_9_F_q3[3]), .ZN(S_9_F_n12) );
  XNOR2_X1 S_9_F_U16 ( .A(S_9_F_n11), .B(FRESH[73]), .ZN(S_9_q3[2]) );
  XNOR2_X1 S_9_F_U15 ( .A(FRESH[72]), .B(S_9_F_q3[2]), .ZN(S_9_F_n11) );
  XOR2_X1 S_9_F_U14 ( .A(FRESH[75]), .B(S_9_F_q2[3]), .Z(S_9_q2[3]) );
  XOR2_X1 S_9_F_U13 ( .A(FRESH[73]), .B(S_9_F_q2[2]), .Z(S_9_q2[2]) );
  XOR2_X1 S_9_F_U12 ( .A(FRESH[74]), .B(S_9_F_q1[3]), .Z(S_9_q1[3]) );
  XOR2_X1 S_9_F_U11 ( .A(FRESH[72]), .B(S_9_F_q1[2]), .Z(S_9_q1[2]) );
  XNOR2_X1 S_9_F_U10 ( .A(S_9_F_n10), .B(FRESH[77]), .ZN(S_9_F_N5) );
  XNOR2_X1 S_9_F_U9 ( .A(S_9_F_in3[3]), .B(FRESH[76]), .ZN(S_9_F_n10) );
  XOR2_X1 S_9_F_U8 ( .A(FRESH[77]), .B(S_9_F_in2[3]), .Z(S_9_F_N4) );
  XOR2_X1 S_9_F_U7 ( .A(FRESH[76]), .B(S_9_F_in1[3]), .Z(S_9_F_N3) );
  XNOR2_X1 S_9_F_U6 ( .A(S_9_F_n9), .B(FRESH[79]), .ZN(S_9_F_N2) );
  XNOR2_X1 S_9_F_U5 ( .A(S_9_F_in3[2]), .B(FRESH[78]), .ZN(S_9_F_n9) );
  XOR2_X1 S_9_F_U4 ( .A(FRESH[79]), .B(S_9_F_in2[2]), .Z(S_9_F_N1) );
  XOR2_X1 S_9_F_U3 ( .A(FRESH[78]), .B(S_9_F_in1[2]), .Z(S_9_F_N0) );
  DFF_X1 S_9_F_CF_Reg_reg_0_ ( .D(S_9_F_CF_Out[0]), .CK(CLK), .Q(
        S_9_F_CF_Reg[0]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_1_ ( .D(S_9_F_CF_Out[1]), .CK(CLK), .Q(
        S_9_F_CF_Reg[1]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_2_ ( .D(S_9_F_CF_Out[2]), .CK(CLK), .Q(
        S_9_F_CF_Reg[2]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_3_ ( .D(S_9_F_CF_Out[3]), .CK(CLK), .Q(
        S_9_F_CF_Reg[3]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_4_ ( .D(S_9_F_CF_Out[4]), .CK(CLK), .Q(
        S_9_F_CF_Reg[4]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_5_ ( .D(S_9_F_CF_Out[5]), .CK(CLK), .Q(
        S_9_F_CF_Reg[5]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_6_ ( .D(S_9_F_CF_Out[6]), .CK(CLK), .Q(
        S_9_F_CF_Reg[6]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_7_ ( .D(S_9_F_CF_Out[7]), .CK(CLK), .Q(
        S_9_F_CF_Reg[7]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_8_ ( .D(S_9_F_CF_Out[8]), .CK(CLK), .Q(
        S_9_F_CF_Reg[8]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_9_ ( .D(S_9_F_CF_Out[9]), .CK(CLK), .Q(
        S_9_F_CF_Reg[9]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_10_ ( .D(S_9_F_CF_Out[10]), .CK(CLK), .Q(
        S_9_F_CF_Reg[10]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_11_ ( .D(S_9_F_CF_Out[11]), .CK(CLK), .Q(
        S_9_F_CF_Reg[11]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_12_ ( .D(S_9_F_CF_Out[12]), .CK(CLK), .Q(
        S_9_F_CF_Reg[12]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_13_ ( .D(S_9_F_CF_Out[13]), .CK(CLK), .Q(
        S_9_F_CF_Reg[13]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_14_ ( .D(S_9_F_CF_Out[14]), .CK(CLK), .Q(
        S_9_F_CF_Reg[14]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_15_ ( .D(S_9_F_CF_Out[15]), .CK(CLK), .Q(
        S_9_F_CF_Reg[15]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_16_ ( .D(S_9_F_CF_Out[16]), .CK(CLK), .Q(
        S_9_F_CF_Reg[16]), .QN() );
  DFF_X1 S_9_F_CF_Reg_reg_17_ ( .D(S_9_F_CF_Out[17]), .CK(CLK), .Q(
        S_9_F_CF_Reg[17]), .QN() );
  DFF_X1 S_9_F_out2_reg_0_ ( .D(S_9_F_N4), .CK(CLK), .Q(S_9_q2[0]), .QN() );
  DFF_X1 S_9_F_out2_reg_1_ ( .D(S_9_F_N1), .CK(CLK), .Q(S_9_q2[1]), .QN() );
  DFF_X1 S_9_F_out3_reg_0_ ( .D(S_9_F_N5), .CK(CLK), .Q(S_9_q3[0]), .QN() );
  DFF_X1 S_9_F_out3_reg_1_ ( .D(S_9_F_N2), .CK(CLK), .Q(S_9_q3[1]), .QN() );
  DFF_X1 S_9_F_out1_reg_0_ ( .D(S_9_F_N3), .CK(CLK), .Q(S_9_q1[0]), .QN() );
  DFF_X1 S_9_F_out1_reg_1_ ( .D(S_9_F_N0), .CK(CLK), .Q(S_9_q1[1]), .QN() );
  NOR2_X1 S_9_F_Inst_0__CF_Inst_U2 ( .A1(S_9_F_in1[2]), .A2(
        S_9_F_Inst_0__CF_Inst_n3), .ZN(S_9_F_CF_Out[0]) );
  INV_X1 S_9_F_Inst_0__CF_Inst_U1 ( .A(S_9_F_in1[3]), .ZN(
        S_9_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_9_F_Inst_1__CF_Inst_U2 ( .A(S_9_F_Inst_1__CF_Inst_n3), .B(
        S_9_F_in1[1]), .ZN(S_9_F_CF_Out[1]) );
  NAND2_X1 S_9_F_Inst_1__CF_Inst_U1 ( .A1(S_9_F_in2[2]), .A2(S_9_F_in1[3]), 
        .ZN(S_9_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_9_F_Inst_2__CF_Inst_U1 ( .A1(S_9_F_in1[3]), .A2(S_9_F_in3[2]), .ZN(
        S_9_F_CF_Out[2]) );
  NOR2_X1 S_9_F_Inst_3__CF_Inst_U2 ( .A1(S_9_F_in2[3]), .A2(
        S_9_F_Inst_3__CF_Inst_n3), .ZN(S_9_F_CF_Out[3]) );
  INV_X1 S_9_F_Inst_3__CF_Inst_U1 ( .A(S_9_F_in1[2]), .ZN(
        S_9_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_9_F_Inst_4__CF_Inst_U2 ( .A(S_9_F_Inst_4__CF_Inst_n3), .B(
        S_9_F_in2[1]), .ZN(S_9_F_CF_Out[4]) );
  NAND2_X1 S_9_F_Inst_4__CF_Inst_U1 ( .A1(S_9_F_in2[2]), .A2(S_9_F_in2[3]), 
        .ZN(S_9_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_9_F_Inst_5__CF_Inst_U1 ( .A1(S_9_F_in3[2]), .A2(S_9_F_in2[3]), 
        .ZN(S_9_F_CF_Out[5]) );
  XNOR2_X1 S_9_F_Inst_6__CF_Inst_U2 ( .A(S_9_F_Inst_6__CF_Inst_n7), .B(
        S_9_F_in3[1]), .ZN(S_9_F_CF_Out[6]) );
  NOR2_X1 S_9_F_Inst_6__CF_Inst_U1 ( .A1(S_9_F_in1[2]), .A2(S_9_F_in3[3]), 
        .ZN(S_9_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_9_F_Inst_7__CF_Inst_U1 ( .A1(S_9_F_in2[2]), .A2(S_9_F_in3[3]), 
        .ZN(S_9_F_CF_Out[7]) );
  OR2_X1 S_9_F_Inst_8__CF_Inst_U1 ( .A1(S_9_F_in3[3]), .A2(S_9_F_in3[2]), .ZN(
        S_9_F_CF_Out[8]) );
  NOR2_X1 S_9_F_Inst_9__CF_Inst_U2 ( .A1(S_9_F_in1[3]), .A2(
        S_9_F_Inst_9__CF_Inst_n3), .ZN(S_9_F_CF_Out[9]) );
  INV_X1 S_9_F_Inst_9__CF_Inst_U1 ( .A(S_9_F_in1[1]), .ZN(
        S_9_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_9_F_Inst_10__CF_Inst_U1 ( .A1(S_9_F_in2[1]), .A2(S_9_F_in1[3]), 
        .ZN(S_9_F_CF_Out[10]) );
  XNOR2_X1 S_9_F_Inst_11__CF_Inst_U2 ( .A(S_9_F_Inst_11__CF_Inst_n3), .B(
        S_9_F_in1[0]), .ZN(S_9_F_CF_Out[11]) );
  NAND2_X1 S_9_F_Inst_11__CF_Inst_U1 ( .A1(S_9_F_in3[1]), .A2(S_9_F_in1[3]), 
        .ZN(S_9_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_9_F_Inst_12__CF_Inst_U2 ( .A(S_9_F_Inst_12__CF_Inst_n3), .B(
        S_9_F_in2[0]), .ZN(S_9_F_CF_Out[12]) );
  NAND2_X1 S_9_F_Inst_12__CF_Inst_U1 ( .A1(S_9_F_in1[1]), .A2(S_9_F_in2[3]), 
        .ZN(S_9_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_9_F_Inst_13__CF_Inst_U2 ( .A1(S_9_F_in2[3]), .A2(
        S_9_F_Inst_13__CF_Inst_n3), .ZN(S_9_F_CF_Out[13]) );
  INV_X1 S_9_F_Inst_13__CF_Inst_U1 ( .A(S_9_F_in2[1]), .ZN(
        S_9_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_9_F_Inst_14__CF_Inst_U1 ( .A1(S_9_F_in3[1]), .A2(S_9_F_in2[3]), 
        .ZN(S_9_F_CF_Out[14]) );
  XNOR2_X1 S_9_F_Inst_15__CF_Inst_U2 ( .A(S_9_F_Inst_15__CF_Inst_n7), .B(
        S_9_F_in3[0]), .ZN(S_9_F_CF_Out[15]) );
  NOR2_X1 S_9_F_Inst_15__CF_Inst_U1 ( .A1(S_9_F_in1[1]), .A2(S_9_F_in3[3]), 
        .ZN(S_9_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_9_F_Inst_16__CF_Inst_U2 ( .A1(S_9_F_in3[3]), .A2(
        S_9_F_Inst_16__CF_Inst_n3), .ZN(S_9_F_CF_Out[16]) );
  INV_X1 S_9_F_Inst_16__CF_Inst_U1 ( .A(S_9_F_in2[1]), .ZN(
        S_9_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_9_F_Inst_17__CF_Inst_U2 ( .A1(S_9_F_in3[1]), .A2(
        S_9_F_Inst_17__CF_Inst_n3), .ZN(S_9_F_CF_Out[17]) );
  INV_X1 S_9_F_Inst_17__CF_Inst_U1 ( .A(S_9_F_in3[3]), .ZN(
        S_9_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_9_F_InstXOR_0__Compression1_U2 ( .A(
        S_9_F_InstXOR_0__Compression1_n3), .B(S_9_F_CF_Reg[2]), .ZN(
        S_9_F_q1[2]) );
  XNOR2_X1 S_9_F_InstXOR_0__Compression1_U1 ( .A(S_9_F_CF_Reg[0]), .B(
        S_9_F_CF_Reg[1]), .ZN(S_9_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_9_F_InstXOR_0__Compression2_U2 ( .A(
        S_9_F_InstXOR_0__Compression2_n3), .B(S_9_F_CF_Reg[5]), .ZN(
        S_9_F_q2[2]) );
  XNOR2_X1 S_9_F_InstXOR_0__Compression2_U1 ( .A(S_9_F_CF_Reg[3]), .B(
        S_9_F_CF_Reg[4]), .ZN(S_9_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_9_F_InstXOR_0__Compression3_U2 ( .A(
        S_9_F_InstXOR_0__Compression3_n3), .B(S_9_F_CF_Reg[8]), .ZN(
        S_9_F_q3[2]) );
  XNOR2_X1 S_9_F_InstXOR_0__Compression3_U1 ( .A(S_9_F_CF_Reg[6]), .B(
        S_9_F_CF_Reg[7]), .ZN(S_9_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_9_F_InstXOR_1__Compression1_U2 ( .A(
        S_9_F_InstXOR_1__Compression1_n3), .B(S_9_F_CF_Reg[11]), .ZN(
        S_9_F_q1[3]) );
  XNOR2_X1 S_9_F_InstXOR_1__Compression1_U1 ( .A(S_9_F_CF_Reg[9]), .B(
        S_9_F_CF_Reg[10]), .ZN(S_9_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_9_F_InstXOR_1__Compression2_U2 ( .A(
        S_9_F_InstXOR_1__Compression2_n3), .B(S_9_F_CF_Reg[14]), .ZN(
        S_9_F_q2[3]) );
  XNOR2_X1 S_9_F_InstXOR_1__Compression2_U1 ( .A(S_9_F_CF_Reg[12]), .B(
        S_9_F_CF_Reg[13]), .ZN(S_9_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_9_F_InstXOR_1__Compression3_U2 ( .A(
        S_9_F_InstXOR_1__Compression3_n3), .B(S_9_F_CF_Reg[17]), .ZN(
        S_9_F_q3[3]) );
  XNOR2_X1 S_9_F_InstXOR_1__Compression3_U1 ( .A(S_9_F_CF_Reg[15]), .B(
        S_9_F_CF_Reg[16]), .ZN(S_9_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_9_G_CF_Reg_reg_0_ ( .D(S_9_G_CF_Out[0]), .CK(CLK), .Q(
        S_9_G_CF_Reg[0]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_1_ ( .D(S_9_G_CF_Out[1]), .CK(CLK), .Q(
        S_9_G_CF_Reg[1]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_2_ ( .D(S_9_G_CF_Out[2]), .CK(CLK), .Q(
        S_9_G_CF_Reg[2]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_3_ ( .D(S_9_G_CF_Out[3]), .CK(CLK), .Q(
        S_9_G_CF_Reg[3]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_4_ ( .D(S_9_G_CF_Out[4]), .CK(CLK), .Q(
        S_9_G_CF_Reg[4]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_5_ ( .D(S_9_G_CF_Out[5]), .CK(CLK), .Q(
        S_9_G_CF_Reg[5]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_6_ ( .D(S_9_G_CF_Out[6]), .CK(CLK), .Q(
        S_9_G_CF_Reg[6]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_7_ ( .D(S_9_G_CF_Out[7]), .CK(CLK), .Q(
        S_9_G_CF_Reg[7]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_8_ ( .D(S_9_G_CF_Out[8]), .CK(CLK), .Q(
        S_9_G_CF_Reg[8]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_9_ ( .D(S_9_G_CF_Out[9]), .CK(CLK), .Q(
        S_9_G_CF_Reg[9]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_10_ ( .D(S_9_G_CF_Out[10]), .CK(CLK), .Q(
        S_9_G_CF_Reg[10]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_11_ ( .D(S_9_G_CF_Out[11]), .CK(CLK), .Q(
        S_9_G_CF_Reg[11]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_12_ ( .D(S_9_G_CF_Out[12]), .CK(CLK), .Q(
        S_9_G_CF_Reg[12]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_13_ ( .D(S_9_G_CF_Out[13]), .CK(CLK), .Q(
        S_9_G_CF_Reg[13]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_14_ ( .D(S_9_G_CF_Out[14]), .CK(CLK), .Q(
        S_9_G_CF_Reg[14]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_15_ ( .D(S_9_G_CF_Out[15]), .CK(CLK), .Q(
        S_9_G_CF_Reg[15]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_16_ ( .D(S_9_G_CF_Out[16]), .CK(CLK), .Q(
        S_9_G_CF_Reg[16]), .QN() );
  DFF_X1 S_9_G_CF_Reg_reg_17_ ( .D(S_9_G_CF_Out[17]), .CK(CLK), .Q(
        S_9_G_CF_Reg[17]), .QN() );
  DFF_X1 S_9_G_out1_reg_2_ ( .D(S_9_Rq1[2]), .CK(CLK), .Q(S_9_G_out1[2]), 
        .QN() );
  DFF_X1 S_9_G_out1_reg_3_ ( .D(S_9_Rq1[3]), .CK(CLK), .Q(S_9_G_out1[3]), 
        .QN() );
  DFF_X1 S_9_G_out2_reg_2_ ( .D(S_9_Rq2[2]), .CK(CLK), .Q(SUB_OUT2[38]), .QN()
         );
  DFF_X1 S_9_G_out2_reg_3_ ( .D(S_9_Rq2[3]), .CK(CLK), .Q(SUB_OUT2[39]), .QN()
         );
  DFF_X1 S_9_G_out3_reg_2_ ( .D(S_9_Rq3[2]), .CK(CLK), .Q(SUB_OUT3[38]), .QN()
         );
  DFF_X1 S_9_G_out3_reg_3_ ( .D(S_9_Rq3[3]), .CK(CLK), .Q(SUB_OUT3[39]), .QN()
         );
  AND2_X1 S_9_G_Inst_0__CF_Inst_U1 ( .A1(S_9_Rq1[1]), .A2(S_9_Rq1[3]), .ZN(
        S_9_G_CF_Out[0]) );
  NOR2_X1 S_9_G_Inst_1__CF_Inst_U2 ( .A1(S_9_Rq1[3]), .A2(
        S_9_G_Inst_1__CF_Inst_n3), .ZN(S_9_G_CF_Out[1]) );
  INV_X1 S_9_G_Inst_1__CF_Inst_U1 ( .A(S_9_Rq2[1]), .ZN(
        S_9_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_9_G_Inst_2__CF_Inst_U2 ( .A(S_9_G_Inst_2__CF_Inst_n3), .B(
        S_9_Rq2[0]), .ZN(S_9_G_CF_Out[2]) );
  NAND2_X1 S_9_G_Inst_2__CF_Inst_U1 ( .A1(S_9_Rq1[1]), .A2(S_9_Rq2[3]), .ZN(
        S_9_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_9_G_Inst_3__CF_Inst_U3 ( .A(S_9_Rq1[0]), .B(
        S_9_G_Inst_3__CF_Inst_n6), .ZN(S_9_G_CF_Out[3]) );
  NAND2_X1 S_9_G_Inst_3__CF_Inst_U2 ( .A1(S_9_Rq3[1]), .A2(
        S_9_G_Inst_3__CF_Inst_n5), .ZN(S_9_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_9_G_Inst_3__CF_Inst_U1 ( .A(S_9_Rq1[3]), .ZN(
        S_9_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_9_G_Inst_4__CF_Inst_U1 ( .A1(S_9_Rq2[1]), .A2(S_9_Rq2[3]), .ZN(
        S_9_G_CF_Out[4]) );
  OR2_X1 S_9_G_Inst_5__CF_Inst_U1 ( .A1(S_9_Rq3[3]), .A2(S_9_Rq2[1]), .ZN(
        S_9_G_CF_Out[5]) );
  AND2_X1 S_9_G_Inst_6__CF_Inst_U1 ( .A1(S_9_Rq3[1]), .A2(S_9_Rq2[3]), .ZN(
        S_9_G_CF_Out[6]) );
  XNOR2_X1 S_9_G_Inst_7__CF_Inst_U2 ( .A(S_9_G_Inst_7__CF_Inst_n3), .B(
        S_9_Rq3[0]), .ZN(S_9_G_CF_Out[7]) );
  NAND2_X1 S_9_G_Inst_7__CF_Inst_U1 ( .A1(S_9_Rq1[1]), .A2(S_9_Rq3[3]), .ZN(
        S_9_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_9_G_Inst_8__CF_Inst_U1 ( .A1(S_9_Rq3[3]), .A2(S_9_Rq3[1]), .ZN(
        S_9_G_CF_Out[8]) );
  NOR2_X1 S_9_G_Inst_9__CF_Inst_U2 ( .A1(S_9_Rq1[3]), .A2(
        S_9_G_Inst_9__CF_Inst_n3), .ZN(S_9_G_CF_Out[9]) );
  INV_X1 S_9_G_Inst_9__CF_Inst_U1 ( .A(S_9_Rq1[2]), .ZN(
        S_9_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_9_G_Inst_10__CF_Inst_U2 ( .A1(S_9_Rq2[2]), .A2(
        S_9_G_Inst_10__CF_Inst_n3), .ZN(S_9_G_CF_Out[10]) );
  INV_X1 S_9_G_Inst_10__CF_Inst_U1 ( .A(S_9_Rq1[3]), .ZN(
        S_9_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_9_G_Inst_11__CF_Inst_U3 ( .A(S_9_Rq1[1]), .B(
        S_9_G_Inst_11__CF_Inst_n6), .ZN(S_9_G_CF_Out[11]) );
  NAND2_X1 S_9_G_Inst_11__CF_Inst_U2 ( .A1(S_9_Rq1[3]), .A2(
        S_9_G_Inst_11__CF_Inst_n5), .ZN(S_9_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_9_G_Inst_11__CF_Inst_U1 ( .A(S_9_Rq3[2]), .ZN(
        S_9_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_9_G_Inst_12__CF_Inst_U2 ( .A1(S_9_Rq2[3]), .A2(
        S_9_G_Inst_12__CF_Inst_n3), .ZN(S_9_G_CF_Out[12]) );
  INV_X1 S_9_G_Inst_12__CF_Inst_U1 ( .A(S_9_Rq1[2]), .ZN(
        S_9_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_9_G_Inst_13__CF_Inst_U1 ( .A1(S_9_Rq2[2]), .A2(S_9_Rq2[3]), .ZN(
        S_9_G_CF_Out[13]) );
  XNOR2_X1 S_9_G_Inst_14__CF_Inst_U3 ( .A(S_9_Rq2[1]), .B(
        S_9_G_Inst_14__CF_Inst_n6), .ZN(S_9_G_CF_Out[14]) );
  NAND2_X1 S_9_G_Inst_14__CF_Inst_U2 ( .A1(S_9_Rq3[2]), .A2(
        S_9_G_Inst_14__CF_Inst_n5), .ZN(S_9_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_9_G_Inst_14__CF_Inst_U1 ( .A(S_9_Rq2[3]), .ZN(
        S_9_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_9_G_Inst_15__CF_Inst_U2 ( .A(S_9_G_Inst_15__CF_Inst_n3), .B(
        S_9_Rq3[1]), .ZN(S_9_G_CF_Out[15]) );
  NAND2_X1 S_9_G_Inst_15__CF_Inst_U1 ( .A1(S_9_Rq1[2]), .A2(S_9_Rq3[3]), .ZN(
        S_9_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_9_G_Inst_16__CF_Inst_U1 ( .A1(S_9_Rq2[2]), .A2(S_9_Rq3[3]), .ZN(
        S_9_G_CF_Out[16]) );
  NOR2_X1 S_9_G_Inst_17__CF_Inst_U2 ( .A1(S_9_Rq3[3]), .A2(
        S_9_G_Inst_17__CF_Inst_n3), .ZN(S_9_G_CF_Out[17]) );
  INV_X1 S_9_G_Inst_17__CF_Inst_U1 ( .A(S_9_Rq3[2]), .ZN(
        S_9_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_9_G_InstXOR_0__Compression1_U2 ( .A(
        S_9_G_InstXOR_0__Compression1_n3), .B(S_9_G_CF_Reg[2]), .ZN(
        S_9_G_out1[0]) );
  XNOR2_X1 S_9_G_InstXOR_0__Compression1_U1 ( .A(S_9_G_CF_Reg[0]), .B(
        S_9_G_CF_Reg[1]), .ZN(S_9_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_9_G_InstXOR_0__Compression2_U2 ( .A(
        S_9_G_InstXOR_0__Compression2_n3), .B(S_9_G_CF_Reg[5]), .ZN(
        SUB_OUT2[37]) );
  XNOR2_X1 S_9_G_InstXOR_0__Compression2_U1 ( .A(S_9_G_CF_Reg[3]), .B(
        S_9_G_CF_Reg[4]), .ZN(S_9_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_9_G_InstXOR_0__Compression3_U2 ( .A(
        S_9_G_InstXOR_0__Compression3_n3), .B(S_9_G_CF_Reg[8]), .ZN(
        SUB_OUT3[37]) );
  XNOR2_X1 S_9_G_InstXOR_0__Compression3_U1 ( .A(S_9_G_CF_Reg[6]), .B(
        S_9_G_CF_Reg[7]), .ZN(S_9_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_9_G_InstXOR_1__Compression1_U2 ( .A(
        S_9_G_InstXOR_1__Compression1_n3), .B(S_9_G_CF_Reg[11]), .ZN(
        S_9_G_out1[1]) );
  XNOR2_X1 S_9_G_InstXOR_1__Compression1_U1 ( .A(S_9_G_CF_Reg[9]), .B(
        S_9_G_CF_Reg[10]), .ZN(S_9_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_9_G_InstXOR_1__Compression2_U2 ( .A(
        S_9_G_InstXOR_1__Compression2_n3), .B(S_9_G_CF_Reg[14]), .ZN(
        SUB_OUT2[36]) );
  XNOR2_X1 S_9_G_InstXOR_1__Compression2_U1 ( .A(S_9_G_CF_Reg[12]), .B(
        S_9_G_CF_Reg[13]), .ZN(S_9_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_9_G_InstXOR_1__Compression3_U2 ( .A(
        S_9_G_InstXOR_1__Compression3_n3), .B(S_9_G_CF_Reg[17]), .ZN(
        SUB_OUT3[36]) );
  XNOR2_X1 S_9_G_InstXOR_1__Compression3_U1 ( .A(S_9_G_CF_Reg[15]), .B(
        S_9_G_CF_Reg[16]), .ZN(S_9_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_9_OutputAffine_U4 ( .A(S_9_G_out1[3]), .ZN(SUB_OUT1[39]) );
  INV_X1 S_9_OutputAffine_U3 ( .A(S_9_G_out1[2]), .ZN(SUB_OUT1[38]) );
  INV_X1 S_9_OutputAffine_U2 ( .A(S_9_G_out1[1]), .ZN(SUB_OUT1[36]) );
  INV_X1 S_9_OutputAffine_U1 ( .A(S_9_G_out1[0]), .ZN(SUB_OUT1[37]) );
  DFF_X1 S_10_Rq3_reg_0_ ( .D(S_10_q3[0]), .CK(CLK), .Q(S_10_Rq3[0]), .QN() );
  DFF_X1 S_10_Rq3_reg_1_ ( .D(S_10_q3[1]), .CK(CLK), .Q(S_10_Rq3[1]), .QN() );
  DFF_X1 S_10_Rq3_reg_2_ ( .D(S_10_q3[2]), .CK(CLK), .Q(S_10_Rq3[2]), .QN() );
  DFF_X1 S_10_Rq3_reg_3_ ( .D(S_10_q3[3]), .CK(CLK), .Q(S_10_Rq3[3]), .QN() );
  DFF_X1 S_10_Rq2_reg_0_ ( .D(S_10_q2[0]), .CK(CLK), .Q(S_10_Rq2[0]), .QN() );
  DFF_X1 S_10_Rq2_reg_1_ ( .D(S_10_q2[1]), .CK(CLK), .Q(S_10_Rq2[1]), .QN() );
  DFF_X1 S_10_Rq2_reg_2_ ( .D(S_10_q2[2]), .CK(CLK), .Q(S_10_Rq2[2]), .QN() );
  DFF_X1 S_10_Rq2_reg_3_ ( .D(S_10_q2[3]), .CK(CLK), .Q(S_10_Rq2[3]), .QN() );
  DFF_X1 S_10_Rq1_reg_0_ ( .D(S_10_q1[0]), .CK(CLK), .Q(S_10_Rq1[0]), .QN() );
  DFF_X1 S_10_Rq1_reg_1_ ( .D(S_10_q1[1]), .CK(CLK), .Q(S_10_Rq1[1]), .QN() );
  DFF_X1 S_10_Rq1_reg_2_ ( .D(S_10_q1[2]), .CK(CLK), .Q(S_10_Rq1[2]), .QN() );
  DFF_X1 S_10_Rq1_reg_3_ ( .D(S_10_q1[3]), .CK(CLK), .Q(S_10_Rq1[3]), .QN() );
  INV_X1 S_10_InputAffine_U4 ( .A(SUB_IN1[40]), .ZN(S_10_F_in1[0]) );
  INV_X1 S_10_InputAffine_U3 ( .A(SUB_IN1[42]), .ZN(S_10_F_in1[3]) );
  INV_X1 S_10_InputAffine_U2 ( .A(SUB_IN1[43]), .ZN(S_10_F_in1[1]) );
  INV_X1 S_10_InputAffine_U1 ( .A(SUB_IN1[41]), .ZN(S_10_F_in1[2]) );
  XNOR2_X1 S_10_F_U18 ( .A(S_10_F_n12), .B(FRESH[83]), .ZN(S_10_q3[3]) );
  XNOR2_X1 S_10_F_U17 ( .A(FRESH[82]), .B(S_10_F_q3[3]), .ZN(S_10_F_n12) );
  XNOR2_X1 S_10_F_U16 ( .A(S_10_F_n11), .B(FRESH[81]), .ZN(S_10_q3[2]) );
  XNOR2_X1 S_10_F_U15 ( .A(FRESH[80]), .B(S_10_F_q3[2]), .ZN(S_10_F_n11) );
  XOR2_X1 S_10_F_U14 ( .A(FRESH[83]), .B(S_10_F_q2[3]), .Z(S_10_q2[3]) );
  XOR2_X1 S_10_F_U13 ( .A(FRESH[81]), .B(S_10_F_q2[2]), .Z(S_10_q2[2]) );
  XOR2_X1 S_10_F_U12 ( .A(FRESH[82]), .B(S_10_F_q1[3]), .Z(S_10_q1[3]) );
  XOR2_X1 S_10_F_U11 ( .A(FRESH[80]), .B(S_10_F_q1[2]), .Z(S_10_q1[2]) );
  XNOR2_X1 S_10_F_U10 ( .A(S_10_F_n10), .B(FRESH[85]), .ZN(S_10_F_N5) );
  XNOR2_X1 S_10_F_U9 ( .A(S_10_F_in3[3]), .B(FRESH[84]), .ZN(S_10_F_n10) );
  XOR2_X1 S_10_F_U8 ( .A(FRESH[85]), .B(S_10_F_in2[3]), .Z(S_10_F_N4) );
  XOR2_X1 S_10_F_U7 ( .A(FRESH[84]), .B(S_10_F_in1[3]), .Z(S_10_F_N3) );
  XNOR2_X1 S_10_F_U6 ( .A(S_10_F_n9), .B(FRESH[87]), .ZN(S_10_F_N2) );
  XNOR2_X1 S_10_F_U5 ( .A(S_10_F_in3[2]), .B(FRESH[86]), .ZN(S_10_F_n9) );
  XOR2_X1 S_10_F_U4 ( .A(FRESH[87]), .B(S_10_F_in2[2]), .Z(S_10_F_N1) );
  XOR2_X1 S_10_F_U3 ( .A(FRESH[86]), .B(S_10_F_in1[2]), .Z(S_10_F_N0) );
  DFF_X1 S_10_F_CF_Reg_reg_0_ ( .D(S_10_F_CF_Out[0]), .CK(CLK), .Q(
        S_10_F_CF_Reg[0]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_1_ ( .D(S_10_F_CF_Out[1]), .CK(CLK), .Q(
        S_10_F_CF_Reg[1]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_2_ ( .D(S_10_F_CF_Out[2]), .CK(CLK), .Q(
        S_10_F_CF_Reg[2]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_3_ ( .D(S_10_F_CF_Out[3]), .CK(CLK), .Q(
        S_10_F_CF_Reg[3]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_4_ ( .D(S_10_F_CF_Out[4]), .CK(CLK), .Q(
        S_10_F_CF_Reg[4]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_5_ ( .D(S_10_F_CF_Out[5]), .CK(CLK), .Q(
        S_10_F_CF_Reg[5]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_6_ ( .D(S_10_F_CF_Out[6]), .CK(CLK), .Q(
        S_10_F_CF_Reg[6]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_7_ ( .D(S_10_F_CF_Out[7]), .CK(CLK), .Q(
        S_10_F_CF_Reg[7]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_8_ ( .D(S_10_F_CF_Out[8]), .CK(CLK), .Q(
        S_10_F_CF_Reg[8]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_9_ ( .D(S_10_F_CF_Out[9]), .CK(CLK), .Q(
        S_10_F_CF_Reg[9]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_10_ ( .D(S_10_F_CF_Out[10]), .CK(CLK), .Q(
        S_10_F_CF_Reg[10]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_11_ ( .D(S_10_F_CF_Out[11]), .CK(CLK), .Q(
        S_10_F_CF_Reg[11]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_12_ ( .D(S_10_F_CF_Out[12]), .CK(CLK), .Q(
        S_10_F_CF_Reg[12]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_13_ ( .D(S_10_F_CF_Out[13]), .CK(CLK), .Q(
        S_10_F_CF_Reg[13]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_14_ ( .D(S_10_F_CF_Out[14]), .CK(CLK), .Q(
        S_10_F_CF_Reg[14]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_15_ ( .D(S_10_F_CF_Out[15]), .CK(CLK), .Q(
        S_10_F_CF_Reg[15]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_16_ ( .D(S_10_F_CF_Out[16]), .CK(CLK), .Q(
        S_10_F_CF_Reg[16]), .QN() );
  DFF_X1 S_10_F_CF_Reg_reg_17_ ( .D(S_10_F_CF_Out[17]), .CK(CLK), .Q(
        S_10_F_CF_Reg[17]), .QN() );
  DFF_X1 S_10_F_out2_reg_0_ ( .D(S_10_F_N4), .CK(CLK), .Q(S_10_q2[0]), .QN()
         );
  DFF_X1 S_10_F_out2_reg_1_ ( .D(S_10_F_N1), .CK(CLK), .Q(S_10_q2[1]), .QN()
         );
  DFF_X1 S_10_F_out3_reg_0_ ( .D(S_10_F_N5), .CK(CLK), .Q(S_10_q3[0]), .QN()
         );
  DFF_X1 S_10_F_out3_reg_1_ ( .D(S_10_F_N2), .CK(CLK), .Q(S_10_q3[1]), .QN()
         );
  DFF_X1 S_10_F_out1_reg_0_ ( .D(S_10_F_N3), .CK(CLK), .Q(S_10_q1[0]), .QN()
         );
  DFF_X1 S_10_F_out1_reg_1_ ( .D(S_10_F_N0), .CK(CLK), .Q(S_10_q1[1]), .QN()
         );
  NOR2_X1 S_10_F_Inst_0__CF_Inst_U2 ( .A1(S_10_F_in1[2]), .A2(
        S_10_F_Inst_0__CF_Inst_n3), .ZN(S_10_F_CF_Out[0]) );
  INV_X1 S_10_F_Inst_0__CF_Inst_U1 ( .A(S_10_F_in1[3]), .ZN(
        S_10_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_10_F_Inst_1__CF_Inst_U2 ( .A(S_10_F_Inst_1__CF_Inst_n3), .B(
        S_10_F_in1[1]), .ZN(S_10_F_CF_Out[1]) );
  NAND2_X1 S_10_F_Inst_1__CF_Inst_U1 ( .A1(S_10_F_in2[2]), .A2(S_10_F_in1[3]), 
        .ZN(S_10_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_10_F_Inst_2__CF_Inst_U1 ( .A1(S_10_F_in1[3]), .A2(S_10_F_in3[2]), 
        .ZN(S_10_F_CF_Out[2]) );
  NOR2_X1 S_10_F_Inst_3__CF_Inst_U2 ( .A1(S_10_F_in2[3]), .A2(
        S_10_F_Inst_3__CF_Inst_n3), .ZN(S_10_F_CF_Out[3]) );
  INV_X1 S_10_F_Inst_3__CF_Inst_U1 ( .A(S_10_F_in1[2]), .ZN(
        S_10_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_10_F_Inst_4__CF_Inst_U2 ( .A(S_10_F_Inst_4__CF_Inst_n3), .B(
        S_10_F_in2[1]), .ZN(S_10_F_CF_Out[4]) );
  NAND2_X1 S_10_F_Inst_4__CF_Inst_U1 ( .A1(S_10_F_in2[2]), .A2(S_10_F_in2[3]), 
        .ZN(S_10_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_10_F_Inst_5__CF_Inst_U1 ( .A1(S_10_F_in3[2]), .A2(S_10_F_in2[3]), 
        .ZN(S_10_F_CF_Out[5]) );
  XNOR2_X1 S_10_F_Inst_6__CF_Inst_U2 ( .A(S_10_F_Inst_6__CF_Inst_n7), .B(
        S_10_F_in3[1]), .ZN(S_10_F_CF_Out[6]) );
  NOR2_X1 S_10_F_Inst_6__CF_Inst_U1 ( .A1(S_10_F_in1[2]), .A2(S_10_F_in3[3]), 
        .ZN(S_10_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_10_F_Inst_7__CF_Inst_U1 ( .A1(S_10_F_in2[2]), .A2(S_10_F_in3[3]), 
        .ZN(S_10_F_CF_Out[7]) );
  OR2_X1 S_10_F_Inst_8__CF_Inst_U1 ( .A1(S_10_F_in3[3]), .A2(S_10_F_in3[2]), 
        .ZN(S_10_F_CF_Out[8]) );
  NOR2_X1 S_10_F_Inst_9__CF_Inst_U2 ( .A1(S_10_F_in1[3]), .A2(
        S_10_F_Inst_9__CF_Inst_n3), .ZN(S_10_F_CF_Out[9]) );
  INV_X1 S_10_F_Inst_9__CF_Inst_U1 ( .A(S_10_F_in1[1]), .ZN(
        S_10_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_10_F_Inst_10__CF_Inst_U1 ( .A1(S_10_F_in2[1]), .A2(S_10_F_in1[3]), 
        .ZN(S_10_F_CF_Out[10]) );
  XNOR2_X1 S_10_F_Inst_11__CF_Inst_U2 ( .A(S_10_F_Inst_11__CF_Inst_n3), .B(
        S_10_F_in1[0]), .ZN(S_10_F_CF_Out[11]) );
  NAND2_X1 S_10_F_Inst_11__CF_Inst_U1 ( .A1(S_10_F_in3[1]), .A2(S_10_F_in1[3]), 
        .ZN(S_10_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_10_F_Inst_12__CF_Inst_U2 ( .A(S_10_F_Inst_12__CF_Inst_n3), .B(
        S_10_F_in2[0]), .ZN(S_10_F_CF_Out[12]) );
  NAND2_X1 S_10_F_Inst_12__CF_Inst_U1 ( .A1(S_10_F_in1[1]), .A2(S_10_F_in2[3]), 
        .ZN(S_10_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_10_F_Inst_13__CF_Inst_U2 ( .A1(S_10_F_in2[3]), .A2(
        S_10_F_Inst_13__CF_Inst_n3), .ZN(S_10_F_CF_Out[13]) );
  INV_X1 S_10_F_Inst_13__CF_Inst_U1 ( .A(S_10_F_in2[1]), .ZN(
        S_10_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_10_F_Inst_14__CF_Inst_U1 ( .A1(S_10_F_in3[1]), .A2(S_10_F_in2[3]), 
        .ZN(S_10_F_CF_Out[14]) );
  XNOR2_X1 S_10_F_Inst_15__CF_Inst_U2 ( .A(S_10_F_Inst_15__CF_Inst_n7), .B(
        S_10_F_in3[0]), .ZN(S_10_F_CF_Out[15]) );
  NOR2_X1 S_10_F_Inst_15__CF_Inst_U1 ( .A1(S_10_F_in1[1]), .A2(S_10_F_in3[3]), 
        .ZN(S_10_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_10_F_Inst_16__CF_Inst_U2 ( .A1(S_10_F_in3[3]), .A2(
        S_10_F_Inst_16__CF_Inst_n3), .ZN(S_10_F_CF_Out[16]) );
  INV_X1 S_10_F_Inst_16__CF_Inst_U1 ( .A(S_10_F_in2[1]), .ZN(
        S_10_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_10_F_Inst_17__CF_Inst_U2 ( .A1(S_10_F_in3[1]), .A2(
        S_10_F_Inst_17__CF_Inst_n3), .ZN(S_10_F_CF_Out[17]) );
  INV_X1 S_10_F_Inst_17__CF_Inst_U1 ( .A(S_10_F_in3[3]), .ZN(
        S_10_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_10_F_InstXOR_0__Compression1_U2 ( .A(
        S_10_F_InstXOR_0__Compression1_n3), .B(S_10_F_CF_Reg[2]), .ZN(
        S_10_F_q1[2]) );
  XNOR2_X1 S_10_F_InstXOR_0__Compression1_U1 ( .A(S_10_F_CF_Reg[0]), .B(
        S_10_F_CF_Reg[1]), .ZN(S_10_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_10_F_InstXOR_0__Compression2_U2 ( .A(
        S_10_F_InstXOR_0__Compression2_n3), .B(S_10_F_CF_Reg[5]), .ZN(
        S_10_F_q2[2]) );
  XNOR2_X1 S_10_F_InstXOR_0__Compression2_U1 ( .A(S_10_F_CF_Reg[3]), .B(
        S_10_F_CF_Reg[4]), .ZN(S_10_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_10_F_InstXOR_0__Compression3_U2 ( .A(
        S_10_F_InstXOR_0__Compression3_n3), .B(S_10_F_CF_Reg[8]), .ZN(
        S_10_F_q3[2]) );
  XNOR2_X1 S_10_F_InstXOR_0__Compression3_U1 ( .A(S_10_F_CF_Reg[6]), .B(
        S_10_F_CF_Reg[7]), .ZN(S_10_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_10_F_InstXOR_1__Compression1_U2 ( .A(
        S_10_F_InstXOR_1__Compression1_n3), .B(S_10_F_CF_Reg[11]), .ZN(
        S_10_F_q1[3]) );
  XNOR2_X1 S_10_F_InstXOR_1__Compression1_U1 ( .A(S_10_F_CF_Reg[9]), .B(
        S_10_F_CF_Reg[10]), .ZN(S_10_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_10_F_InstXOR_1__Compression2_U2 ( .A(
        S_10_F_InstXOR_1__Compression2_n3), .B(S_10_F_CF_Reg[14]), .ZN(
        S_10_F_q2[3]) );
  XNOR2_X1 S_10_F_InstXOR_1__Compression2_U1 ( .A(S_10_F_CF_Reg[12]), .B(
        S_10_F_CF_Reg[13]), .ZN(S_10_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_10_F_InstXOR_1__Compression3_U2 ( .A(
        S_10_F_InstXOR_1__Compression3_n3), .B(S_10_F_CF_Reg[17]), .ZN(
        S_10_F_q3[3]) );
  XNOR2_X1 S_10_F_InstXOR_1__Compression3_U1 ( .A(S_10_F_CF_Reg[15]), .B(
        S_10_F_CF_Reg[16]), .ZN(S_10_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_10_G_CF_Reg_reg_0_ ( .D(S_10_G_CF_Out[0]), .CK(CLK), .Q(
        S_10_G_CF_Reg[0]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_1_ ( .D(S_10_G_CF_Out[1]), .CK(CLK), .Q(
        S_10_G_CF_Reg[1]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_2_ ( .D(S_10_G_CF_Out[2]), .CK(CLK), .Q(
        S_10_G_CF_Reg[2]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_3_ ( .D(S_10_G_CF_Out[3]), .CK(CLK), .Q(
        S_10_G_CF_Reg[3]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_4_ ( .D(S_10_G_CF_Out[4]), .CK(CLK), .Q(
        S_10_G_CF_Reg[4]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_5_ ( .D(S_10_G_CF_Out[5]), .CK(CLK), .Q(
        S_10_G_CF_Reg[5]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_6_ ( .D(S_10_G_CF_Out[6]), .CK(CLK), .Q(
        S_10_G_CF_Reg[6]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_7_ ( .D(S_10_G_CF_Out[7]), .CK(CLK), .Q(
        S_10_G_CF_Reg[7]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_8_ ( .D(S_10_G_CF_Out[8]), .CK(CLK), .Q(
        S_10_G_CF_Reg[8]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_9_ ( .D(S_10_G_CF_Out[9]), .CK(CLK), .Q(
        S_10_G_CF_Reg[9]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_10_ ( .D(S_10_G_CF_Out[10]), .CK(CLK), .Q(
        S_10_G_CF_Reg[10]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_11_ ( .D(S_10_G_CF_Out[11]), .CK(CLK), .Q(
        S_10_G_CF_Reg[11]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_12_ ( .D(S_10_G_CF_Out[12]), .CK(CLK), .Q(
        S_10_G_CF_Reg[12]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_13_ ( .D(S_10_G_CF_Out[13]), .CK(CLK), .Q(
        S_10_G_CF_Reg[13]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_14_ ( .D(S_10_G_CF_Out[14]), .CK(CLK), .Q(
        S_10_G_CF_Reg[14]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_15_ ( .D(S_10_G_CF_Out[15]), .CK(CLK), .Q(
        S_10_G_CF_Reg[15]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_16_ ( .D(S_10_G_CF_Out[16]), .CK(CLK), .Q(
        S_10_G_CF_Reg[16]), .QN() );
  DFF_X1 S_10_G_CF_Reg_reg_17_ ( .D(S_10_G_CF_Out[17]), .CK(CLK), .Q(
        S_10_G_CF_Reg[17]), .QN() );
  DFF_X1 S_10_G_out1_reg_2_ ( .D(S_10_Rq1[2]), .CK(CLK), .Q(S_10_G_out1[2]), 
        .QN() );
  DFF_X1 S_10_G_out1_reg_3_ ( .D(S_10_Rq1[3]), .CK(CLK), .Q(S_10_G_out1[3]), 
        .QN() );
  DFF_X1 S_10_G_out2_reg_2_ ( .D(S_10_Rq2[2]), .CK(CLK), .Q(SUB_OUT2[42]), 
        .QN() );
  DFF_X1 S_10_G_out2_reg_3_ ( .D(S_10_Rq2[3]), .CK(CLK), .Q(SUB_OUT2[43]), 
        .QN() );
  DFF_X1 S_10_G_out3_reg_2_ ( .D(S_10_Rq3[2]), .CK(CLK), .Q(SUB_OUT3[42]), 
        .QN() );
  DFF_X1 S_10_G_out3_reg_3_ ( .D(S_10_Rq3[3]), .CK(CLK), .Q(SUB_OUT3[43]), 
        .QN() );
  AND2_X1 S_10_G_Inst_0__CF_Inst_U1 ( .A1(S_10_Rq1[1]), .A2(S_10_Rq1[3]), .ZN(
        S_10_G_CF_Out[0]) );
  NOR2_X1 S_10_G_Inst_1__CF_Inst_U2 ( .A1(S_10_Rq1[3]), .A2(
        S_10_G_Inst_1__CF_Inst_n3), .ZN(S_10_G_CF_Out[1]) );
  INV_X1 S_10_G_Inst_1__CF_Inst_U1 ( .A(S_10_Rq2[1]), .ZN(
        S_10_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_10_G_Inst_2__CF_Inst_U2 ( .A(S_10_G_Inst_2__CF_Inst_n3), .B(
        S_10_Rq2[0]), .ZN(S_10_G_CF_Out[2]) );
  NAND2_X1 S_10_G_Inst_2__CF_Inst_U1 ( .A1(S_10_Rq1[1]), .A2(S_10_Rq2[3]), 
        .ZN(S_10_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_10_G_Inst_3__CF_Inst_U3 ( .A(S_10_Rq1[0]), .B(
        S_10_G_Inst_3__CF_Inst_n6), .ZN(S_10_G_CF_Out[3]) );
  NAND2_X1 S_10_G_Inst_3__CF_Inst_U2 ( .A1(S_10_Rq3[1]), .A2(
        S_10_G_Inst_3__CF_Inst_n5), .ZN(S_10_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_10_G_Inst_3__CF_Inst_U1 ( .A(S_10_Rq1[3]), .ZN(
        S_10_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_10_G_Inst_4__CF_Inst_U1 ( .A1(S_10_Rq2[1]), .A2(S_10_Rq2[3]), .ZN(
        S_10_G_CF_Out[4]) );
  OR2_X1 S_10_G_Inst_5__CF_Inst_U1 ( .A1(S_10_Rq3[3]), .A2(S_10_Rq2[1]), .ZN(
        S_10_G_CF_Out[5]) );
  AND2_X1 S_10_G_Inst_6__CF_Inst_U1 ( .A1(S_10_Rq3[1]), .A2(S_10_Rq2[3]), .ZN(
        S_10_G_CF_Out[6]) );
  XNOR2_X1 S_10_G_Inst_7__CF_Inst_U2 ( .A(S_10_G_Inst_7__CF_Inst_n3), .B(
        S_10_Rq3[0]), .ZN(S_10_G_CF_Out[7]) );
  NAND2_X1 S_10_G_Inst_7__CF_Inst_U1 ( .A1(S_10_Rq1[1]), .A2(S_10_Rq3[3]), 
        .ZN(S_10_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_10_G_Inst_8__CF_Inst_U1 ( .A1(S_10_Rq3[3]), .A2(S_10_Rq3[1]), .ZN(
        S_10_G_CF_Out[8]) );
  NOR2_X1 S_10_G_Inst_9__CF_Inst_U2 ( .A1(S_10_Rq1[3]), .A2(
        S_10_G_Inst_9__CF_Inst_n3), .ZN(S_10_G_CF_Out[9]) );
  INV_X1 S_10_G_Inst_9__CF_Inst_U1 ( .A(S_10_Rq1[2]), .ZN(
        S_10_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_10_G_Inst_10__CF_Inst_U2 ( .A1(S_10_Rq2[2]), .A2(
        S_10_G_Inst_10__CF_Inst_n3), .ZN(S_10_G_CF_Out[10]) );
  INV_X1 S_10_G_Inst_10__CF_Inst_U1 ( .A(S_10_Rq1[3]), .ZN(
        S_10_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_10_G_Inst_11__CF_Inst_U3 ( .A(S_10_Rq1[1]), .B(
        S_10_G_Inst_11__CF_Inst_n6), .ZN(S_10_G_CF_Out[11]) );
  NAND2_X1 S_10_G_Inst_11__CF_Inst_U2 ( .A1(S_10_Rq1[3]), .A2(
        S_10_G_Inst_11__CF_Inst_n5), .ZN(S_10_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_10_G_Inst_11__CF_Inst_U1 ( .A(S_10_Rq3[2]), .ZN(
        S_10_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_10_G_Inst_12__CF_Inst_U2 ( .A1(S_10_Rq2[3]), .A2(
        S_10_G_Inst_12__CF_Inst_n3), .ZN(S_10_G_CF_Out[12]) );
  INV_X1 S_10_G_Inst_12__CF_Inst_U1 ( .A(S_10_Rq1[2]), .ZN(
        S_10_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_10_G_Inst_13__CF_Inst_U1 ( .A1(S_10_Rq2[2]), .A2(S_10_Rq2[3]), 
        .ZN(S_10_G_CF_Out[13]) );
  XNOR2_X1 S_10_G_Inst_14__CF_Inst_U3 ( .A(S_10_Rq2[1]), .B(
        S_10_G_Inst_14__CF_Inst_n6), .ZN(S_10_G_CF_Out[14]) );
  NAND2_X1 S_10_G_Inst_14__CF_Inst_U2 ( .A1(S_10_Rq3[2]), .A2(
        S_10_G_Inst_14__CF_Inst_n5), .ZN(S_10_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_10_G_Inst_14__CF_Inst_U1 ( .A(S_10_Rq2[3]), .ZN(
        S_10_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_10_G_Inst_15__CF_Inst_U2 ( .A(S_10_G_Inst_15__CF_Inst_n3), .B(
        S_10_Rq3[1]), .ZN(S_10_G_CF_Out[15]) );
  NAND2_X1 S_10_G_Inst_15__CF_Inst_U1 ( .A1(S_10_Rq1[2]), .A2(S_10_Rq3[3]), 
        .ZN(S_10_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_10_G_Inst_16__CF_Inst_U1 ( .A1(S_10_Rq2[2]), .A2(S_10_Rq3[3]), 
        .ZN(S_10_G_CF_Out[16]) );
  NOR2_X1 S_10_G_Inst_17__CF_Inst_U2 ( .A1(S_10_Rq3[3]), .A2(
        S_10_G_Inst_17__CF_Inst_n3), .ZN(S_10_G_CF_Out[17]) );
  INV_X1 S_10_G_Inst_17__CF_Inst_U1 ( .A(S_10_Rq3[2]), .ZN(
        S_10_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_10_G_InstXOR_0__Compression1_U2 ( .A(
        S_10_G_InstXOR_0__Compression1_n3), .B(S_10_G_CF_Reg[2]), .ZN(
        S_10_G_out1[0]) );
  XNOR2_X1 S_10_G_InstXOR_0__Compression1_U1 ( .A(S_10_G_CF_Reg[0]), .B(
        S_10_G_CF_Reg[1]), .ZN(S_10_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_10_G_InstXOR_0__Compression2_U2 ( .A(
        S_10_G_InstXOR_0__Compression2_n3), .B(S_10_G_CF_Reg[5]), .ZN(
        SUB_OUT2[41]) );
  XNOR2_X1 S_10_G_InstXOR_0__Compression2_U1 ( .A(S_10_G_CF_Reg[3]), .B(
        S_10_G_CF_Reg[4]), .ZN(S_10_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_10_G_InstXOR_0__Compression3_U2 ( .A(
        S_10_G_InstXOR_0__Compression3_n3), .B(S_10_G_CF_Reg[8]), .ZN(
        SUB_OUT3[41]) );
  XNOR2_X1 S_10_G_InstXOR_0__Compression3_U1 ( .A(S_10_G_CF_Reg[6]), .B(
        S_10_G_CF_Reg[7]), .ZN(S_10_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_10_G_InstXOR_1__Compression1_U2 ( .A(
        S_10_G_InstXOR_1__Compression1_n3), .B(S_10_G_CF_Reg[11]), .ZN(
        S_10_G_out1[1]) );
  XNOR2_X1 S_10_G_InstXOR_1__Compression1_U1 ( .A(S_10_G_CF_Reg[9]), .B(
        S_10_G_CF_Reg[10]), .ZN(S_10_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_10_G_InstXOR_1__Compression2_U2 ( .A(
        S_10_G_InstXOR_1__Compression2_n3), .B(S_10_G_CF_Reg[14]), .ZN(
        SUB_OUT2[40]) );
  XNOR2_X1 S_10_G_InstXOR_1__Compression2_U1 ( .A(S_10_G_CF_Reg[12]), .B(
        S_10_G_CF_Reg[13]), .ZN(S_10_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_10_G_InstXOR_1__Compression3_U2 ( .A(
        S_10_G_InstXOR_1__Compression3_n3), .B(S_10_G_CF_Reg[17]), .ZN(
        SUB_OUT3[40]) );
  XNOR2_X1 S_10_G_InstXOR_1__Compression3_U1 ( .A(S_10_G_CF_Reg[15]), .B(
        S_10_G_CF_Reg[16]), .ZN(S_10_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_10_OutputAffine_U4 ( .A(S_10_G_out1[3]), .ZN(SUB_OUT1[43]) );
  INV_X1 S_10_OutputAffine_U3 ( .A(S_10_G_out1[2]), .ZN(SUB_OUT1[42]) );
  INV_X1 S_10_OutputAffine_U2 ( .A(S_10_G_out1[1]), .ZN(SUB_OUT1[40]) );
  INV_X1 S_10_OutputAffine_U1 ( .A(S_10_G_out1[0]), .ZN(SUB_OUT1[41]) );
  DFF_X1 S_11_Rq3_reg_0_ ( .D(S_11_q3[0]), .CK(CLK), .Q(S_11_Rq3[0]), .QN() );
  DFF_X1 S_11_Rq3_reg_1_ ( .D(S_11_q3[1]), .CK(CLK), .Q(S_11_Rq3[1]), .QN() );
  DFF_X1 S_11_Rq3_reg_2_ ( .D(S_11_q3[2]), .CK(CLK), .Q(S_11_Rq3[2]), .QN() );
  DFF_X1 S_11_Rq3_reg_3_ ( .D(S_11_q3[3]), .CK(CLK), .Q(S_11_Rq3[3]), .QN() );
  DFF_X1 S_11_Rq2_reg_0_ ( .D(S_11_q2[0]), .CK(CLK), .Q(S_11_Rq2[0]), .QN() );
  DFF_X1 S_11_Rq2_reg_1_ ( .D(S_11_q2[1]), .CK(CLK), .Q(S_11_Rq2[1]), .QN() );
  DFF_X1 S_11_Rq2_reg_2_ ( .D(S_11_q2[2]), .CK(CLK), .Q(S_11_Rq2[2]), .QN() );
  DFF_X1 S_11_Rq2_reg_3_ ( .D(S_11_q2[3]), .CK(CLK), .Q(S_11_Rq2[3]), .QN() );
  DFF_X1 S_11_Rq1_reg_0_ ( .D(S_11_q1[0]), .CK(CLK), .Q(S_11_Rq1[0]), .QN() );
  DFF_X1 S_11_Rq1_reg_1_ ( .D(S_11_q1[1]), .CK(CLK), .Q(S_11_Rq1[1]), .QN() );
  DFF_X1 S_11_Rq1_reg_2_ ( .D(S_11_q1[2]), .CK(CLK), .Q(S_11_Rq1[2]), .QN() );
  DFF_X1 S_11_Rq1_reg_3_ ( .D(S_11_q1[3]), .CK(CLK), .Q(S_11_Rq1[3]), .QN() );
  INV_X1 S_11_InputAffine_U4 ( .A(SUB_IN1[44]), .ZN(S_11_F_in1[0]) );
  INV_X1 S_11_InputAffine_U3 ( .A(SUB_IN1[46]), .ZN(S_11_F_in1[3]) );
  INV_X1 S_11_InputAffine_U2 ( .A(SUB_IN1[47]), .ZN(S_11_F_in1[1]) );
  INV_X1 S_11_InputAffine_U1 ( .A(SUB_IN1[45]), .ZN(S_11_F_in1[2]) );
  XNOR2_X1 S_11_F_U18 ( .A(S_11_F_n12), .B(FRESH[91]), .ZN(S_11_q3[3]) );
  XNOR2_X1 S_11_F_U17 ( .A(FRESH[90]), .B(S_11_F_q3[3]), .ZN(S_11_F_n12) );
  XNOR2_X1 S_11_F_U16 ( .A(S_11_F_n11), .B(FRESH[89]), .ZN(S_11_q3[2]) );
  XNOR2_X1 S_11_F_U15 ( .A(FRESH[88]), .B(S_11_F_q3[2]), .ZN(S_11_F_n11) );
  XOR2_X1 S_11_F_U14 ( .A(FRESH[91]), .B(S_11_F_q2[3]), .Z(S_11_q2[3]) );
  XOR2_X1 S_11_F_U13 ( .A(FRESH[89]), .B(S_11_F_q2[2]), .Z(S_11_q2[2]) );
  XOR2_X1 S_11_F_U12 ( .A(FRESH[90]), .B(S_11_F_q1[3]), .Z(S_11_q1[3]) );
  XOR2_X1 S_11_F_U11 ( .A(FRESH[88]), .B(S_11_F_q1[2]), .Z(S_11_q1[2]) );
  XNOR2_X1 S_11_F_U10 ( .A(S_11_F_n10), .B(FRESH[93]), .ZN(S_11_F_N5) );
  XNOR2_X1 S_11_F_U9 ( .A(S_11_F_in3[3]), .B(FRESH[92]), .ZN(S_11_F_n10) );
  XOR2_X1 S_11_F_U8 ( .A(FRESH[93]), .B(S_11_F_in2[3]), .Z(S_11_F_N4) );
  XOR2_X1 S_11_F_U7 ( .A(FRESH[92]), .B(S_11_F_in1[3]), .Z(S_11_F_N3) );
  XNOR2_X1 S_11_F_U6 ( .A(S_11_F_n9), .B(FRESH[95]), .ZN(S_11_F_N2) );
  XNOR2_X1 S_11_F_U5 ( .A(S_11_F_in3[2]), .B(FRESH[94]), .ZN(S_11_F_n9) );
  XOR2_X1 S_11_F_U4 ( .A(FRESH[95]), .B(S_11_F_in2[2]), .Z(S_11_F_N1) );
  XOR2_X1 S_11_F_U3 ( .A(FRESH[94]), .B(S_11_F_in1[2]), .Z(S_11_F_N0) );
  DFF_X1 S_11_F_CF_Reg_reg_0_ ( .D(S_11_F_CF_Out[0]), .CK(CLK), .Q(
        S_11_F_CF_Reg[0]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_1_ ( .D(S_11_F_CF_Out[1]), .CK(CLK), .Q(
        S_11_F_CF_Reg[1]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_2_ ( .D(S_11_F_CF_Out[2]), .CK(CLK), .Q(
        S_11_F_CF_Reg[2]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_3_ ( .D(S_11_F_CF_Out[3]), .CK(CLK), .Q(
        S_11_F_CF_Reg[3]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_4_ ( .D(S_11_F_CF_Out[4]), .CK(CLK), .Q(
        S_11_F_CF_Reg[4]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_5_ ( .D(S_11_F_CF_Out[5]), .CK(CLK), .Q(
        S_11_F_CF_Reg[5]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_6_ ( .D(S_11_F_CF_Out[6]), .CK(CLK), .Q(
        S_11_F_CF_Reg[6]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_7_ ( .D(S_11_F_CF_Out[7]), .CK(CLK), .Q(
        S_11_F_CF_Reg[7]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_8_ ( .D(S_11_F_CF_Out[8]), .CK(CLK), .Q(
        S_11_F_CF_Reg[8]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_9_ ( .D(S_11_F_CF_Out[9]), .CK(CLK), .Q(
        S_11_F_CF_Reg[9]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_10_ ( .D(S_11_F_CF_Out[10]), .CK(CLK), .Q(
        S_11_F_CF_Reg[10]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_11_ ( .D(S_11_F_CF_Out[11]), .CK(CLK), .Q(
        S_11_F_CF_Reg[11]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_12_ ( .D(S_11_F_CF_Out[12]), .CK(CLK), .Q(
        S_11_F_CF_Reg[12]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_13_ ( .D(S_11_F_CF_Out[13]), .CK(CLK), .Q(
        S_11_F_CF_Reg[13]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_14_ ( .D(S_11_F_CF_Out[14]), .CK(CLK), .Q(
        S_11_F_CF_Reg[14]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_15_ ( .D(S_11_F_CF_Out[15]), .CK(CLK), .Q(
        S_11_F_CF_Reg[15]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_16_ ( .D(S_11_F_CF_Out[16]), .CK(CLK), .Q(
        S_11_F_CF_Reg[16]), .QN() );
  DFF_X1 S_11_F_CF_Reg_reg_17_ ( .D(S_11_F_CF_Out[17]), .CK(CLK), .Q(
        S_11_F_CF_Reg[17]), .QN() );
  DFF_X1 S_11_F_out2_reg_0_ ( .D(S_11_F_N4), .CK(CLK), .Q(S_11_q2[0]), .QN()
         );
  DFF_X1 S_11_F_out2_reg_1_ ( .D(S_11_F_N1), .CK(CLK), .Q(S_11_q2[1]), .QN()
         );
  DFF_X1 S_11_F_out3_reg_0_ ( .D(S_11_F_N5), .CK(CLK), .Q(S_11_q3[0]), .QN()
         );
  DFF_X1 S_11_F_out3_reg_1_ ( .D(S_11_F_N2), .CK(CLK), .Q(S_11_q3[1]), .QN()
         );
  DFF_X1 S_11_F_out1_reg_0_ ( .D(S_11_F_N3), .CK(CLK), .Q(S_11_q1[0]), .QN()
         );
  DFF_X1 S_11_F_out1_reg_1_ ( .D(S_11_F_N0), .CK(CLK), .Q(S_11_q1[1]), .QN()
         );
  NOR2_X1 S_11_F_Inst_0__CF_Inst_U2 ( .A1(S_11_F_in1[2]), .A2(
        S_11_F_Inst_0__CF_Inst_n3), .ZN(S_11_F_CF_Out[0]) );
  INV_X1 S_11_F_Inst_0__CF_Inst_U1 ( .A(S_11_F_in1[3]), .ZN(
        S_11_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_11_F_Inst_1__CF_Inst_U2 ( .A(S_11_F_Inst_1__CF_Inst_n3), .B(
        S_11_F_in1[1]), .ZN(S_11_F_CF_Out[1]) );
  NAND2_X1 S_11_F_Inst_1__CF_Inst_U1 ( .A1(S_11_F_in2[2]), .A2(S_11_F_in1[3]), 
        .ZN(S_11_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_11_F_Inst_2__CF_Inst_U1 ( .A1(S_11_F_in1[3]), .A2(S_11_F_in3[2]), 
        .ZN(S_11_F_CF_Out[2]) );
  NOR2_X1 S_11_F_Inst_3__CF_Inst_U2 ( .A1(S_11_F_in2[3]), .A2(
        S_11_F_Inst_3__CF_Inst_n3), .ZN(S_11_F_CF_Out[3]) );
  INV_X1 S_11_F_Inst_3__CF_Inst_U1 ( .A(S_11_F_in1[2]), .ZN(
        S_11_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_11_F_Inst_4__CF_Inst_U2 ( .A(S_11_F_Inst_4__CF_Inst_n3), .B(
        S_11_F_in2[1]), .ZN(S_11_F_CF_Out[4]) );
  NAND2_X1 S_11_F_Inst_4__CF_Inst_U1 ( .A1(S_11_F_in2[2]), .A2(S_11_F_in2[3]), 
        .ZN(S_11_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_11_F_Inst_5__CF_Inst_U1 ( .A1(S_11_F_in3[2]), .A2(S_11_F_in2[3]), 
        .ZN(S_11_F_CF_Out[5]) );
  XNOR2_X1 S_11_F_Inst_6__CF_Inst_U2 ( .A(S_11_F_Inst_6__CF_Inst_n7), .B(
        S_11_F_in3[1]), .ZN(S_11_F_CF_Out[6]) );
  NOR2_X1 S_11_F_Inst_6__CF_Inst_U1 ( .A1(S_11_F_in1[2]), .A2(S_11_F_in3[3]), 
        .ZN(S_11_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_11_F_Inst_7__CF_Inst_U1 ( .A1(S_11_F_in2[2]), .A2(S_11_F_in3[3]), 
        .ZN(S_11_F_CF_Out[7]) );
  OR2_X1 S_11_F_Inst_8__CF_Inst_U1 ( .A1(S_11_F_in3[3]), .A2(S_11_F_in3[2]), 
        .ZN(S_11_F_CF_Out[8]) );
  NOR2_X1 S_11_F_Inst_9__CF_Inst_U2 ( .A1(S_11_F_in1[3]), .A2(
        S_11_F_Inst_9__CF_Inst_n3), .ZN(S_11_F_CF_Out[9]) );
  INV_X1 S_11_F_Inst_9__CF_Inst_U1 ( .A(S_11_F_in1[1]), .ZN(
        S_11_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_11_F_Inst_10__CF_Inst_U1 ( .A1(S_11_F_in2[1]), .A2(S_11_F_in1[3]), 
        .ZN(S_11_F_CF_Out[10]) );
  XNOR2_X1 S_11_F_Inst_11__CF_Inst_U2 ( .A(S_11_F_Inst_11__CF_Inst_n3), .B(
        S_11_F_in1[0]), .ZN(S_11_F_CF_Out[11]) );
  NAND2_X1 S_11_F_Inst_11__CF_Inst_U1 ( .A1(S_11_F_in3[1]), .A2(S_11_F_in1[3]), 
        .ZN(S_11_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_11_F_Inst_12__CF_Inst_U2 ( .A(S_11_F_Inst_12__CF_Inst_n3), .B(
        S_11_F_in2[0]), .ZN(S_11_F_CF_Out[12]) );
  NAND2_X1 S_11_F_Inst_12__CF_Inst_U1 ( .A1(S_11_F_in1[1]), .A2(S_11_F_in2[3]), 
        .ZN(S_11_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_11_F_Inst_13__CF_Inst_U2 ( .A1(S_11_F_in2[3]), .A2(
        S_11_F_Inst_13__CF_Inst_n3), .ZN(S_11_F_CF_Out[13]) );
  INV_X1 S_11_F_Inst_13__CF_Inst_U1 ( .A(S_11_F_in2[1]), .ZN(
        S_11_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_11_F_Inst_14__CF_Inst_U1 ( .A1(S_11_F_in3[1]), .A2(S_11_F_in2[3]), 
        .ZN(S_11_F_CF_Out[14]) );
  XNOR2_X1 S_11_F_Inst_15__CF_Inst_U2 ( .A(S_11_F_Inst_15__CF_Inst_n7), .B(
        S_11_F_in3[0]), .ZN(S_11_F_CF_Out[15]) );
  NOR2_X1 S_11_F_Inst_15__CF_Inst_U1 ( .A1(S_11_F_in1[1]), .A2(S_11_F_in3[3]), 
        .ZN(S_11_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_11_F_Inst_16__CF_Inst_U2 ( .A1(S_11_F_in3[3]), .A2(
        S_11_F_Inst_16__CF_Inst_n3), .ZN(S_11_F_CF_Out[16]) );
  INV_X1 S_11_F_Inst_16__CF_Inst_U1 ( .A(S_11_F_in2[1]), .ZN(
        S_11_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_11_F_Inst_17__CF_Inst_U2 ( .A1(S_11_F_in3[1]), .A2(
        S_11_F_Inst_17__CF_Inst_n3), .ZN(S_11_F_CF_Out[17]) );
  INV_X1 S_11_F_Inst_17__CF_Inst_U1 ( .A(S_11_F_in3[3]), .ZN(
        S_11_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_11_F_InstXOR_0__Compression1_U2 ( .A(
        S_11_F_InstXOR_0__Compression1_n3), .B(S_11_F_CF_Reg[2]), .ZN(
        S_11_F_q1[2]) );
  XNOR2_X1 S_11_F_InstXOR_0__Compression1_U1 ( .A(S_11_F_CF_Reg[0]), .B(
        S_11_F_CF_Reg[1]), .ZN(S_11_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_11_F_InstXOR_0__Compression2_U2 ( .A(
        S_11_F_InstXOR_0__Compression2_n3), .B(S_11_F_CF_Reg[5]), .ZN(
        S_11_F_q2[2]) );
  XNOR2_X1 S_11_F_InstXOR_0__Compression2_U1 ( .A(S_11_F_CF_Reg[3]), .B(
        S_11_F_CF_Reg[4]), .ZN(S_11_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_11_F_InstXOR_0__Compression3_U2 ( .A(
        S_11_F_InstXOR_0__Compression3_n3), .B(S_11_F_CF_Reg[8]), .ZN(
        S_11_F_q3[2]) );
  XNOR2_X1 S_11_F_InstXOR_0__Compression3_U1 ( .A(S_11_F_CF_Reg[6]), .B(
        S_11_F_CF_Reg[7]), .ZN(S_11_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_11_F_InstXOR_1__Compression1_U2 ( .A(
        S_11_F_InstXOR_1__Compression1_n3), .B(S_11_F_CF_Reg[11]), .ZN(
        S_11_F_q1[3]) );
  XNOR2_X1 S_11_F_InstXOR_1__Compression1_U1 ( .A(S_11_F_CF_Reg[9]), .B(
        S_11_F_CF_Reg[10]), .ZN(S_11_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_11_F_InstXOR_1__Compression2_U2 ( .A(
        S_11_F_InstXOR_1__Compression2_n3), .B(S_11_F_CF_Reg[14]), .ZN(
        S_11_F_q2[3]) );
  XNOR2_X1 S_11_F_InstXOR_1__Compression2_U1 ( .A(S_11_F_CF_Reg[12]), .B(
        S_11_F_CF_Reg[13]), .ZN(S_11_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_11_F_InstXOR_1__Compression3_U2 ( .A(
        S_11_F_InstXOR_1__Compression3_n3), .B(S_11_F_CF_Reg[17]), .ZN(
        S_11_F_q3[3]) );
  XNOR2_X1 S_11_F_InstXOR_1__Compression3_U1 ( .A(S_11_F_CF_Reg[15]), .B(
        S_11_F_CF_Reg[16]), .ZN(S_11_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_11_G_CF_Reg_reg_0_ ( .D(S_11_G_CF_Out[0]), .CK(CLK), .Q(
        S_11_G_CF_Reg[0]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_1_ ( .D(S_11_G_CF_Out[1]), .CK(CLK), .Q(
        S_11_G_CF_Reg[1]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_2_ ( .D(S_11_G_CF_Out[2]), .CK(CLK), .Q(
        S_11_G_CF_Reg[2]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_3_ ( .D(S_11_G_CF_Out[3]), .CK(CLK), .Q(
        S_11_G_CF_Reg[3]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_4_ ( .D(S_11_G_CF_Out[4]), .CK(CLK), .Q(
        S_11_G_CF_Reg[4]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_5_ ( .D(S_11_G_CF_Out[5]), .CK(CLK), .Q(
        S_11_G_CF_Reg[5]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_6_ ( .D(S_11_G_CF_Out[6]), .CK(CLK), .Q(
        S_11_G_CF_Reg[6]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_7_ ( .D(S_11_G_CF_Out[7]), .CK(CLK), .Q(
        S_11_G_CF_Reg[7]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_8_ ( .D(S_11_G_CF_Out[8]), .CK(CLK), .Q(
        S_11_G_CF_Reg[8]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_9_ ( .D(S_11_G_CF_Out[9]), .CK(CLK), .Q(
        S_11_G_CF_Reg[9]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_10_ ( .D(S_11_G_CF_Out[10]), .CK(CLK), .Q(
        S_11_G_CF_Reg[10]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_11_ ( .D(S_11_G_CF_Out[11]), .CK(CLK), .Q(
        S_11_G_CF_Reg[11]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_12_ ( .D(S_11_G_CF_Out[12]), .CK(CLK), .Q(
        S_11_G_CF_Reg[12]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_13_ ( .D(S_11_G_CF_Out[13]), .CK(CLK), .Q(
        S_11_G_CF_Reg[13]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_14_ ( .D(S_11_G_CF_Out[14]), .CK(CLK), .Q(
        S_11_G_CF_Reg[14]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_15_ ( .D(S_11_G_CF_Out[15]), .CK(CLK), .Q(
        S_11_G_CF_Reg[15]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_16_ ( .D(S_11_G_CF_Out[16]), .CK(CLK), .Q(
        S_11_G_CF_Reg[16]), .QN() );
  DFF_X1 S_11_G_CF_Reg_reg_17_ ( .D(S_11_G_CF_Out[17]), .CK(CLK), .Q(
        S_11_G_CF_Reg[17]), .QN() );
  DFF_X1 S_11_G_out1_reg_2_ ( .D(S_11_Rq1[2]), .CK(CLK), .Q(S_11_G_out1[2]), 
        .QN() );
  DFF_X1 S_11_G_out1_reg_3_ ( .D(S_11_Rq1[3]), .CK(CLK), .Q(S_11_G_out1[3]), 
        .QN() );
  DFF_X1 S_11_G_out2_reg_2_ ( .D(S_11_Rq2[2]), .CK(CLK), .Q(SUB_OUT2[46]), 
        .QN() );
  DFF_X1 S_11_G_out2_reg_3_ ( .D(S_11_Rq2[3]), .CK(CLK), .Q(SUB_OUT2[47]), 
        .QN() );
  DFF_X1 S_11_G_out3_reg_2_ ( .D(S_11_Rq3[2]), .CK(CLK), .Q(SUB_OUT3[46]), 
        .QN() );
  DFF_X1 S_11_G_out3_reg_3_ ( .D(S_11_Rq3[3]), .CK(CLK), .Q(SUB_OUT3[47]), 
        .QN() );
  AND2_X1 S_11_G_Inst_0__CF_Inst_U1 ( .A1(S_11_Rq1[1]), .A2(S_11_Rq1[3]), .ZN(
        S_11_G_CF_Out[0]) );
  NOR2_X1 S_11_G_Inst_1__CF_Inst_U2 ( .A1(S_11_Rq1[3]), .A2(
        S_11_G_Inst_1__CF_Inst_n3), .ZN(S_11_G_CF_Out[1]) );
  INV_X1 S_11_G_Inst_1__CF_Inst_U1 ( .A(S_11_Rq2[1]), .ZN(
        S_11_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_11_G_Inst_2__CF_Inst_U2 ( .A(S_11_G_Inst_2__CF_Inst_n3), .B(
        S_11_Rq2[0]), .ZN(S_11_G_CF_Out[2]) );
  NAND2_X1 S_11_G_Inst_2__CF_Inst_U1 ( .A1(S_11_Rq1[1]), .A2(S_11_Rq2[3]), 
        .ZN(S_11_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_11_G_Inst_3__CF_Inst_U3 ( .A(S_11_Rq1[0]), .B(
        S_11_G_Inst_3__CF_Inst_n6), .ZN(S_11_G_CF_Out[3]) );
  NAND2_X1 S_11_G_Inst_3__CF_Inst_U2 ( .A1(S_11_Rq3[1]), .A2(
        S_11_G_Inst_3__CF_Inst_n5), .ZN(S_11_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_11_G_Inst_3__CF_Inst_U1 ( .A(S_11_Rq1[3]), .ZN(
        S_11_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_11_G_Inst_4__CF_Inst_U1 ( .A1(S_11_Rq2[1]), .A2(S_11_Rq2[3]), .ZN(
        S_11_G_CF_Out[4]) );
  OR2_X1 S_11_G_Inst_5__CF_Inst_U1 ( .A1(S_11_Rq3[3]), .A2(S_11_Rq2[1]), .ZN(
        S_11_G_CF_Out[5]) );
  AND2_X1 S_11_G_Inst_6__CF_Inst_U1 ( .A1(S_11_Rq3[1]), .A2(S_11_Rq2[3]), .ZN(
        S_11_G_CF_Out[6]) );
  XNOR2_X1 S_11_G_Inst_7__CF_Inst_U2 ( .A(S_11_G_Inst_7__CF_Inst_n3), .B(
        S_11_Rq3[0]), .ZN(S_11_G_CF_Out[7]) );
  NAND2_X1 S_11_G_Inst_7__CF_Inst_U1 ( .A1(S_11_Rq1[1]), .A2(S_11_Rq3[3]), 
        .ZN(S_11_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_11_G_Inst_8__CF_Inst_U1 ( .A1(S_11_Rq3[3]), .A2(S_11_Rq3[1]), .ZN(
        S_11_G_CF_Out[8]) );
  NOR2_X1 S_11_G_Inst_9__CF_Inst_U2 ( .A1(S_11_Rq1[3]), .A2(
        S_11_G_Inst_9__CF_Inst_n3), .ZN(S_11_G_CF_Out[9]) );
  INV_X1 S_11_G_Inst_9__CF_Inst_U1 ( .A(S_11_Rq1[2]), .ZN(
        S_11_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_11_G_Inst_10__CF_Inst_U2 ( .A1(S_11_Rq2[2]), .A2(
        S_11_G_Inst_10__CF_Inst_n3), .ZN(S_11_G_CF_Out[10]) );
  INV_X1 S_11_G_Inst_10__CF_Inst_U1 ( .A(S_11_Rq1[3]), .ZN(
        S_11_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_11_G_Inst_11__CF_Inst_U3 ( .A(S_11_Rq1[1]), .B(
        S_11_G_Inst_11__CF_Inst_n6), .ZN(S_11_G_CF_Out[11]) );
  NAND2_X1 S_11_G_Inst_11__CF_Inst_U2 ( .A1(S_11_Rq1[3]), .A2(
        S_11_G_Inst_11__CF_Inst_n5), .ZN(S_11_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_11_G_Inst_11__CF_Inst_U1 ( .A(S_11_Rq3[2]), .ZN(
        S_11_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_11_G_Inst_12__CF_Inst_U2 ( .A1(S_11_Rq2[3]), .A2(
        S_11_G_Inst_12__CF_Inst_n3), .ZN(S_11_G_CF_Out[12]) );
  INV_X1 S_11_G_Inst_12__CF_Inst_U1 ( .A(S_11_Rq1[2]), .ZN(
        S_11_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_11_G_Inst_13__CF_Inst_U1 ( .A1(S_11_Rq2[2]), .A2(S_11_Rq2[3]), 
        .ZN(S_11_G_CF_Out[13]) );
  XNOR2_X1 S_11_G_Inst_14__CF_Inst_U3 ( .A(S_11_Rq2[1]), .B(
        S_11_G_Inst_14__CF_Inst_n6), .ZN(S_11_G_CF_Out[14]) );
  NAND2_X1 S_11_G_Inst_14__CF_Inst_U2 ( .A1(S_11_Rq3[2]), .A2(
        S_11_G_Inst_14__CF_Inst_n5), .ZN(S_11_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_11_G_Inst_14__CF_Inst_U1 ( .A(S_11_Rq2[3]), .ZN(
        S_11_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_11_G_Inst_15__CF_Inst_U2 ( .A(S_11_G_Inst_15__CF_Inst_n3), .B(
        S_11_Rq3[1]), .ZN(S_11_G_CF_Out[15]) );
  NAND2_X1 S_11_G_Inst_15__CF_Inst_U1 ( .A1(S_11_Rq1[2]), .A2(S_11_Rq3[3]), 
        .ZN(S_11_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_11_G_Inst_16__CF_Inst_U1 ( .A1(S_11_Rq2[2]), .A2(S_11_Rq3[3]), 
        .ZN(S_11_G_CF_Out[16]) );
  NOR2_X1 S_11_G_Inst_17__CF_Inst_U2 ( .A1(S_11_Rq3[3]), .A2(
        S_11_G_Inst_17__CF_Inst_n3), .ZN(S_11_G_CF_Out[17]) );
  INV_X1 S_11_G_Inst_17__CF_Inst_U1 ( .A(S_11_Rq3[2]), .ZN(
        S_11_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_11_G_InstXOR_0__Compression1_U2 ( .A(
        S_11_G_InstXOR_0__Compression1_n3), .B(S_11_G_CF_Reg[2]), .ZN(
        S_11_G_out1[0]) );
  XNOR2_X1 S_11_G_InstXOR_0__Compression1_U1 ( .A(S_11_G_CF_Reg[0]), .B(
        S_11_G_CF_Reg[1]), .ZN(S_11_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_11_G_InstXOR_0__Compression2_U2 ( .A(
        S_11_G_InstXOR_0__Compression2_n3), .B(S_11_G_CF_Reg[5]), .ZN(
        SUB_OUT2[45]) );
  XNOR2_X1 S_11_G_InstXOR_0__Compression2_U1 ( .A(S_11_G_CF_Reg[3]), .B(
        S_11_G_CF_Reg[4]), .ZN(S_11_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_11_G_InstXOR_0__Compression3_U2 ( .A(
        S_11_G_InstXOR_0__Compression3_n3), .B(S_11_G_CF_Reg[8]), .ZN(
        SUB_OUT3[45]) );
  XNOR2_X1 S_11_G_InstXOR_0__Compression3_U1 ( .A(S_11_G_CF_Reg[6]), .B(
        S_11_G_CF_Reg[7]), .ZN(S_11_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_11_G_InstXOR_1__Compression1_U2 ( .A(
        S_11_G_InstXOR_1__Compression1_n3), .B(S_11_G_CF_Reg[11]), .ZN(
        S_11_G_out1[1]) );
  XNOR2_X1 S_11_G_InstXOR_1__Compression1_U1 ( .A(S_11_G_CF_Reg[9]), .B(
        S_11_G_CF_Reg[10]), .ZN(S_11_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_11_G_InstXOR_1__Compression2_U2 ( .A(
        S_11_G_InstXOR_1__Compression2_n3), .B(S_11_G_CF_Reg[14]), .ZN(
        SUB_OUT2[44]) );
  XNOR2_X1 S_11_G_InstXOR_1__Compression2_U1 ( .A(S_11_G_CF_Reg[12]), .B(
        S_11_G_CF_Reg[13]), .ZN(S_11_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_11_G_InstXOR_1__Compression3_U2 ( .A(
        S_11_G_InstXOR_1__Compression3_n3), .B(S_11_G_CF_Reg[17]), .ZN(
        SUB_OUT3[44]) );
  XNOR2_X1 S_11_G_InstXOR_1__Compression3_U1 ( .A(S_11_G_CF_Reg[15]), .B(
        S_11_G_CF_Reg[16]), .ZN(S_11_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_11_OutputAffine_U4 ( .A(S_11_G_out1[3]), .ZN(SUB_OUT1[47]) );
  INV_X1 S_11_OutputAffine_U3 ( .A(S_11_G_out1[2]), .ZN(SUB_OUT1[46]) );
  INV_X1 S_11_OutputAffine_U2 ( .A(S_11_G_out1[1]), .ZN(SUB_OUT1[44]) );
  INV_X1 S_11_OutputAffine_U1 ( .A(S_11_G_out1[0]), .ZN(SUB_OUT1[45]) );
  DFF_X1 S_12_Rq3_reg_0_ ( .D(S_12_q3[0]), .CK(CLK), .Q(S_12_Rq3[0]), .QN() );
  DFF_X1 S_12_Rq3_reg_1_ ( .D(S_12_q3[1]), .CK(CLK), .Q(S_12_Rq3[1]), .QN() );
  DFF_X1 S_12_Rq3_reg_2_ ( .D(S_12_q3[2]), .CK(CLK), .Q(S_12_Rq3[2]), .QN() );
  DFF_X1 S_12_Rq3_reg_3_ ( .D(S_12_q3[3]), .CK(CLK), .Q(S_12_Rq3[3]), .QN() );
  DFF_X1 S_12_Rq2_reg_0_ ( .D(S_12_q2[0]), .CK(CLK), .Q(S_12_Rq2[0]), .QN() );
  DFF_X1 S_12_Rq2_reg_1_ ( .D(S_12_q2[1]), .CK(CLK), .Q(S_12_Rq2[1]), .QN() );
  DFF_X1 S_12_Rq2_reg_2_ ( .D(S_12_q2[2]), .CK(CLK), .Q(S_12_Rq2[2]), .QN() );
  DFF_X1 S_12_Rq2_reg_3_ ( .D(S_12_q2[3]), .CK(CLK), .Q(S_12_Rq2[3]), .QN() );
  DFF_X1 S_12_Rq1_reg_0_ ( .D(S_12_q1[0]), .CK(CLK), .Q(S_12_Rq1[0]), .QN() );
  DFF_X1 S_12_Rq1_reg_1_ ( .D(S_12_q1[1]), .CK(CLK), .Q(S_12_Rq1[1]), .QN() );
  DFF_X1 S_12_Rq1_reg_2_ ( .D(S_12_q1[2]), .CK(CLK), .Q(S_12_Rq1[2]), .QN() );
  DFF_X1 S_12_Rq1_reg_3_ ( .D(S_12_q1[3]), .CK(CLK), .Q(S_12_Rq1[3]), .QN() );
  INV_X1 S_12_InputAffine_U4 ( .A(SUB_IN1[48]), .ZN(S_12_F_in1[0]) );
  INV_X1 S_12_InputAffine_U3 ( .A(SUB_IN1[50]), .ZN(S_12_F_in1[3]) );
  INV_X1 S_12_InputAffine_U2 ( .A(SUB_IN1[51]), .ZN(S_12_F_in1[1]) );
  INV_X1 S_12_InputAffine_U1 ( .A(SUB_IN1[49]), .ZN(S_12_F_in1[2]) );
  XNOR2_X1 S_12_F_U18 ( .A(S_12_F_n12), .B(FRESH[99]), .ZN(S_12_q3[3]) );
  XNOR2_X1 S_12_F_U17 ( .A(FRESH[98]), .B(S_12_F_q3[3]), .ZN(S_12_F_n12) );
  XNOR2_X1 S_12_F_U16 ( .A(S_12_F_n11), .B(FRESH[97]), .ZN(S_12_q3[2]) );
  XNOR2_X1 S_12_F_U15 ( .A(FRESH[96]), .B(S_12_F_q3[2]), .ZN(S_12_F_n11) );
  XOR2_X1 S_12_F_U14 ( .A(FRESH[99]), .B(S_12_F_q2[3]), .Z(S_12_q2[3]) );
  XOR2_X1 S_12_F_U13 ( .A(FRESH[97]), .B(S_12_F_q2[2]), .Z(S_12_q2[2]) );
  XOR2_X1 S_12_F_U12 ( .A(FRESH[98]), .B(S_12_F_q1[3]), .Z(S_12_q1[3]) );
  XOR2_X1 S_12_F_U11 ( .A(FRESH[96]), .B(S_12_F_q1[2]), .Z(S_12_q1[2]) );
  XNOR2_X1 S_12_F_U10 ( .A(S_12_F_n10), .B(FRESH[101]), .ZN(S_12_F_N5) );
  XNOR2_X1 S_12_F_U9 ( .A(S_12_F_in3[3]), .B(FRESH[100]), .ZN(S_12_F_n10) );
  XOR2_X1 S_12_F_U8 ( .A(FRESH[101]), .B(S_12_F_in2[3]), .Z(S_12_F_N4) );
  XOR2_X1 S_12_F_U7 ( .A(FRESH[100]), .B(S_12_F_in1[3]), .Z(S_12_F_N3) );
  XNOR2_X1 S_12_F_U6 ( .A(S_12_F_n9), .B(FRESH[103]), .ZN(S_12_F_N2) );
  XNOR2_X1 S_12_F_U5 ( .A(S_12_F_in3[2]), .B(FRESH[102]), .ZN(S_12_F_n9) );
  XOR2_X1 S_12_F_U4 ( .A(FRESH[103]), .B(S_12_F_in2[2]), .Z(S_12_F_N1) );
  XOR2_X1 S_12_F_U3 ( .A(FRESH[102]), .B(S_12_F_in1[2]), .Z(S_12_F_N0) );
  DFF_X1 S_12_F_CF_Reg_reg_0_ ( .D(S_12_F_CF_Out[0]), .CK(CLK), .Q(
        S_12_F_CF_Reg[0]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_1_ ( .D(S_12_F_CF_Out[1]), .CK(CLK), .Q(
        S_12_F_CF_Reg[1]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_2_ ( .D(S_12_F_CF_Out[2]), .CK(CLK), .Q(
        S_12_F_CF_Reg[2]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_3_ ( .D(S_12_F_CF_Out[3]), .CK(CLK), .Q(
        S_12_F_CF_Reg[3]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_4_ ( .D(S_12_F_CF_Out[4]), .CK(CLK), .Q(
        S_12_F_CF_Reg[4]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_5_ ( .D(S_12_F_CF_Out[5]), .CK(CLK), .Q(
        S_12_F_CF_Reg[5]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_6_ ( .D(S_12_F_CF_Out[6]), .CK(CLK), .Q(
        S_12_F_CF_Reg[6]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_7_ ( .D(S_12_F_CF_Out[7]), .CK(CLK), .Q(
        S_12_F_CF_Reg[7]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_8_ ( .D(S_12_F_CF_Out[8]), .CK(CLK), .Q(
        S_12_F_CF_Reg[8]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_9_ ( .D(S_12_F_CF_Out[9]), .CK(CLK), .Q(
        S_12_F_CF_Reg[9]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_10_ ( .D(S_12_F_CF_Out[10]), .CK(CLK), .Q(
        S_12_F_CF_Reg[10]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_11_ ( .D(S_12_F_CF_Out[11]), .CK(CLK), .Q(
        S_12_F_CF_Reg[11]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_12_ ( .D(S_12_F_CF_Out[12]), .CK(CLK), .Q(
        S_12_F_CF_Reg[12]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_13_ ( .D(S_12_F_CF_Out[13]), .CK(CLK), .Q(
        S_12_F_CF_Reg[13]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_14_ ( .D(S_12_F_CF_Out[14]), .CK(CLK), .Q(
        S_12_F_CF_Reg[14]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_15_ ( .D(S_12_F_CF_Out[15]), .CK(CLK), .Q(
        S_12_F_CF_Reg[15]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_16_ ( .D(S_12_F_CF_Out[16]), .CK(CLK), .Q(
        S_12_F_CF_Reg[16]), .QN() );
  DFF_X1 S_12_F_CF_Reg_reg_17_ ( .D(S_12_F_CF_Out[17]), .CK(CLK), .Q(
        S_12_F_CF_Reg[17]), .QN() );
  DFF_X1 S_12_F_out2_reg_0_ ( .D(S_12_F_N4), .CK(CLK), .Q(S_12_q2[0]), .QN()
         );
  DFF_X1 S_12_F_out2_reg_1_ ( .D(S_12_F_N1), .CK(CLK), .Q(S_12_q2[1]), .QN()
         );
  DFF_X1 S_12_F_out3_reg_0_ ( .D(S_12_F_N5), .CK(CLK), .Q(S_12_q3[0]), .QN()
         );
  DFF_X1 S_12_F_out3_reg_1_ ( .D(S_12_F_N2), .CK(CLK), .Q(S_12_q3[1]), .QN()
         );
  DFF_X1 S_12_F_out1_reg_0_ ( .D(S_12_F_N3), .CK(CLK), .Q(S_12_q1[0]), .QN()
         );
  DFF_X1 S_12_F_out1_reg_1_ ( .D(S_12_F_N0), .CK(CLK), .Q(S_12_q1[1]), .QN()
         );
  NOR2_X1 S_12_F_Inst_0__CF_Inst_U2 ( .A1(S_12_F_in1[2]), .A2(
        S_12_F_Inst_0__CF_Inst_n3), .ZN(S_12_F_CF_Out[0]) );
  INV_X1 S_12_F_Inst_0__CF_Inst_U1 ( .A(S_12_F_in1[3]), .ZN(
        S_12_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_12_F_Inst_1__CF_Inst_U2 ( .A(S_12_F_Inst_1__CF_Inst_n3), .B(
        S_12_F_in1[1]), .ZN(S_12_F_CF_Out[1]) );
  NAND2_X1 S_12_F_Inst_1__CF_Inst_U1 ( .A1(S_12_F_in2[2]), .A2(S_12_F_in1[3]), 
        .ZN(S_12_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_12_F_Inst_2__CF_Inst_U1 ( .A1(S_12_F_in1[3]), .A2(S_12_F_in3[2]), 
        .ZN(S_12_F_CF_Out[2]) );
  NOR2_X1 S_12_F_Inst_3__CF_Inst_U2 ( .A1(S_12_F_in2[3]), .A2(
        S_12_F_Inst_3__CF_Inst_n3), .ZN(S_12_F_CF_Out[3]) );
  INV_X1 S_12_F_Inst_3__CF_Inst_U1 ( .A(S_12_F_in1[2]), .ZN(
        S_12_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_12_F_Inst_4__CF_Inst_U2 ( .A(S_12_F_Inst_4__CF_Inst_n3), .B(
        S_12_F_in2[1]), .ZN(S_12_F_CF_Out[4]) );
  NAND2_X1 S_12_F_Inst_4__CF_Inst_U1 ( .A1(S_12_F_in2[2]), .A2(S_12_F_in2[3]), 
        .ZN(S_12_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_12_F_Inst_5__CF_Inst_U1 ( .A1(S_12_F_in3[2]), .A2(S_12_F_in2[3]), 
        .ZN(S_12_F_CF_Out[5]) );
  XNOR2_X1 S_12_F_Inst_6__CF_Inst_U2 ( .A(S_12_F_Inst_6__CF_Inst_n7), .B(
        S_12_F_in3[1]), .ZN(S_12_F_CF_Out[6]) );
  NOR2_X1 S_12_F_Inst_6__CF_Inst_U1 ( .A1(S_12_F_in1[2]), .A2(S_12_F_in3[3]), 
        .ZN(S_12_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_12_F_Inst_7__CF_Inst_U1 ( .A1(S_12_F_in2[2]), .A2(S_12_F_in3[3]), 
        .ZN(S_12_F_CF_Out[7]) );
  OR2_X1 S_12_F_Inst_8__CF_Inst_U1 ( .A1(S_12_F_in3[3]), .A2(S_12_F_in3[2]), 
        .ZN(S_12_F_CF_Out[8]) );
  NOR2_X1 S_12_F_Inst_9__CF_Inst_U2 ( .A1(S_12_F_in1[3]), .A2(
        S_12_F_Inst_9__CF_Inst_n3), .ZN(S_12_F_CF_Out[9]) );
  INV_X1 S_12_F_Inst_9__CF_Inst_U1 ( .A(S_12_F_in1[1]), .ZN(
        S_12_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_12_F_Inst_10__CF_Inst_U1 ( .A1(S_12_F_in2[1]), .A2(S_12_F_in1[3]), 
        .ZN(S_12_F_CF_Out[10]) );
  XNOR2_X1 S_12_F_Inst_11__CF_Inst_U2 ( .A(S_12_F_Inst_11__CF_Inst_n3), .B(
        S_12_F_in1[0]), .ZN(S_12_F_CF_Out[11]) );
  NAND2_X1 S_12_F_Inst_11__CF_Inst_U1 ( .A1(S_12_F_in3[1]), .A2(S_12_F_in1[3]), 
        .ZN(S_12_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_12_F_Inst_12__CF_Inst_U2 ( .A(S_12_F_Inst_12__CF_Inst_n3), .B(
        S_12_F_in2[0]), .ZN(S_12_F_CF_Out[12]) );
  NAND2_X1 S_12_F_Inst_12__CF_Inst_U1 ( .A1(S_12_F_in1[1]), .A2(S_12_F_in2[3]), 
        .ZN(S_12_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_12_F_Inst_13__CF_Inst_U2 ( .A1(S_12_F_in2[3]), .A2(
        S_12_F_Inst_13__CF_Inst_n3), .ZN(S_12_F_CF_Out[13]) );
  INV_X1 S_12_F_Inst_13__CF_Inst_U1 ( .A(S_12_F_in2[1]), .ZN(
        S_12_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_12_F_Inst_14__CF_Inst_U1 ( .A1(S_12_F_in3[1]), .A2(S_12_F_in2[3]), 
        .ZN(S_12_F_CF_Out[14]) );
  XNOR2_X1 S_12_F_Inst_15__CF_Inst_U2 ( .A(S_12_F_Inst_15__CF_Inst_n7), .B(
        S_12_F_in3[0]), .ZN(S_12_F_CF_Out[15]) );
  NOR2_X1 S_12_F_Inst_15__CF_Inst_U1 ( .A1(S_12_F_in1[1]), .A2(S_12_F_in3[3]), 
        .ZN(S_12_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_12_F_Inst_16__CF_Inst_U2 ( .A1(S_12_F_in3[3]), .A2(
        S_12_F_Inst_16__CF_Inst_n3), .ZN(S_12_F_CF_Out[16]) );
  INV_X1 S_12_F_Inst_16__CF_Inst_U1 ( .A(S_12_F_in2[1]), .ZN(
        S_12_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_12_F_Inst_17__CF_Inst_U2 ( .A1(S_12_F_in3[1]), .A2(
        S_12_F_Inst_17__CF_Inst_n3), .ZN(S_12_F_CF_Out[17]) );
  INV_X1 S_12_F_Inst_17__CF_Inst_U1 ( .A(S_12_F_in3[3]), .ZN(
        S_12_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_12_F_InstXOR_0__Compression1_U2 ( .A(
        S_12_F_InstXOR_0__Compression1_n3), .B(S_12_F_CF_Reg[2]), .ZN(
        S_12_F_q1[2]) );
  XNOR2_X1 S_12_F_InstXOR_0__Compression1_U1 ( .A(S_12_F_CF_Reg[0]), .B(
        S_12_F_CF_Reg[1]), .ZN(S_12_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_12_F_InstXOR_0__Compression2_U2 ( .A(
        S_12_F_InstXOR_0__Compression2_n3), .B(S_12_F_CF_Reg[5]), .ZN(
        S_12_F_q2[2]) );
  XNOR2_X1 S_12_F_InstXOR_0__Compression2_U1 ( .A(S_12_F_CF_Reg[3]), .B(
        S_12_F_CF_Reg[4]), .ZN(S_12_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_12_F_InstXOR_0__Compression3_U2 ( .A(
        S_12_F_InstXOR_0__Compression3_n3), .B(S_12_F_CF_Reg[8]), .ZN(
        S_12_F_q3[2]) );
  XNOR2_X1 S_12_F_InstXOR_0__Compression3_U1 ( .A(S_12_F_CF_Reg[6]), .B(
        S_12_F_CF_Reg[7]), .ZN(S_12_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_12_F_InstXOR_1__Compression1_U2 ( .A(
        S_12_F_InstXOR_1__Compression1_n3), .B(S_12_F_CF_Reg[11]), .ZN(
        S_12_F_q1[3]) );
  XNOR2_X1 S_12_F_InstXOR_1__Compression1_U1 ( .A(S_12_F_CF_Reg[9]), .B(
        S_12_F_CF_Reg[10]), .ZN(S_12_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_12_F_InstXOR_1__Compression2_U2 ( .A(
        S_12_F_InstXOR_1__Compression2_n3), .B(S_12_F_CF_Reg[14]), .ZN(
        S_12_F_q2[3]) );
  XNOR2_X1 S_12_F_InstXOR_1__Compression2_U1 ( .A(S_12_F_CF_Reg[12]), .B(
        S_12_F_CF_Reg[13]), .ZN(S_12_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_12_F_InstXOR_1__Compression3_U2 ( .A(
        S_12_F_InstXOR_1__Compression3_n3), .B(S_12_F_CF_Reg[17]), .ZN(
        S_12_F_q3[3]) );
  XNOR2_X1 S_12_F_InstXOR_1__Compression3_U1 ( .A(S_12_F_CF_Reg[15]), .B(
        S_12_F_CF_Reg[16]), .ZN(S_12_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_12_G_CF_Reg_reg_0_ ( .D(S_12_G_CF_Out[0]), .CK(CLK), .Q(
        S_12_G_CF_Reg[0]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_1_ ( .D(S_12_G_CF_Out[1]), .CK(CLK), .Q(
        S_12_G_CF_Reg[1]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_2_ ( .D(S_12_G_CF_Out[2]), .CK(CLK), .Q(
        S_12_G_CF_Reg[2]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_3_ ( .D(S_12_G_CF_Out[3]), .CK(CLK), .Q(
        S_12_G_CF_Reg[3]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_4_ ( .D(S_12_G_CF_Out[4]), .CK(CLK), .Q(
        S_12_G_CF_Reg[4]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_5_ ( .D(S_12_G_CF_Out[5]), .CK(CLK), .Q(
        S_12_G_CF_Reg[5]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_6_ ( .D(S_12_G_CF_Out[6]), .CK(CLK), .Q(
        S_12_G_CF_Reg[6]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_7_ ( .D(S_12_G_CF_Out[7]), .CK(CLK), .Q(
        S_12_G_CF_Reg[7]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_8_ ( .D(S_12_G_CF_Out[8]), .CK(CLK), .Q(
        S_12_G_CF_Reg[8]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_9_ ( .D(S_12_G_CF_Out[9]), .CK(CLK), .Q(
        S_12_G_CF_Reg[9]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_10_ ( .D(S_12_G_CF_Out[10]), .CK(CLK), .Q(
        S_12_G_CF_Reg[10]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_11_ ( .D(S_12_G_CF_Out[11]), .CK(CLK), .Q(
        S_12_G_CF_Reg[11]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_12_ ( .D(S_12_G_CF_Out[12]), .CK(CLK), .Q(
        S_12_G_CF_Reg[12]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_13_ ( .D(S_12_G_CF_Out[13]), .CK(CLK), .Q(
        S_12_G_CF_Reg[13]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_14_ ( .D(S_12_G_CF_Out[14]), .CK(CLK), .Q(
        S_12_G_CF_Reg[14]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_15_ ( .D(S_12_G_CF_Out[15]), .CK(CLK), .Q(
        S_12_G_CF_Reg[15]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_16_ ( .D(S_12_G_CF_Out[16]), .CK(CLK), .Q(
        S_12_G_CF_Reg[16]), .QN() );
  DFF_X1 S_12_G_CF_Reg_reg_17_ ( .D(S_12_G_CF_Out[17]), .CK(CLK), .Q(
        S_12_G_CF_Reg[17]), .QN() );
  DFF_X1 S_12_G_out1_reg_2_ ( .D(S_12_Rq1[2]), .CK(CLK), .Q(S_12_G_out1[2]), 
        .QN() );
  DFF_X1 S_12_G_out1_reg_3_ ( .D(S_12_Rq1[3]), .CK(CLK), .Q(S_12_G_out1[3]), 
        .QN() );
  DFF_X1 S_12_G_out2_reg_2_ ( .D(S_12_Rq2[2]), .CK(CLK), .Q(SUB_OUT2[50]), 
        .QN() );
  DFF_X1 S_12_G_out2_reg_3_ ( .D(S_12_Rq2[3]), .CK(CLK), .Q(SUB_OUT2[51]), 
        .QN() );
  DFF_X1 S_12_G_out3_reg_2_ ( .D(S_12_Rq3[2]), .CK(CLK), .Q(SUB_OUT3[50]), 
        .QN() );
  DFF_X1 S_12_G_out3_reg_3_ ( .D(S_12_Rq3[3]), .CK(CLK), .Q(SUB_OUT3[51]), 
        .QN() );
  AND2_X1 S_12_G_Inst_0__CF_Inst_U1 ( .A1(S_12_Rq1[1]), .A2(S_12_Rq1[3]), .ZN(
        S_12_G_CF_Out[0]) );
  NOR2_X1 S_12_G_Inst_1__CF_Inst_U2 ( .A1(S_12_Rq1[3]), .A2(
        S_12_G_Inst_1__CF_Inst_n3), .ZN(S_12_G_CF_Out[1]) );
  INV_X1 S_12_G_Inst_1__CF_Inst_U1 ( .A(S_12_Rq2[1]), .ZN(
        S_12_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_12_G_Inst_2__CF_Inst_U2 ( .A(S_12_G_Inst_2__CF_Inst_n3), .B(
        S_12_Rq2[0]), .ZN(S_12_G_CF_Out[2]) );
  NAND2_X1 S_12_G_Inst_2__CF_Inst_U1 ( .A1(S_12_Rq1[1]), .A2(S_12_Rq2[3]), 
        .ZN(S_12_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_12_G_Inst_3__CF_Inst_U3 ( .A(S_12_Rq1[0]), .B(
        S_12_G_Inst_3__CF_Inst_n6), .ZN(S_12_G_CF_Out[3]) );
  NAND2_X1 S_12_G_Inst_3__CF_Inst_U2 ( .A1(S_12_Rq3[1]), .A2(
        S_12_G_Inst_3__CF_Inst_n5), .ZN(S_12_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_12_G_Inst_3__CF_Inst_U1 ( .A(S_12_Rq1[3]), .ZN(
        S_12_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_12_G_Inst_4__CF_Inst_U1 ( .A1(S_12_Rq2[1]), .A2(S_12_Rq2[3]), .ZN(
        S_12_G_CF_Out[4]) );
  OR2_X1 S_12_G_Inst_5__CF_Inst_U1 ( .A1(S_12_Rq3[3]), .A2(S_12_Rq2[1]), .ZN(
        S_12_G_CF_Out[5]) );
  AND2_X1 S_12_G_Inst_6__CF_Inst_U1 ( .A1(S_12_Rq3[1]), .A2(S_12_Rq2[3]), .ZN(
        S_12_G_CF_Out[6]) );
  XNOR2_X1 S_12_G_Inst_7__CF_Inst_U2 ( .A(S_12_G_Inst_7__CF_Inst_n3), .B(
        S_12_Rq3[0]), .ZN(S_12_G_CF_Out[7]) );
  NAND2_X1 S_12_G_Inst_7__CF_Inst_U1 ( .A1(S_12_Rq1[1]), .A2(S_12_Rq3[3]), 
        .ZN(S_12_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_12_G_Inst_8__CF_Inst_U1 ( .A1(S_12_Rq3[3]), .A2(S_12_Rq3[1]), .ZN(
        S_12_G_CF_Out[8]) );
  NOR2_X1 S_12_G_Inst_9__CF_Inst_U2 ( .A1(S_12_Rq1[3]), .A2(
        S_12_G_Inst_9__CF_Inst_n3), .ZN(S_12_G_CF_Out[9]) );
  INV_X1 S_12_G_Inst_9__CF_Inst_U1 ( .A(S_12_Rq1[2]), .ZN(
        S_12_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_12_G_Inst_10__CF_Inst_U2 ( .A1(S_12_Rq2[2]), .A2(
        S_12_G_Inst_10__CF_Inst_n3), .ZN(S_12_G_CF_Out[10]) );
  INV_X1 S_12_G_Inst_10__CF_Inst_U1 ( .A(S_12_Rq1[3]), .ZN(
        S_12_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_12_G_Inst_11__CF_Inst_U3 ( .A(S_12_Rq1[1]), .B(
        S_12_G_Inst_11__CF_Inst_n6), .ZN(S_12_G_CF_Out[11]) );
  NAND2_X1 S_12_G_Inst_11__CF_Inst_U2 ( .A1(S_12_Rq1[3]), .A2(
        S_12_G_Inst_11__CF_Inst_n5), .ZN(S_12_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_12_G_Inst_11__CF_Inst_U1 ( .A(S_12_Rq3[2]), .ZN(
        S_12_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_12_G_Inst_12__CF_Inst_U2 ( .A1(S_12_Rq2[3]), .A2(
        S_12_G_Inst_12__CF_Inst_n3), .ZN(S_12_G_CF_Out[12]) );
  INV_X1 S_12_G_Inst_12__CF_Inst_U1 ( .A(S_12_Rq1[2]), .ZN(
        S_12_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_12_G_Inst_13__CF_Inst_U1 ( .A1(S_12_Rq2[2]), .A2(S_12_Rq2[3]), 
        .ZN(S_12_G_CF_Out[13]) );
  XNOR2_X1 S_12_G_Inst_14__CF_Inst_U3 ( .A(S_12_Rq2[1]), .B(
        S_12_G_Inst_14__CF_Inst_n6), .ZN(S_12_G_CF_Out[14]) );
  NAND2_X1 S_12_G_Inst_14__CF_Inst_U2 ( .A1(S_12_Rq3[2]), .A2(
        S_12_G_Inst_14__CF_Inst_n5), .ZN(S_12_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_12_G_Inst_14__CF_Inst_U1 ( .A(S_12_Rq2[3]), .ZN(
        S_12_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_12_G_Inst_15__CF_Inst_U2 ( .A(S_12_G_Inst_15__CF_Inst_n3), .B(
        S_12_Rq3[1]), .ZN(S_12_G_CF_Out[15]) );
  NAND2_X1 S_12_G_Inst_15__CF_Inst_U1 ( .A1(S_12_Rq1[2]), .A2(S_12_Rq3[3]), 
        .ZN(S_12_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_12_G_Inst_16__CF_Inst_U1 ( .A1(S_12_Rq2[2]), .A2(S_12_Rq3[3]), 
        .ZN(S_12_G_CF_Out[16]) );
  NOR2_X1 S_12_G_Inst_17__CF_Inst_U2 ( .A1(S_12_Rq3[3]), .A2(
        S_12_G_Inst_17__CF_Inst_n3), .ZN(S_12_G_CF_Out[17]) );
  INV_X1 S_12_G_Inst_17__CF_Inst_U1 ( .A(S_12_Rq3[2]), .ZN(
        S_12_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_12_G_InstXOR_0__Compression1_U2 ( .A(
        S_12_G_InstXOR_0__Compression1_n3), .B(S_12_G_CF_Reg[2]), .ZN(
        S_12_G_out1[0]) );
  XNOR2_X1 S_12_G_InstXOR_0__Compression1_U1 ( .A(S_12_G_CF_Reg[0]), .B(
        S_12_G_CF_Reg[1]), .ZN(S_12_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_12_G_InstXOR_0__Compression2_U2 ( .A(
        S_12_G_InstXOR_0__Compression2_n3), .B(S_12_G_CF_Reg[5]), .ZN(
        SUB_OUT2[49]) );
  XNOR2_X1 S_12_G_InstXOR_0__Compression2_U1 ( .A(S_12_G_CF_Reg[3]), .B(
        S_12_G_CF_Reg[4]), .ZN(S_12_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_12_G_InstXOR_0__Compression3_U2 ( .A(
        S_12_G_InstXOR_0__Compression3_n3), .B(S_12_G_CF_Reg[8]), .ZN(
        SUB_OUT3[49]) );
  XNOR2_X1 S_12_G_InstXOR_0__Compression3_U1 ( .A(S_12_G_CF_Reg[6]), .B(
        S_12_G_CF_Reg[7]), .ZN(S_12_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_12_G_InstXOR_1__Compression1_U2 ( .A(
        S_12_G_InstXOR_1__Compression1_n3), .B(S_12_G_CF_Reg[11]), .ZN(
        S_12_G_out1[1]) );
  XNOR2_X1 S_12_G_InstXOR_1__Compression1_U1 ( .A(S_12_G_CF_Reg[9]), .B(
        S_12_G_CF_Reg[10]), .ZN(S_12_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_12_G_InstXOR_1__Compression2_U2 ( .A(
        S_12_G_InstXOR_1__Compression2_n3), .B(S_12_G_CF_Reg[14]), .ZN(
        SUB_OUT2[48]) );
  XNOR2_X1 S_12_G_InstXOR_1__Compression2_U1 ( .A(S_12_G_CF_Reg[12]), .B(
        S_12_G_CF_Reg[13]), .ZN(S_12_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_12_G_InstXOR_1__Compression3_U2 ( .A(
        S_12_G_InstXOR_1__Compression3_n3), .B(S_12_G_CF_Reg[17]), .ZN(
        SUB_OUT3[48]) );
  XNOR2_X1 S_12_G_InstXOR_1__Compression3_U1 ( .A(S_12_G_CF_Reg[15]), .B(
        S_12_G_CF_Reg[16]), .ZN(S_12_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_12_OutputAffine_U4 ( .A(S_12_G_out1[3]), .ZN(SUB_OUT1[51]) );
  INV_X1 S_12_OutputAffine_U3 ( .A(S_12_G_out1[2]), .ZN(SUB_OUT1[50]) );
  INV_X1 S_12_OutputAffine_U2 ( .A(S_12_G_out1[1]), .ZN(SUB_OUT1[48]) );
  INV_X1 S_12_OutputAffine_U1 ( .A(S_12_G_out1[0]), .ZN(SUB_OUT1[49]) );
  DFF_X1 S_13_Rq3_reg_0_ ( .D(S_13_q3[0]), .CK(CLK), .Q(S_13_Rq3[0]), .QN() );
  DFF_X1 S_13_Rq3_reg_1_ ( .D(S_13_q3[1]), .CK(CLK), .Q(S_13_Rq3[1]), .QN() );
  DFF_X1 S_13_Rq3_reg_2_ ( .D(S_13_q3[2]), .CK(CLK), .Q(S_13_Rq3[2]), .QN() );
  DFF_X1 S_13_Rq3_reg_3_ ( .D(S_13_q3[3]), .CK(CLK), .Q(S_13_Rq3[3]), .QN() );
  DFF_X1 S_13_Rq2_reg_0_ ( .D(S_13_q2[0]), .CK(CLK), .Q(S_13_Rq2[0]), .QN() );
  DFF_X1 S_13_Rq2_reg_1_ ( .D(S_13_q2[1]), .CK(CLK), .Q(S_13_Rq2[1]), .QN() );
  DFF_X1 S_13_Rq2_reg_2_ ( .D(S_13_q2[2]), .CK(CLK), .Q(S_13_Rq2[2]), .QN() );
  DFF_X1 S_13_Rq2_reg_3_ ( .D(S_13_q2[3]), .CK(CLK), .Q(S_13_Rq2[3]), .QN() );
  DFF_X1 S_13_Rq1_reg_0_ ( .D(S_13_q1[0]), .CK(CLK), .Q(S_13_Rq1[0]), .QN() );
  DFF_X1 S_13_Rq1_reg_1_ ( .D(S_13_q1[1]), .CK(CLK), .Q(S_13_Rq1[1]), .QN() );
  DFF_X1 S_13_Rq1_reg_2_ ( .D(S_13_q1[2]), .CK(CLK), .Q(S_13_Rq1[2]), .QN() );
  DFF_X1 S_13_Rq1_reg_3_ ( .D(S_13_q1[3]), .CK(CLK), .Q(S_13_Rq1[3]), .QN() );
  INV_X1 S_13_InputAffine_U4 ( .A(SUB_IN1[52]), .ZN(S_13_F_in1[0]) );
  INV_X1 S_13_InputAffine_U3 ( .A(SUB_IN1[54]), .ZN(S_13_F_in1[3]) );
  INV_X1 S_13_InputAffine_U2 ( .A(SUB_IN1[55]), .ZN(S_13_F_in1[1]) );
  INV_X1 S_13_InputAffine_U1 ( .A(SUB_IN1[53]), .ZN(S_13_F_in1[2]) );
  XNOR2_X1 S_13_F_U18 ( .A(S_13_F_n12), .B(FRESH[107]), .ZN(S_13_q3[3]) );
  XNOR2_X1 S_13_F_U17 ( .A(FRESH[106]), .B(S_13_F_q3[3]), .ZN(S_13_F_n12) );
  XNOR2_X1 S_13_F_U16 ( .A(S_13_F_n11), .B(FRESH[105]), .ZN(S_13_q3[2]) );
  XNOR2_X1 S_13_F_U15 ( .A(FRESH[104]), .B(S_13_F_q3[2]), .ZN(S_13_F_n11) );
  XOR2_X1 S_13_F_U14 ( .A(FRESH[107]), .B(S_13_F_q2[3]), .Z(S_13_q2[3]) );
  XOR2_X1 S_13_F_U13 ( .A(FRESH[105]), .B(S_13_F_q2[2]), .Z(S_13_q2[2]) );
  XOR2_X1 S_13_F_U12 ( .A(FRESH[106]), .B(S_13_F_q1[3]), .Z(S_13_q1[3]) );
  XOR2_X1 S_13_F_U11 ( .A(FRESH[104]), .B(S_13_F_q1[2]), .Z(S_13_q1[2]) );
  XNOR2_X1 S_13_F_U10 ( .A(S_13_F_n10), .B(FRESH[109]), .ZN(S_13_F_N5) );
  XNOR2_X1 S_13_F_U9 ( .A(S_13_F_in3[3]), .B(FRESH[108]), .ZN(S_13_F_n10) );
  XOR2_X1 S_13_F_U8 ( .A(FRESH[109]), .B(S_13_F_in2[3]), .Z(S_13_F_N4) );
  XOR2_X1 S_13_F_U7 ( .A(FRESH[108]), .B(S_13_F_in1[3]), .Z(S_13_F_N3) );
  XNOR2_X1 S_13_F_U6 ( .A(S_13_F_n9), .B(FRESH[111]), .ZN(S_13_F_N2) );
  XNOR2_X1 S_13_F_U5 ( .A(S_13_F_in3[2]), .B(FRESH[110]), .ZN(S_13_F_n9) );
  XOR2_X1 S_13_F_U4 ( .A(FRESH[111]), .B(S_13_F_in2[2]), .Z(S_13_F_N1) );
  XOR2_X1 S_13_F_U3 ( .A(FRESH[110]), .B(S_13_F_in1[2]), .Z(S_13_F_N0) );
  DFF_X1 S_13_F_CF_Reg_reg_0_ ( .D(S_13_F_CF_Out[0]), .CK(CLK), .Q(
        S_13_F_CF_Reg[0]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_1_ ( .D(S_13_F_CF_Out[1]), .CK(CLK), .Q(
        S_13_F_CF_Reg[1]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_2_ ( .D(S_13_F_CF_Out[2]), .CK(CLK), .Q(
        S_13_F_CF_Reg[2]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_3_ ( .D(S_13_F_CF_Out[3]), .CK(CLK), .Q(
        S_13_F_CF_Reg[3]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_4_ ( .D(S_13_F_CF_Out[4]), .CK(CLK), .Q(
        S_13_F_CF_Reg[4]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_5_ ( .D(S_13_F_CF_Out[5]), .CK(CLK), .Q(
        S_13_F_CF_Reg[5]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_6_ ( .D(S_13_F_CF_Out[6]), .CK(CLK), .Q(
        S_13_F_CF_Reg[6]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_7_ ( .D(S_13_F_CF_Out[7]), .CK(CLK), .Q(
        S_13_F_CF_Reg[7]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_8_ ( .D(S_13_F_CF_Out[8]), .CK(CLK), .Q(
        S_13_F_CF_Reg[8]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_9_ ( .D(S_13_F_CF_Out[9]), .CK(CLK), .Q(
        S_13_F_CF_Reg[9]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_10_ ( .D(S_13_F_CF_Out[10]), .CK(CLK), .Q(
        S_13_F_CF_Reg[10]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_11_ ( .D(S_13_F_CF_Out[11]), .CK(CLK), .Q(
        S_13_F_CF_Reg[11]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_12_ ( .D(S_13_F_CF_Out[12]), .CK(CLK), .Q(
        S_13_F_CF_Reg[12]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_13_ ( .D(S_13_F_CF_Out[13]), .CK(CLK), .Q(
        S_13_F_CF_Reg[13]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_14_ ( .D(S_13_F_CF_Out[14]), .CK(CLK), .Q(
        S_13_F_CF_Reg[14]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_15_ ( .D(S_13_F_CF_Out[15]), .CK(CLK), .Q(
        S_13_F_CF_Reg[15]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_16_ ( .D(S_13_F_CF_Out[16]), .CK(CLK), .Q(
        S_13_F_CF_Reg[16]), .QN() );
  DFF_X1 S_13_F_CF_Reg_reg_17_ ( .D(S_13_F_CF_Out[17]), .CK(CLK), .Q(
        S_13_F_CF_Reg[17]), .QN() );
  DFF_X1 S_13_F_out2_reg_0_ ( .D(S_13_F_N4), .CK(CLK), .Q(S_13_q2[0]), .QN()
         );
  DFF_X1 S_13_F_out2_reg_1_ ( .D(S_13_F_N1), .CK(CLK), .Q(S_13_q2[1]), .QN()
         );
  DFF_X1 S_13_F_out3_reg_0_ ( .D(S_13_F_N5), .CK(CLK), .Q(S_13_q3[0]), .QN()
         );
  DFF_X1 S_13_F_out3_reg_1_ ( .D(S_13_F_N2), .CK(CLK), .Q(S_13_q3[1]), .QN()
         );
  DFF_X1 S_13_F_out1_reg_0_ ( .D(S_13_F_N3), .CK(CLK), .Q(S_13_q1[0]), .QN()
         );
  DFF_X1 S_13_F_out1_reg_1_ ( .D(S_13_F_N0), .CK(CLK), .Q(S_13_q1[1]), .QN()
         );
  NOR2_X1 S_13_F_Inst_0__CF_Inst_U2 ( .A1(S_13_F_in1[2]), .A2(
        S_13_F_Inst_0__CF_Inst_n3), .ZN(S_13_F_CF_Out[0]) );
  INV_X1 S_13_F_Inst_0__CF_Inst_U1 ( .A(S_13_F_in1[3]), .ZN(
        S_13_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_13_F_Inst_1__CF_Inst_U2 ( .A(S_13_F_Inst_1__CF_Inst_n3), .B(
        S_13_F_in1[1]), .ZN(S_13_F_CF_Out[1]) );
  NAND2_X1 S_13_F_Inst_1__CF_Inst_U1 ( .A1(S_13_F_in2[2]), .A2(S_13_F_in1[3]), 
        .ZN(S_13_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_13_F_Inst_2__CF_Inst_U1 ( .A1(S_13_F_in1[3]), .A2(S_13_F_in3[2]), 
        .ZN(S_13_F_CF_Out[2]) );
  NOR2_X1 S_13_F_Inst_3__CF_Inst_U2 ( .A1(S_13_F_in2[3]), .A2(
        S_13_F_Inst_3__CF_Inst_n3), .ZN(S_13_F_CF_Out[3]) );
  INV_X1 S_13_F_Inst_3__CF_Inst_U1 ( .A(S_13_F_in1[2]), .ZN(
        S_13_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_13_F_Inst_4__CF_Inst_U2 ( .A(S_13_F_Inst_4__CF_Inst_n3), .B(
        S_13_F_in2[1]), .ZN(S_13_F_CF_Out[4]) );
  NAND2_X1 S_13_F_Inst_4__CF_Inst_U1 ( .A1(S_13_F_in2[2]), .A2(S_13_F_in2[3]), 
        .ZN(S_13_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_13_F_Inst_5__CF_Inst_U1 ( .A1(S_13_F_in3[2]), .A2(S_13_F_in2[3]), 
        .ZN(S_13_F_CF_Out[5]) );
  XNOR2_X1 S_13_F_Inst_6__CF_Inst_U2 ( .A(S_13_F_Inst_6__CF_Inst_n7), .B(
        S_13_F_in3[1]), .ZN(S_13_F_CF_Out[6]) );
  NOR2_X1 S_13_F_Inst_6__CF_Inst_U1 ( .A1(S_13_F_in1[2]), .A2(S_13_F_in3[3]), 
        .ZN(S_13_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_13_F_Inst_7__CF_Inst_U1 ( .A1(S_13_F_in2[2]), .A2(S_13_F_in3[3]), 
        .ZN(S_13_F_CF_Out[7]) );
  OR2_X1 S_13_F_Inst_8__CF_Inst_U1 ( .A1(S_13_F_in3[3]), .A2(S_13_F_in3[2]), 
        .ZN(S_13_F_CF_Out[8]) );
  NOR2_X1 S_13_F_Inst_9__CF_Inst_U2 ( .A1(S_13_F_in1[3]), .A2(
        S_13_F_Inst_9__CF_Inst_n3), .ZN(S_13_F_CF_Out[9]) );
  INV_X1 S_13_F_Inst_9__CF_Inst_U1 ( .A(S_13_F_in1[1]), .ZN(
        S_13_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_13_F_Inst_10__CF_Inst_U1 ( .A1(S_13_F_in2[1]), .A2(S_13_F_in1[3]), 
        .ZN(S_13_F_CF_Out[10]) );
  XNOR2_X1 S_13_F_Inst_11__CF_Inst_U2 ( .A(S_13_F_Inst_11__CF_Inst_n3), .B(
        S_13_F_in1[0]), .ZN(S_13_F_CF_Out[11]) );
  NAND2_X1 S_13_F_Inst_11__CF_Inst_U1 ( .A1(S_13_F_in3[1]), .A2(S_13_F_in1[3]), 
        .ZN(S_13_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_13_F_Inst_12__CF_Inst_U2 ( .A(S_13_F_Inst_12__CF_Inst_n3), .B(
        S_13_F_in2[0]), .ZN(S_13_F_CF_Out[12]) );
  NAND2_X1 S_13_F_Inst_12__CF_Inst_U1 ( .A1(S_13_F_in1[1]), .A2(S_13_F_in2[3]), 
        .ZN(S_13_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_13_F_Inst_13__CF_Inst_U2 ( .A1(S_13_F_in2[3]), .A2(
        S_13_F_Inst_13__CF_Inst_n3), .ZN(S_13_F_CF_Out[13]) );
  INV_X1 S_13_F_Inst_13__CF_Inst_U1 ( .A(S_13_F_in2[1]), .ZN(
        S_13_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_13_F_Inst_14__CF_Inst_U1 ( .A1(S_13_F_in3[1]), .A2(S_13_F_in2[3]), 
        .ZN(S_13_F_CF_Out[14]) );
  XNOR2_X1 S_13_F_Inst_15__CF_Inst_U2 ( .A(S_13_F_Inst_15__CF_Inst_n7), .B(
        S_13_F_in3[0]), .ZN(S_13_F_CF_Out[15]) );
  NOR2_X1 S_13_F_Inst_15__CF_Inst_U1 ( .A1(S_13_F_in1[1]), .A2(S_13_F_in3[3]), 
        .ZN(S_13_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_13_F_Inst_16__CF_Inst_U2 ( .A1(S_13_F_in3[3]), .A2(
        S_13_F_Inst_16__CF_Inst_n3), .ZN(S_13_F_CF_Out[16]) );
  INV_X1 S_13_F_Inst_16__CF_Inst_U1 ( .A(S_13_F_in2[1]), .ZN(
        S_13_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_13_F_Inst_17__CF_Inst_U2 ( .A1(S_13_F_in3[1]), .A2(
        S_13_F_Inst_17__CF_Inst_n3), .ZN(S_13_F_CF_Out[17]) );
  INV_X1 S_13_F_Inst_17__CF_Inst_U1 ( .A(S_13_F_in3[3]), .ZN(
        S_13_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_13_F_InstXOR_0__Compression1_U2 ( .A(
        S_13_F_InstXOR_0__Compression1_n3), .B(S_13_F_CF_Reg[2]), .ZN(
        S_13_F_q1[2]) );
  XNOR2_X1 S_13_F_InstXOR_0__Compression1_U1 ( .A(S_13_F_CF_Reg[0]), .B(
        S_13_F_CF_Reg[1]), .ZN(S_13_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_13_F_InstXOR_0__Compression2_U2 ( .A(
        S_13_F_InstXOR_0__Compression2_n3), .B(S_13_F_CF_Reg[5]), .ZN(
        S_13_F_q2[2]) );
  XNOR2_X1 S_13_F_InstXOR_0__Compression2_U1 ( .A(S_13_F_CF_Reg[3]), .B(
        S_13_F_CF_Reg[4]), .ZN(S_13_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_13_F_InstXOR_0__Compression3_U2 ( .A(
        S_13_F_InstXOR_0__Compression3_n3), .B(S_13_F_CF_Reg[8]), .ZN(
        S_13_F_q3[2]) );
  XNOR2_X1 S_13_F_InstXOR_0__Compression3_U1 ( .A(S_13_F_CF_Reg[6]), .B(
        S_13_F_CF_Reg[7]), .ZN(S_13_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_13_F_InstXOR_1__Compression1_U2 ( .A(
        S_13_F_InstXOR_1__Compression1_n3), .B(S_13_F_CF_Reg[11]), .ZN(
        S_13_F_q1[3]) );
  XNOR2_X1 S_13_F_InstXOR_1__Compression1_U1 ( .A(S_13_F_CF_Reg[9]), .B(
        S_13_F_CF_Reg[10]), .ZN(S_13_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_13_F_InstXOR_1__Compression2_U2 ( .A(
        S_13_F_InstXOR_1__Compression2_n3), .B(S_13_F_CF_Reg[14]), .ZN(
        S_13_F_q2[3]) );
  XNOR2_X1 S_13_F_InstXOR_1__Compression2_U1 ( .A(S_13_F_CF_Reg[12]), .B(
        S_13_F_CF_Reg[13]), .ZN(S_13_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_13_F_InstXOR_1__Compression3_U2 ( .A(
        S_13_F_InstXOR_1__Compression3_n3), .B(S_13_F_CF_Reg[17]), .ZN(
        S_13_F_q3[3]) );
  XNOR2_X1 S_13_F_InstXOR_1__Compression3_U1 ( .A(S_13_F_CF_Reg[15]), .B(
        S_13_F_CF_Reg[16]), .ZN(S_13_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_13_G_CF_Reg_reg_0_ ( .D(S_13_G_CF_Out[0]), .CK(CLK), .Q(
        S_13_G_CF_Reg[0]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_1_ ( .D(S_13_G_CF_Out[1]), .CK(CLK), .Q(
        S_13_G_CF_Reg[1]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_2_ ( .D(S_13_G_CF_Out[2]), .CK(CLK), .Q(
        S_13_G_CF_Reg[2]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_3_ ( .D(S_13_G_CF_Out[3]), .CK(CLK), .Q(
        S_13_G_CF_Reg[3]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_4_ ( .D(S_13_G_CF_Out[4]), .CK(CLK), .Q(
        S_13_G_CF_Reg[4]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_5_ ( .D(S_13_G_CF_Out[5]), .CK(CLK), .Q(
        S_13_G_CF_Reg[5]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_6_ ( .D(S_13_G_CF_Out[6]), .CK(CLK), .Q(
        S_13_G_CF_Reg[6]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_7_ ( .D(S_13_G_CF_Out[7]), .CK(CLK), .Q(
        S_13_G_CF_Reg[7]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_8_ ( .D(S_13_G_CF_Out[8]), .CK(CLK), .Q(
        S_13_G_CF_Reg[8]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_9_ ( .D(S_13_G_CF_Out[9]), .CK(CLK), .Q(
        S_13_G_CF_Reg[9]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_10_ ( .D(S_13_G_CF_Out[10]), .CK(CLK), .Q(
        S_13_G_CF_Reg[10]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_11_ ( .D(S_13_G_CF_Out[11]), .CK(CLK), .Q(
        S_13_G_CF_Reg[11]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_12_ ( .D(S_13_G_CF_Out[12]), .CK(CLK), .Q(
        S_13_G_CF_Reg[12]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_13_ ( .D(S_13_G_CF_Out[13]), .CK(CLK), .Q(
        S_13_G_CF_Reg[13]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_14_ ( .D(S_13_G_CF_Out[14]), .CK(CLK), .Q(
        S_13_G_CF_Reg[14]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_15_ ( .D(S_13_G_CF_Out[15]), .CK(CLK), .Q(
        S_13_G_CF_Reg[15]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_16_ ( .D(S_13_G_CF_Out[16]), .CK(CLK), .Q(
        S_13_G_CF_Reg[16]), .QN() );
  DFF_X1 S_13_G_CF_Reg_reg_17_ ( .D(S_13_G_CF_Out[17]), .CK(CLK), .Q(
        S_13_G_CF_Reg[17]), .QN() );
  DFF_X1 S_13_G_out1_reg_2_ ( .D(S_13_Rq1[2]), .CK(CLK), .Q(S_13_G_out1[2]), 
        .QN() );
  DFF_X1 S_13_G_out1_reg_3_ ( .D(S_13_Rq1[3]), .CK(CLK), .Q(S_13_G_out1[3]), 
        .QN() );
  DFF_X1 S_13_G_out2_reg_2_ ( .D(S_13_Rq2[2]), .CK(CLK), .Q(SUB_OUT2[54]), 
        .QN() );
  DFF_X1 S_13_G_out2_reg_3_ ( .D(S_13_Rq2[3]), .CK(CLK), .Q(SUB_OUT2[55]), 
        .QN() );
  DFF_X1 S_13_G_out3_reg_2_ ( .D(S_13_Rq3[2]), .CK(CLK), .Q(SUB_OUT3[54]), 
        .QN() );
  DFF_X1 S_13_G_out3_reg_3_ ( .D(S_13_Rq3[3]), .CK(CLK), .Q(SUB_OUT3[55]), 
        .QN() );
  AND2_X1 S_13_G_Inst_0__CF_Inst_U1 ( .A1(S_13_Rq1[1]), .A2(S_13_Rq1[3]), .ZN(
        S_13_G_CF_Out[0]) );
  NOR2_X1 S_13_G_Inst_1__CF_Inst_U2 ( .A1(S_13_Rq1[3]), .A2(
        S_13_G_Inst_1__CF_Inst_n3), .ZN(S_13_G_CF_Out[1]) );
  INV_X1 S_13_G_Inst_1__CF_Inst_U1 ( .A(S_13_Rq2[1]), .ZN(
        S_13_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_13_G_Inst_2__CF_Inst_U2 ( .A(S_13_G_Inst_2__CF_Inst_n3), .B(
        S_13_Rq2[0]), .ZN(S_13_G_CF_Out[2]) );
  NAND2_X1 S_13_G_Inst_2__CF_Inst_U1 ( .A1(S_13_Rq1[1]), .A2(S_13_Rq2[3]), 
        .ZN(S_13_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_13_G_Inst_3__CF_Inst_U3 ( .A(S_13_Rq1[0]), .B(
        S_13_G_Inst_3__CF_Inst_n6), .ZN(S_13_G_CF_Out[3]) );
  NAND2_X1 S_13_G_Inst_3__CF_Inst_U2 ( .A1(S_13_Rq3[1]), .A2(
        S_13_G_Inst_3__CF_Inst_n5), .ZN(S_13_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_13_G_Inst_3__CF_Inst_U1 ( .A(S_13_Rq1[3]), .ZN(
        S_13_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_13_G_Inst_4__CF_Inst_U1 ( .A1(S_13_Rq2[1]), .A2(S_13_Rq2[3]), .ZN(
        S_13_G_CF_Out[4]) );
  OR2_X1 S_13_G_Inst_5__CF_Inst_U1 ( .A1(S_13_Rq3[3]), .A2(S_13_Rq2[1]), .ZN(
        S_13_G_CF_Out[5]) );
  AND2_X1 S_13_G_Inst_6__CF_Inst_U1 ( .A1(S_13_Rq3[1]), .A2(S_13_Rq2[3]), .ZN(
        S_13_G_CF_Out[6]) );
  XNOR2_X1 S_13_G_Inst_7__CF_Inst_U2 ( .A(S_13_G_Inst_7__CF_Inst_n3), .B(
        S_13_Rq3[0]), .ZN(S_13_G_CF_Out[7]) );
  NAND2_X1 S_13_G_Inst_7__CF_Inst_U1 ( .A1(S_13_Rq1[1]), .A2(S_13_Rq3[3]), 
        .ZN(S_13_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_13_G_Inst_8__CF_Inst_U1 ( .A1(S_13_Rq3[3]), .A2(S_13_Rq3[1]), .ZN(
        S_13_G_CF_Out[8]) );
  NOR2_X1 S_13_G_Inst_9__CF_Inst_U2 ( .A1(S_13_Rq1[3]), .A2(
        S_13_G_Inst_9__CF_Inst_n3), .ZN(S_13_G_CF_Out[9]) );
  INV_X1 S_13_G_Inst_9__CF_Inst_U1 ( .A(S_13_Rq1[2]), .ZN(
        S_13_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_13_G_Inst_10__CF_Inst_U2 ( .A1(S_13_Rq2[2]), .A2(
        S_13_G_Inst_10__CF_Inst_n3), .ZN(S_13_G_CF_Out[10]) );
  INV_X1 S_13_G_Inst_10__CF_Inst_U1 ( .A(S_13_Rq1[3]), .ZN(
        S_13_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_13_G_Inst_11__CF_Inst_U3 ( .A(S_13_Rq1[1]), .B(
        S_13_G_Inst_11__CF_Inst_n6), .ZN(S_13_G_CF_Out[11]) );
  NAND2_X1 S_13_G_Inst_11__CF_Inst_U2 ( .A1(S_13_Rq1[3]), .A2(
        S_13_G_Inst_11__CF_Inst_n5), .ZN(S_13_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_13_G_Inst_11__CF_Inst_U1 ( .A(S_13_Rq3[2]), .ZN(
        S_13_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_13_G_Inst_12__CF_Inst_U2 ( .A1(S_13_Rq2[3]), .A2(
        S_13_G_Inst_12__CF_Inst_n3), .ZN(S_13_G_CF_Out[12]) );
  INV_X1 S_13_G_Inst_12__CF_Inst_U1 ( .A(S_13_Rq1[2]), .ZN(
        S_13_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_13_G_Inst_13__CF_Inst_U1 ( .A1(S_13_Rq2[2]), .A2(S_13_Rq2[3]), 
        .ZN(S_13_G_CF_Out[13]) );
  XNOR2_X1 S_13_G_Inst_14__CF_Inst_U3 ( .A(S_13_Rq2[1]), .B(
        S_13_G_Inst_14__CF_Inst_n6), .ZN(S_13_G_CF_Out[14]) );
  NAND2_X1 S_13_G_Inst_14__CF_Inst_U2 ( .A1(S_13_Rq3[2]), .A2(
        S_13_G_Inst_14__CF_Inst_n5), .ZN(S_13_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_13_G_Inst_14__CF_Inst_U1 ( .A(S_13_Rq2[3]), .ZN(
        S_13_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_13_G_Inst_15__CF_Inst_U2 ( .A(S_13_G_Inst_15__CF_Inst_n3), .B(
        S_13_Rq3[1]), .ZN(S_13_G_CF_Out[15]) );
  NAND2_X1 S_13_G_Inst_15__CF_Inst_U1 ( .A1(S_13_Rq1[2]), .A2(S_13_Rq3[3]), 
        .ZN(S_13_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_13_G_Inst_16__CF_Inst_U1 ( .A1(S_13_Rq2[2]), .A2(S_13_Rq3[3]), 
        .ZN(S_13_G_CF_Out[16]) );
  NOR2_X1 S_13_G_Inst_17__CF_Inst_U2 ( .A1(S_13_Rq3[3]), .A2(
        S_13_G_Inst_17__CF_Inst_n3), .ZN(S_13_G_CF_Out[17]) );
  INV_X1 S_13_G_Inst_17__CF_Inst_U1 ( .A(S_13_Rq3[2]), .ZN(
        S_13_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_13_G_InstXOR_0__Compression1_U2 ( .A(
        S_13_G_InstXOR_0__Compression1_n3), .B(S_13_G_CF_Reg[2]), .ZN(
        S_13_G_out1[0]) );
  XNOR2_X1 S_13_G_InstXOR_0__Compression1_U1 ( .A(S_13_G_CF_Reg[0]), .B(
        S_13_G_CF_Reg[1]), .ZN(S_13_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_13_G_InstXOR_0__Compression2_U2 ( .A(
        S_13_G_InstXOR_0__Compression2_n3), .B(S_13_G_CF_Reg[5]), .ZN(
        SUB_OUT2[53]) );
  XNOR2_X1 S_13_G_InstXOR_0__Compression2_U1 ( .A(S_13_G_CF_Reg[3]), .B(
        S_13_G_CF_Reg[4]), .ZN(S_13_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_13_G_InstXOR_0__Compression3_U2 ( .A(
        S_13_G_InstXOR_0__Compression3_n3), .B(S_13_G_CF_Reg[8]), .ZN(
        SUB_OUT3[53]) );
  XNOR2_X1 S_13_G_InstXOR_0__Compression3_U1 ( .A(S_13_G_CF_Reg[6]), .B(
        S_13_G_CF_Reg[7]), .ZN(S_13_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_13_G_InstXOR_1__Compression1_U2 ( .A(
        S_13_G_InstXOR_1__Compression1_n3), .B(S_13_G_CF_Reg[11]), .ZN(
        S_13_G_out1[1]) );
  XNOR2_X1 S_13_G_InstXOR_1__Compression1_U1 ( .A(S_13_G_CF_Reg[9]), .B(
        S_13_G_CF_Reg[10]), .ZN(S_13_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_13_G_InstXOR_1__Compression2_U2 ( .A(
        S_13_G_InstXOR_1__Compression2_n3), .B(S_13_G_CF_Reg[14]), .ZN(
        SUB_OUT2[52]) );
  XNOR2_X1 S_13_G_InstXOR_1__Compression2_U1 ( .A(S_13_G_CF_Reg[12]), .B(
        S_13_G_CF_Reg[13]), .ZN(S_13_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_13_G_InstXOR_1__Compression3_U2 ( .A(
        S_13_G_InstXOR_1__Compression3_n3), .B(S_13_G_CF_Reg[17]), .ZN(
        SUB_OUT3[52]) );
  XNOR2_X1 S_13_G_InstXOR_1__Compression3_U1 ( .A(S_13_G_CF_Reg[15]), .B(
        S_13_G_CF_Reg[16]), .ZN(S_13_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_13_OutputAffine_U4 ( .A(S_13_G_out1[3]), .ZN(SUB_OUT1[55]) );
  INV_X1 S_13_OutputAffine_U3 ( .A(S_13_G_out1[2]), .ZN(SUB_OUT1[54]) );
  INV_X1 S_13_OutputAffine_U2 ( .A(S_13_G_out1[1]), .ZN(SUB_OUT1[52]) );
  INV_X1 S_13_OutputAffine_U1 ( .A(S_13_G_out1[0]), .ZN(SUB_OUT1[53]) );
  DFF_X1 S_14_Rq3_reg_0_ ( .D(S_14_q3[0]), .CK(CLK), .Q(S_14_Rq3[0]), .QN() );
  DFF_X1 S_14_Rq3_reg_1_ ( .D(S_14_q3[1]), .CK(CLK), .Q(S_14_Rq3[1]), .QN() );
  DFF_X1 S_14_Rq3_reg_2_ ( .D(S_14_q3[2]), .CK(CLK), .Q(S_14_Rq3[2]), .QN() );
  DFF_X1 S_14_Rq3_reg_3_ ( .D(S_14_q3[3]), .CK(CLK), .Q(S_14_Rq3[3]), .QN() );
  DFF_X1 S_14_Rq2_reg_0_ ( .D(S_14_q2[0]), .CK(CLK), .Q(S_14_Rq2[0]), .QN() );
  DFF_X1 S_14_Rq2_reg_1_ ( .D(S_14_q2[1]), .CK(CLK), .Q(S_14_Rq2[1]), .QN() );
  DFF_X1 S_14_Rq2_reg_2_ ( .D(S_14_q2[2]), .CK(CLK), .Q(S_14_Rq2[2]), .QN() );
  DFF_X1 S_14_Rq2_reg_3_ ( .D(S_14_q2[3]), .CK(CLK), .Q(S_14_Rq2[3]), .QN() );
  DFF_X1 S_14_Rq1_reg_0_ ( .D(S_14_q1[0]), .CK(CLK), .Q(S_14_Rq1[0]), .QN() );
  DFF_X1 S_14_Rq1_reg_1_ ( .D(S_14_q1[1]), .CK(CLK), .Q(S_14_Rq1[1]), .QN() );
  DFF_X1 S_14_Rq1_reg_2_ ( .D(S_14_q1[2]), .CK(CLK), .Q(S_14_Rq1[2]), .QN() );
  DFF_X1 S_14_Rq1_reg_3_ ( .D(S_14_q1[3]), .CK(CLK), .Q(S_14_Rq1[3]), .QN() );
  INV_X1 S_14_InputAffine_U4 ( .A(SUB_IN1[56]), .ZN(S_14_F_in1[0]) );
  INV_X1 S_14_InputAffine_U3 ( .A(SUB_IN1[58]), .ZN(S_14_F_in1[3]) );
  INV_X1 S_14_InputAffine_U2 ( .A(SUB_IN1[59]), .ZN(S_14_F_in1[1]) );
  INV_X1 S_14_InputAffine_U1 ( .A(SUB_IN1[57]), .ZN(S_14_F_in1[2]) );
  XNOR2_X1 S_14_F_U18 ( .A(S_14_F_n12), .B(FRESH[115]), .ZN(S_14_q3[3]) );
  XNOR2_X1 S_14_F_U17 ( .A(FRESH[114]), .B(S_14_F_q3[3]), .ZN(S_14_F_n12) );
  XNOR2_X1 S_14_F_U16 ( .A(S_14_F_n11), .B(FRESH[113]), .ZN(S_14_q3[2]) );
  XNOR2_X1 S_14_F_U15 ( .A(FRESH[112]), .B(S_14_F_q3[2]), .ZN(S_14_F_n11) );
  XOR2_X1 S_14_F_U14 ( .A(FRESH[115]), .B(S_14_F_q2[3]), .Z(S_14_q2[3]) );
  XOR2_X1 S_14_F_U13 ( .A(FRESH[113]), .B(S_14_F_q2[2]), .Z(S_14_q2[2]) );
  XOR2_X1 S_14_F_U12 ( .A(FRESH[114]), .B(S_14_F_q1[3]), .Z(S_14_q1[3]) );
  XOR2_X1 S_14_F_U11 ( .A(FRESH[112]), .B(S_14_F_q1[2]), .Z(S_14_q1[2]) );
  XNOR2_X1 S_14_F_U10 ( .A(S_14_F_n10), .B(FRESH[117]), .ZN(S_14_F_N5) );
  XNOR2_X1 S_14_F_U9 ( .A(S_14_F_in3[3]), .B(FRESH[116]), .ZN(S_14_F_n10) );
  XOR2_X1 S_14_F_U8 ( .A(FRESH[117]), .B(S_14_F_in2[3]), .Z(S_14_F_N4) );
  XOR2_X1 S_14_F_U7 ( .A(FRESH[116]), .B(S_14_F_in1[3]), .Z(S_14_F_N3) );
  XNOR2_X1 S_14_F_U6 ( .A(S_14_F_n9), .B(FRESH[119]), .ZN(S_14_F_N2) );
  XNOR2_X1 S_14_F_U5 ( .A(S_14_F_in3[2]), .B(FRESH[118]), .ZN(S_14_F_n9) );
  XOR2_X1 S_14_F_U4 ( .A(FRESH[119]), .B(S_14_F_in2[2]), .Z(S_14_F_N1) );
  XOR2_X1 S_14_F_U3 ( .A(FRESH[118]), .B(S_14_F_in1[2]), .Z(S_14_F_N0) );
  DFF_X1 S_14_F_CF_Reg_reg_0_ ( .D(S_14_F_CF_Out[0]), .CK(CLK), .Q(
        S_14_F_CF_Reg[0]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_1_ ( .D(S_14_F_CF_Out[1]), .CK(CLK), .Q(
        S_14_F_CF_Reg[1]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_2_ ( .D(S_14_F_CF_Out[2]), .CK(CLK), .Q(
        S_14_F_CF_Reg[2]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_3_ ( .D(S_14_F_CF_Out[3]), .CK(CLK), .Q(
        S_14_F_CF_Reg[3]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_4_ ( .D(S_14_F_CF_Out[4]), .CK(CLK), .Q(
        S_14_F_CF_Reg[4]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_5_ ( .D(S_14_F_CF_Out[5]), .CK(CLK), .Q(
        S_14_F_CF_Reg[5]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_6_ ( .D(S_14_F_CF_Out[6]), .CK(CLK), .Q(
        S_14_F_CF_Reg[6]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_7_ ( .D(S_14_F_CF_Out[7]), .CK(CLK), .Q(
        S_14_F_CF_Reg[7]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_8_ ( .D(S_14_F_CF_Out[8]), .CK(CLK), .Q(
        S_14_F_CF_Reg[8]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_9_ ( .D(S_14_F_CF_Out[9]), .CK(CLK), .Q(
        S_14_F_CF_Reg[9]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_10_ ( .D(S_14_F_CF_Out[10]), .CK(CLK), .Q(
        S_14_F_CF_Reg[10]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_11_ ( .D(S_14_F_CF_Out[11]), .CK(CLK), .Q(
        S_14_F_CF_Reg[11]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_12_ ( .D(S_14_F_CF_Out[12]), .CK(CLK), .Q(
        S_14_F_CF_Reg[12]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_13_ ( .D(S_14_F_CF_Out[13]), .CK(CLK), .Q(
        S_14_F_CF_Reg[13]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_14_ ( .D(S_14_F_CF_Out[14]), .CK(CLK), .Q(
        S_14_F_CF_Reg[14]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_15_ ( .D(S_14_F_CF_Out[15]), .CK(CLK), .Q(
        S_14_F_CF_Reg[15]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_16_ ( .D(S_14_F_CF_Out[16]), .CK(CLK), .Q(
        S_14_F_CF_Reg[16]), .QN() );
  DFF_X1 S_14_F_CF_Reg_reg_17_ ( .D(S_14_F_CF_Out[17]), .CK(CLK), .Q(
        S_14_F_CF_Reg[17]), .QN() );
  DFF_X1 S_14_F_out2_reg_0_ ( .D(S_14_F_N4), .CK(CLK), .Q(S_14_q2[0]), .QN()
         );
  DFF_X1 S_14_F_out2_reg_1_ ( .D(S_14_F_N1), .CK(CLK), .Q(S_14_q2[1]), .QN()
         );
  DFF_X1 S_14_F_out3_reg_0_ ( .D(S_14_F_N5), .CK(CLK), .Q(S_14_q3[0]), .QN()
         );
  DFF_X1 S_14_F_out3_reg_1_ ( .D(S_14_F_N2), .CK(CLK), .Q(S_14_q3[1]), .QN()
         );
  DFF_X1 S_14_F_out1_reg_0_ ( .D(S_14_F_N3), .CK(CLK), .Q(S_14_q1[0]), .QN()
         );
  DFF_X1 S_14_F_out1_reg_1_ ( .D(S_14_F_N0), .CK(CLK), .Q(S_14_q1[1]), .QN()
         );
  NOR2_X1 S_14_F_Inst_0__CF_Inst_U2 ( .A1(S_14_F_in1[2]), .A2(
        S_14_F_Inst_0__CF_Inst_n3), .ZN(S_14_F_CF_Out[0]) );
  INV_X1 S_14_F_Inst_0__CF_Inst_U1 ( .A(S_14_F_in1[3]), .ZN(
        S_14_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_14_F_Inst_1__CF_Inst_U2 ( .A(S_14_F_Inst_1__CF_Inst_n3), .B(
        S_14_F_in1[1]), .ZN(S_14_F_CF_Out[1]) );
  NAND2_X1 S_14_F_Inst_1__CF_Inst_U1 ( .A1(S_14_F_in2[2]), .A2(S_14_F_in1[3]), 
        .ZN(S_14_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_14_F_Inst_2__CF_Inst_U1 ( .A1(S_14_F_in1[3]), .A2(S_14_F_in3[2]), 
        .ZN(S_14_F_CF_Out[2]) );
  NOR2_X1 S_14_F_Inst_3__CF_Inst_U2 ( .A1(S_14_F_in2[3]), .A2(
        S_14_F_Inst_3__CF_Inst_n3), .ZN(S_14_F_CF_Out[3]) );
  INV_X1 S_14_F_Inst_3__CF_Inst_U1 ( .A(S_14_F_in1[2]), .ZN(
        S_14_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_14_F_Inst_4__CF_Inst_U2 ( .A(S_14_F_Inst_4__CF_Inst_n3), .B(
        S_14_F_in2[1]), .ZN(S_14_F_CF_Out[4]) );
  NAND2_X1 S_14_F_Inst_4__CF_Inst_U1 ( .A1(S_14_F_in2[2]), .A2(S_14_F_in2[3]), 
        .ZN(S_14_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_14_F_Inst_5__CF_Inst_U1 ( .A1(S_14_F_in3[2]), .A2(S_14_F_in2[3]), 
        .ZN(S_14_F_CF_Out[5]) );
  XNOR2_X1 S_14_F_Inst_6__CF_Inst_U2 ( .A(S_14_F_Inst_6__CF_Inst_n7), .B(
        S_14_F_in3[1]), .ZN(S_14_F_CF_Out[6]) );
  NOR2_X1 S_14_F_Inst_6__CF_Inst_U1 ( .A1(S_14_F_in1[2]), .A2(S_14_F_in3[3]), 
        .ZN(S_14_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_14_F_Inst_7__CF_Inst_U1 ( .A1(S_14_F_in2[2]), .A2(S_14_F_in3[3]), 
        .ZN(S_14_F_CF_Out[7]) );
  OR2_X1 S_14_F_Inst_8__CF_Inst_U1 ( .A1(S_14_F_in3[3]), .A2(S_14_F_in3[2]), 
        .ZN(S_14_F_CF_Out[8]) );
  NOR2_X1 S_14_F_Inst_9__CF_Inst_U2 ( .A1(S_14_F_in1[3]), .A2(
        S_14_F_Inst_9__CF_Inst_n3), .ZN(S_14_F_CF_Out[9]) );
  INV_X1 S_14_F_Inst_9__CF_Inst_U1 ( .A(S_14_F_in1[1]), .ZN(
        S_14_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_14_F_Inst_10__CF_Inst_U1 ( .A1(S_14_F_in2[1]), .A2(S_14_F_in1[3]), 
        .ZN(S_14_F_CF_Out[10]) );
  XNOR2_X1 S_14_F_Inst_11__CF_Inst_U2 ( .A(S_14_F_Inst_11__CF_Inst_n3), .B(
        S_14_F_in1[0]), .ZN(S_14_F_CF_Out[11]) );
  NAND2_X1 S_14_F_Inst_11__CF_Inst_U1 ( .A1(S_14_F_in3[1]), .A2(S_14_F_in1[3]), 
        .ZN(S_14_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_14_F_Inst_12__CF_Inst_U2 ( .A(S_14_F_Inst_12__CF_Inst_n3), .B(
        S_14_F_in2[0]), .ZN(S_14_F_CF_Out[12]) );
  NAND2_X1 S_14_F_Inst_12__CF_Inst_U1 ( .A1(S_14_F_in1[1]), .A2(S_14_F_in2[3]), 
        .ZN(S_14_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_14_F_Inst_13__CF_Inst_U2 ( .A1(S_14_F_in2[3]), .A2(
        S_14_F_Inst_13__CF_Inst_n3), .ZN(S_14_F_CF_Out[13]) );
  INV_X1 S_14_F_Inst_13__CF_Inst_U1 ( .A(S_14_F_in2[1]), .ZN(
        S_14_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_14_F_Inst_14__CF_Inst_U1 ( .A1(S_14_F_in3[1]), .A2(S_14_F_in2[3]), 
        .ZN(S_14_F_CF_Out[14]) );
  XNOR2_X1 S_14_F_Inst_15__CF_Inst_U2 ( .A(S_14_F_Inst_15__CF_Inst_n7), .B(
        S_14_F_in3[0]), .ZN(S_14_F_CF_Out[15]) );
  NOR2_X1 S_14_F_Inst_15__CF_Inst_U1 ( .A1(S_14_F_in1[1]), .A2(S_14_F_in3[3]), 
        .ZN(S_14_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_14_F_Inst_16__CF_Inst_U2 ( .A1(S_14_F_in3[3]), .A2(
        S_14_F_Inst_16__CF_Inst_n3), .ZN(S_14_F_CF_Out[16]) );
  INV_X1 S_14_F_Inst_16__CF_Inst_U1 ( .A(S_14_F_in2[1]), .ZN(
        S_14_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_14_F_Inst_17__CF_Inst_U2 ( .A1(S_14_F_in3[1]), .A2(
        S_14_F_Inst_17__CF_Inst_n3), .ZN(S_14_F_CF_Out[17]) );
  INV_X1 S_14_F_Inst_17__CF_Inst_U1 ( .A(S_14_F_in3[3]), .ZN(
        S_14_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_14_F_InstXOR_0__Compression1_U2 ( .A(
        S_14_F_InstXOR_0__Compression1_n3), .B(S_14_F_CF_Reg[2]), .ZN(
        S_14_F_q1[2]) );
  XNOR2_X1 S_14_F_InstXOR_0__Compression1_U1 ( .A(S_14_F_CF_Reg[0]), .B(
        S_14_F_CF_Reg[1]), .ZN(S_14_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_14_F_InstXOR_0__Compression2_U2 ( .A(
        S_14_F_InstXOR_0__Compression2_n3), .B(S_14_F_CF_Reg[5]), .ZN(
        S_14_F_q2[2]) );
  XNOR2_X1 S_14_F_InstXOR_0__Compression2_U1 ( .A(S_14_F_CF_Reg[3]), .B(
        S_14_F_CF_Reg[4]), .ZN(S_14_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_14_F_InstXOR_0__Compression3_U2 ( .A(
        S_14_F_InstXOR_0__Compression3_n3), .B(S_14_F_CF_Reg[8]), .ZN(
        S_14_F_q3[2]) );
  XNOR2_X1 S_14_F_InstXOR_0__Compression3_U1 ( .A(S_14_F_CF_Reg[6]), .B(
        S_14_F_CF_Reg[7]), .ZN(S_14_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_14_F_InstXOR_1__Compression1_U2 ( .A(
        S_14_F_InstXOR_1__Compression1_n3), .B(S_14_F_CF_Reg[11]), .ZN(
        S_14_F_q1[3]) );
  XNOR2_X1 S_14_F_InstXOR_1__Compression1_U1 ( .A(S_14_F_CF_Reg[9]), .B(
        S_14_F_CF_Reg[10]), .ZN(S_14_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_14_F_InstXOR_1__Compression2_U2 ( .A(
        S_14_F_InstXOR_1__Compression2_n3), .B(S_14_F_CF_Reg[14]), .ZN(
        S_14_F_q2[3]) );
  XNOR2_X1 S_14_F_InstXOR_1__Compression2_U1 ( .A(S_14_F_CF_Reg[12]), .B(
        S_14_F_CF_Reg[13]), .ZN(S_14_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_14_F_InstXOR_1__Compression3_U2 ( .A(
        S_14_F_InstXOR_1__Compression3_n3), .B(S_14_F_CF_Reg[17]), .ZN(
        S_14_F_q3[3]) );
  XNOR2_X1 S_14_F_InstXOR_1__Compression3_U1 ( .A(S_14_F_CF_Reg[15]), .B(
        S_14_F_CF_Reg[16]), .ZN(S_14_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_14_G_CF_Reg_reg_0_ ( .D(S_14_G_CF_Out[0]), .CK(CLK), .Q(
        S_14_G_CF_Reg[0]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_1_ ( .D(S_14_G_CF_Out[1]), .CK(CLK), .Q(
        S_14_G_CF_Reg[1]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_2_ ( .D(S_14_G_CF_Out[2]), .CK(CLK), .Q(
        S_14_G_CF_Reg[2]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_3_ ( .D(S_14_G_CF_Out[3]), .CK(CLK), .Q(
        S_14_G_CF_Reg[3]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_4_ ( .D(S_14_G_CF_Out[4]), .CK(CLK), .Q(
        S_14_G_CF_Reg[4]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_5_ ( .D(S_14_G_CF_Out[5]), .CK(CLK), .Q(
        S_14_G_CF_Reg[5]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_6_ ( .D(S_14_G_CF_Out[6]), .CK(CLK), .Q(
        S_14_G_CF_Reg[6]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_7_ ( .D(S_14_G_CF_Out[7]), .CK(CLK), .Q(
        S_14_G_CF_Reg[7]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_8_ ( .D(S_14_G_CF_Out[8]), .CK(CLK), .Q(
        S_14_G_CF_Reg[8]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_9_ ( .D(S_14_G_CF_Out[9]), .CK(CLK), .Q(
        S_14_G_CF_Reg[9]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_10_ ( .D(S_14_G_CF_Out[10]), .CK(CLK), .Q(
        S_14_G_CF_Reg[10]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_11_ ( .D(S_14_G_CF_Out[11]), .CK(CLK), .Q(
        S_14_G_CF_Reg[11]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_12_ ( .D(S_14_G_CF_Out[12]), .CK(CLK), .Q(
        S_14_G_CF_Reg[12]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_13_ ( .D(S_14_G_CF_Out[13]), .CK(CLK), .Q(
        S_14_G_CF_Reg[13]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_14_ ( .D(S_14_G_CF_Out[14]), .CK(CLK), .Q(
        S_14_G_CF_Reg[14]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_15_ ( .D(S_14_G_CF_Out[15]), .CK(CLK), .Q(
        S_14_G_CF_Reg[15]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_16_ ( .D(S_14_G_CF_Out[16]), .CK(CLK), .Q(
        S_14_G_CF_Reg[16]), .QN() );
  DFF_X1 S_14_G_CF_Reg_reg_17_ ( .D(S_14_G_CF_Out[17]), .CK(CLK), .Q(
        S_14_G_CF_Reg[17]), .QN() );
  DFF_X1 S_14_G_out1_reg_2_ ( .D(S_14_Rq1[2]), .CK(CLK), .Q(S_14_G_out1[2]), 
        .QN() );
  DFF_X1 S_14_G_out1_reg_3_ ( .D(S_14_Rq1[3]), .CK(CLK), .Q(S_14_G_out1[3]), 
        .QN() );
  DFF_X1 S_14_G_out2_reg_2_ ( .D(S_14_Rq2[2]), .CK(CLK), .Q(SUB_OUT2[58]), 
        .QN() );
  DFF_X1 S_14_G_out2_reg_3_ ( .D(S_14_Rq2[3]), .CK(CLK), .Q(SUB_OUT2[59]), 
        .QN() );
  DFF_X1 S_14_G_out3_reg_2_ ( .D(S_14_Rq3[2]), .CK(CLK), .Q(SUB_OUT3[58]), 
        .QN() );
  DFF_X1 S_14_G_out3_reg_3_ ( .D(S_14_Rq3[3]), .CK(CLK), .Q(SUB_OUT3[59]), 
        .QN() );
  AND2_X1 S_14_G_Inst_0__CF_Inst_U1 ( .A1(S_14_Rq1[1]), .A2(S_14_Rq1[3]), .ZN(
        S_14_G_CF_Out[0]) );
  NOR2_X1 S_14_G_Inst_1__CF_Inst_U2 ( .A1(S_14_Rq1[3]), .A2(
        S_14_G_Inst_1__CF_Inst_n3), .ZN(S_14_G_CF_Out[1]) );
  INV_X1 S_14_G_Inst_1__CF_Inst_U1 ( .A(S_14_Rq2[1]), .ZN(
        S_14_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_14_G_Inst_2__CF_Inst_U2 ( .A(S_14_G_Inst_2__CF_Inst_n3), .B(
        S_14_Rq2[0]), .ZN(S_14_G_CF_Out[2]) );
  NAND2_X1 S_14_G_Inst_2__CF_Inst_U1 ( .A1(S_14_Rq1[1]), .A2(S_14_Rq2[3]), 
        .ZN(S_14_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_14_G_Inst_3__CF_Inst_U3 ( .A(S_14_Rq1[0]), .B(
        S_14_G_Inst_3__CF_Inst_n6), .ZN(S_14_G_CF_Out[3]) );
  NAND2_X1 S_14_G_Inst_3__CF_Inst_U2 ( .A1(S_14_Rq3[1]), .A2(
        S_14_G_Inst_3__CF_Inst_n5), .ZN(S_14_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_14_G_Inst_3__CF_Inst_U1 ( .A(S_14_Rq1[3]), .ZN(
        S_14_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_14_G_Inst_4__CF_Inst_U1 ( .A1(S_14_Rq2[1]), .A2(S_14_Rq2[3]), .ZN(
        S_14_G_CF_Out[4]) );
  OR2_X1 S_14_G_Inst_5__CF_Inst_U1 ( .A1(S_14_Rq3[3]), .A2(S_14_Rq2[1]), .ZN(
        S_14_G_CF_Out[5]) );
  AND2_X1 S_14_G_Inst_6__CF_Inst_U1 ( .A1(S_14_Rq3[1]), .A2(S_14_Rq2[3]), .ZN(
        S_14_G_CF_Out[6]) );
  XNOR2_X1 S_14_G_Inst_7__CF_Inst_U2 ( .A(S_14_G_Inst_7__CF_Inst_n3), .B(
        S_14_Rq3[0]), .ZN(S_14_G_CF_Out[7]) );
  NAND2_X1 S_14_G_Inst_7__CF_Inst_U1 ( .A1(S_14_Rq1[1]), .A2(S_14_Rq3[3]), 
        .ZN(S_14_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_14_G_Inst_8__CF_Inst_U1 ( .A1(S_14_Rq3[3]), .A2(S_14_Rq3[1]), .ZN(
        S_14_G_CF_Out[8]) );
  NOR2_X1 S_14_G_Inst_9__CF_Inst_U2 ( .A1(S_14_Rq1[3]), .A2(
        S_14_G_Inst_9__CF_Inst_n3), .ZN(S_14_G_CF_Out[9]) );
  INV_X1 S_14_G_Inst_9__CF_Inst_U1 ( .A(S_14_Rq1[2]), .ZN(
        S_14_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_14_G_Inst_10__CF_Inst_U2 ( .A1(S_14_Rq2[2]), .A2(
        S_14_G_Inst_10__CF_Inst_n3), .ZN(S_14_G_CF_Out[10]) );
  INV_X1 S_14_G_Inst_10__CF_Inst_U1 ( .A(S_14_Rq1[3]), .ZN(
        S_14_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_14_G_Inst_11__CF_Inst_U3 ( .A(S_14_Rq1[1]), .B(
        S_14_G_Inst_11__CF_Inst_n6), .ZN(S_14_G_CF_Out[11]) );
  NAND2_X1 S_14_G_Inst_11__CF_Inst_U2 ( .A1(S_14_Rq1[3]), .A2(
        S_14_G_Inst_11__CF_Inst_n5), .ZN(S_14_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_14_G_Inst_11__CF_Inst_U1 ( .A(S_14_Rq3[2]), .ZN(
        S_14_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_14_G_Inst_12__CF_Inst_U2 ( .A1(S_14_Rq2[3]), .A2(
        S_14_G_Inst_12__CF_Inst_n3), .ZN(S_14_G_CF_Out[12]) );
  INV_X1 S_14_G_Inst_12__CF_Inst_U1 ( .A(S_14_Rq1[2]), .ZN(
        S_14_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_14_G_Inst_13__CF_Inst_U1 ( .A1(S_14_Rq2[2]), .A2(S_14_Rq2[3]), 
        .ZN(S_14_G_CF_Out[13]) );
  XNOR2_X1 S_14_G_Inst_14__CF_Inst_U3 ( .A(S_14_Rq2[1]), .B(
        S_14_G_Inst_14__CF_Inst_n6), .ZN(S_14_G_CF_Out[14]) );
  NAND2_X1 S_14_G_Inst_14__CF_Inst_U2 ( .A1(S_14_Rq3[2]), .A2(
        S_14_G_Inst_14__CF_Inst_n5), .ZN(S_14_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_14_G_Inst_14__CF_Inst_U1 ( .A(S_14_Rq2[3]), .ZN(
        S_14_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_14_G_Inst_15__CF_Inst_U2 ( .A(S_14_G_Inst_15__CF_Inst_n3), .B(
        S_14_Rq3[1]), .ZN(S_14_G_CF_Out[15]) );
  NAND2_X1 S_14_G_Inst_15__CF_Inst_U1 ( .A1(S_14_Rq1[2]), .A2(S_14_Rq3[3]), 
        .ZN(S_14_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_14_G_Inst_16__CF_Inst_U1 ( .A1(S_14_Rq2[2]), .A2(S_14_Rq3[3]), 
        .ZN(S_14_G_CF_Out[16]) );
  NOR2_X1 S_14_G_Inst_17__CF_Inst_U2 ( .A1(S_14_Rq3[3]), .A2(
        S_14_G_Inst_17__CF_Inst_n3), .ZN(S_14_G_CF_Out[17]) );
  INV_X1 S_14_G_Inst_17__CF_Inst_U1 ( .A(S_14_Rq3[2]), .ZN(
        S_14_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_14_G_InstXOR_0__Compression1_U2 ( .A(
        S_14_G_InstXOR_0__Compression1_n3), .B(S_14_G_CF_Reg[2]), .ZN(
        S_14_G_out1[0]) );
  XNOR2_X1 S_14_G_InstXOR_0__Compression1_U1 ( .A(S_14_G_CF_Reg[0]), .B(
        S_14_G_CF_Reg[1]), .ZN(S_14_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_14_G_InstXOR_0__Compression2_U2 ( .A(
        S_14_G_InstXOR_0__Compression2_n3), .B(S_14_G_CF_Reg[5]), .ZN(
        SUB_OUT2[57]) );
  XNOR2_X1 S_14_G_InstXOR_0__Compression2_U1 ( .A(S_14_G_CF_Reg[3]), .B(
        S_14_G_CF_Reg[4]), .ZN(S_14_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_14_G_InstXOR_0__Compression3_U2 ( .A(
        S_14_G_InstXOR_0__Compression3_n3), .B(S_14_G_CF_Reg[8]), .ZN(
        SUB_OUT3[57]) );
  XNOR2_X1 S_14_G_InstXOR_0__Compression3_U1 ( .A(S_14_G_CF_Reg[6]), .B(
        S_14_G_CF_Reg[7]), .ZN(S_14_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_14_G_InstXOR_1__Compression1_U2 ( .A(
        S_14_G_InstXOR_1__Compression1_n3), .B(S_14_G_CF_Reg[11]), .ZN(
        S_14_G_out1[1]) );
  XNOR2_X1 S_14_G_InstXOR_1__Compression1_U1 ( .A(S_14_G_CF_Reg[9]), .B(
        S_14_G_CF_Reg[10]), .ZN(S_14_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_14_G_InstXOR_1__Compression2_U2 ( .A(
        S_14_G_InstXOR_1__Compression2_n3), .B(S_14_G_CF_Reg[14]), .ZN(
        SUB_OUT2[56]) );
  XNOR2_X1 S_14_G_InstXOR_1__Compression2_U1 ( .A(S_14_G_CF_Reg[12]), .B(
        S_14_G_CF_Reg[13]), .ZN(S_14_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_14_G_InstXOR_1__Compression3_U2 ( .A(
        S_14_G_InstXOR_1__Compression3_n3), .B(S_14_G_CF_Reg[17]), .ZN(
        SUB_OUT3[56]) );
  XNOR2_X1 S_14_G_InstXOR_1__Compression3_U1 ( .A(S_14_G_CF_Reg[15]), .B(
        S_14_G_CF_Reg[16]), .ZN(S_14_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_14_OutputAffine_U4 ( .A(S_14_G_out1[3]), .ZN(SUB_OUT1[59]) );
  INV_X1 S_14_OutputAffine_U3 ( .A(S_14_G_out1[2]), .ZN(SUB_OUT1[58]) );
  INV_X1 S_14_OutputAffine_U2 ( .A(S_14_G_out1[1]), .ZN(SUB_OUT1[56]) );
  INV_X1 S_14_OutputAffine_U1 ( .A(S_14_G_out1[0]), .ZN(SUB_OUT1[57]) );
  DFF_X1 S_15_Rq3_reg_0_ ( .D(S_15_q3[0]), .CK(CLK), .Q(S_15_Rq3[0]), .QN() );
  DFF_X1 S_15_Rq3_reg_1_ ( .D(S_15_q3[1]), .CK(CLK), .Q(S_15_Rq3[1]), .QN() );
  DFF_X1 S_15_Rq3_reg_2_ ( .D(S_15_q3[2]), .CK(CLK), .Q(S_15_Rq3[2]), .QN() );
  DFF_X1 S_15_Rq3_reg_3_ ( .D(S_15_q3[3]), .CK(CLK), .Q(S_15_Rq3[3]), .QN() );
  DFF_X1 S_15_Rq2_reg_0_ ( .D(S_15_q2[0]), .CK(CLK), .Q(S_15_Rq2[0]), .QN() );
  DFF_X1 S_15_Rq2_reg_1_ ( .D(S_15_q2[1]), .CK(CLK), .Q(S_15_Rq2[1]), .QN() );
  DFF_X1 S_15_Rq2_reg_2_ ( .D(S_15_q2[2]), .CK(CLK), .Q(S_15_Rq2[2]), .QN() );
  DFF_X1 S_15_Rq2_reg_3_ ( .D(S_15_q2[3]), .CK(CLK), .Q(S_15_Rq2[3]), .QN() );
  DFF_X1 S_15_Rq1_reg_0_ ( .D(S_15_q1[0]), .CK(CLK), .Q(S_15_Rq1[0]), .QN() );
  DFF_X1 S_15_Rq1_reg_1_ ( .D(S_15_q1[1]), .CK(CLK), .Q(S_15_Rq1[1]), .QN() );
  DFF_X1 S_15_Rq1_reg_2_ ( .D(S_15_q1[2]), .CK(CLK), .Q(S_15_Rq1[2]), .QN() );
  DFF_X1 S_15_Rq1_reg_3_ ( .D(S_15_q1[3]), .CK(CLK), .Q(S_15_Rq1[3]), .QN() );
  INV_X1 S_15_InputAffine_U4 ( .A(SUB_IN1[60]), .ZN(S_15_F_in1[0]) );
  INV_X1 S_15_InputAffine_U3 ( .A(SUB_IN1[62]), .ZN(S_15_F_in1[3]) );
  INV_X1 S_15_InputAffine_U2 ( .A(SUB_IN1[63]), .ZN(S_15_F_in1[1]) );
  INV_X1 S_15_InputAffine_U1 ( .A(SUB_IN1[61]), .ZN(S_15_F_in1[2]) );
  XNOR2_X1 S_15_F_U18 ( .A(S_15_F_n12), .B(FRESH[123]), .ZN(S_15_q3[3]) );
  XNOR2_X1 S_15_F_U17 ( .A(FRESH[122]), .B(S_15_F_q3[3]), .ZN(S_15_F_n12) );
  XNOR2_X1 S_15_F_U16 ( .A(S_15_F_n11), .B(FRESH[121]), .ZN(S_15_q3[2]) );
  XNOR2_X1 S_15_F_U15 ( .A(FRESH[120]), .B(S_15_F_q3[2]), .ZN(S_15_F_n11) );
  XOR2_X1 S_15_F_U14 ( .A(FRESH[123]), .B(S_15_F_q2[3]), .Z(S_15_q2[3]) );
  XOR2_X1 S_15_F_U13 ( .A(FRESH[121]), .B(S_15_F_q2[2]), .Z(S_15_q2[2]) );
  XOR2_X1 S_15_F_U12 ( .A(FRESH[122]), .B(S_15_F_q1[3]), .Z(S_15_q1[3]) );
  XOR2_X1 S_15_F_U11 ( .A(FRESH[120]), .B(S_15_F_q1[2]), .Z(S_15_q1[2]) );
  XNOR2_X1 S_15_F_U10 ( .A(S_15_F_n10), .B(FRESH[125]), .ZN(S_15_F_N5) );
  XNOR2_X1 S_15_F_U9 ( .A(S_15_F_in3[3]), .B(FRESH[124]), .ZN(S_15_F_n10) );
  XOR2_X1 S_15_F_U8 ( .A(FRESH[125]), .B(S_15_F_in2[3]), .Z(S_15_F_N4) );
  XOR2_X1 S_15_F_U7 ( .A(FRESH[124]), .B(S_15_F_in1[3]), .Z(S_15_F_N3) );
  XNOR2_X1 S_15_F_U6 ( .A(S_15_F_n9), .B(FRESH[127]), .ZN(S_15_F_N2) );
  XNOR2_X1 S_15_F_U5 ( .A(S_15_F_in3[2]), .B(FRESH[126]), .ZN(S_15_F_n9) );
  XOR2_X1 S_15_F_U4 ( .A(FRESH[127]), .B(S_15_F_in2[2]), .Z(S_15_F_N1) );
  XOR2_X1 S_15_F_U3 ( .A(FRESH[126]), .B(S_15_F_in1[2]), .Z(S_15_F_N0) );
  DFF_X1 S_15_F_CF_Reg_reg_0_ ( .D(S_15_F_CF_Out[0]), .CK(CLK), .Q(
        S_15_F_CF_Reg[0]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_1_ ( .D(S_15_F_CF_Out[1]), .CK(CLK), .Q(
        S_15_F_CF_Reg[1]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_2_ ( .D(S_15_F_CF_Out[2]), .CK(CLK), .Q(
        S_15_F_CF_Reg[2]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_3_ ( .D(S_15_F_CF_Out[3]), .CK(CLK), .Q(
        S_15_F_CF_Reg[3]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_4_ ( .D(S_15_F_CF_Out[4]), .CK(CLK), .Q(
        S_15_F_CF_Reg[4]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_5_ ( .D(S_15_F_CF_Out[5]), .CK(CLK), .Q(
        S_15_F_CF_Reg[5]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_6_ ( .D(S_15_F_CF_Out[6]), .CK(CLK), .Q(
        S_15_F_CF_Reg[6]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_7_ ( .D(S_15_F_CF_Out[7]), .CK(CLK), .Q(
        S_15_F_CF_Reg[7]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_8_ ( .D(S_15_F_CF_Out[8]), .CK(CLK), .Q(
        S_15_F_CF_Reg[8]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_9_ ( .D(S_15_F_CF_Out[9]), .CK(CLK), .Q(
        S_15_F_CF_Reg[9]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_10_ ( .D(S_15_F_CF_Out[10]), .CK(CLK), .Q(
        S_15_F_CF_Reg[10]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_11_ ( .D(S_15_F_CF_Out[11]), .CK(CLK), .Q(
        S_15_F_CF_Reg[11]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_12_ ( .D(S_15_F_CF_Out[12]), .CK(CLK), .Q(
        S_15_F_CF_Reg[12]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_13_ ( .D(S_15_F_CF_Out[13]), .CK(CLK), .Q(
        S_15_F_CF_Reg[13]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_14_ ( .D(S_15_F_CF_Out[14]), .CK(CLK), .Q(
        S_15_F_CF_Reg[14]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_15_ ( .D(S_15_F_CF_Out[15]), .CK(CLK), .Q(
        S_15_F_CF_Reg[15]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_16_ ( .D(S_15_F_CF_Out[16]), .CK(CLK), .Q(
        S_15_F_CF_Reg[16]), .QN() );
  DFF_X1 S_15_F_CF_Reg_reg_17_ ( .D(S_15_F_CF_Out[17]), .CK(CLK), .Q(
        S_15_F_CF_Reg[17]), .QN() );
  DFF_X1 S_15_F_out2_reg_0_ ( .D(S_15_F_N4), .CK(CLK), .Q(S_15_q2[0]), .QN()
         );
  DFF_X1 S_15_F_out2_reg_1_ ( .D(S_15_F_N1), .CK(CLK), .Q(S_15_q2[1]), .QN()
         );
  DFF_X1 S_15_F_out3_reg_0_ ( .D(S_15_F_N5), .CK(CLK), .Q(S_15_q3[0]), .QN()
         );
  DFF_X1 S_15_F_out3_reg_1_ ( .D(S_15_F_N2), .CK(CLK), .Q(S_15_q3[1]), .QN()
         );
  DFF_X1 S_15_F_out1_reg_0_ ( .D(S_15_F_N3), .CK(CLK), .Q(S_15_q1[0]), .QN()
         );
  DFF_X1 S_15_F_out1_reg_1_ ( .D(S_15_F_N0), .CK(CLK), .Q(S_15_q1[1]), .QN()
         );
  NOR2_X1 S_15_F_Inst_0__CF_Inst_U2 ( .A1(S_15_F_in1[2]), .A2(
        S_15_F_Inst_0__CF_Inst_n3), .ZN(S_15_F_CF_Out[0]) );
  INV_X1 S_15_F_Inst_0__CF_Inst_U1 ( .A(S_15_F_in1[3]), .ZN(
        S_15_F_Inst_0__CF_Inst_n3) );
  XNOR2_X1 S_15_F_Inst_1__CF_Inst_U2 ( .A(S_15_F_Inst_1__CF_Inst_n3), .B(
        S_15_F_in1[1]), .ZN(S_15_F_CF_Out[1]) );
  NAND2_X1 S_15_F_Inst_1__CF_Inst_U1 ( .A1(S_15_F_in2[2]), .A2(S_15_F_in1[3]), 
        .ZN(S_15_F_Inst_1__CF_Inst_n3) );
  OR2_X1 S_15_F_Inst_2__CF_Inst_U1 ( .A1(S_15_F_in1[3]), .A2(S_15_F_in3[2]), 
        .ZN(S_15_F_CF_Out[2]) );
  NOR2_X1 S_15_F_Inst_3__CF_Inst_U2 ( .A1(S_15_F_in2[3]), .A2(
        S_15_F_Inst_3__CF_Inst_n3), .ZN(S_15_F_CF_Out[3]) );
  INV_X1 S_15_F_Inst_3__CF_Inst_U1 ( .A(S_15_F_in1[2]), .ZN(
        S_15_F_Inst_3__CF_Inst_n3) );
  XNOR2_X1 S_15_F_Inst_4__CF_Inst_U2 ( .A(S_15_F_Inst_4__CF_Inst_n3), .B(
        S_15_F_in2[1]), .ZN(S_15_F_CF_Out[4]) );
  NAND2_X1 S_15_F_Inst_4__CF_Inst_U1 ( .A1(S_15_F_in2[2]), .A2(S_15_F_in2[3]), 
        .ZN(S_15_F_Inst_4__CF_Inst_n3) );
  AND2_X1 S_15_F_Inst_5__CF_Inst_U1 ( .A1(S_15_F_in3[2]), .A2(S_15_F_in2[3]), 
        .ZN(S_15_F_CF_Out[5]) );
  XNOR2_X1 S_15_F_Inst_6__CF_Inst_U2 ( .A(S_15_F_Inst_6__CF_Inst_n7), .B(
        S_15_F_in3[1]), .ZN(S_15_F_CF_Out[6]) );
  NOR2_X1 S_15_F_Inst_6__CF_Inst_U1 ( .A1(S_15_F_in1[2]), .A2(S_15_F_in3[3]), 
        .ZN(S_15_F_Inst_6__CF_Inst_n7) );
  AND2_X1 S_15_F_Inst_7__CF_Inst_U1 ( .A1(S_15_F_in2[2]), .A2(S_15_F_in3[3]), 
        .ZN(S_15_F_CF_Out[7]) );
  OR2_X1 S_15_F_Inst_8__CF_Inst_U1 ( .A1(S_15_F_in3[3]), .A2(S_15_F_in3[2]), 
        .ZN(S_15_F_CF_Out[8]) );
  NOR2_X1 S_15_F_Inst_9__CF_Inst_U2 ( .A1(S_15_F_in1[3]), .A2(
        S_15_F_Inst_9__CF_Inst_n3), .ZN(S_15_F_CF_Out[9]) );
  INV_X1 S_15_F_Inst_9__CF_Inst_U1 ( .A(S_15_F_in1[1]), .ZN(
        S_15_F_Inst_9__CF_Inst_n3) );
  AND2_X1 S_15_F_Inst_10__CF_Inst_U1 ( .A1(S_15_F_in2[1]), .A2(S_15_F_in1[3]), 
        .ZN(S_15_F_CF_Out[10]) );
  XNOR2_X1 S_15_F_Inst_11__CF_Inst_U2 ( .A(S_15_F_Inst_11__CF_Inst_n3), .B(
        S_15_F_in1[0]), .ZN(S_15_F_CF_Out[11]) );
  NAND2_X1 S_15_F_Inst_11__CF_Inst_U1 ( .A1(S_15_F_in3[1]), .A2(S_15_F_in1[3]), 
        .ZN(S_15_F_Inst_11__CF_Inst_n3) );
  XNOR2_X1 S_15_F_Inst_12__CF_Inst_U2 ( .A(S_15_F_Inst_12__CF_Inst_n3), .B(
        S_15_F_in2[0]), .ZN(S_15_F_CF_Out[12]) );
  NAND2_X1 S_15_F_Inst_12__CF_Inst_U1 ( .A1(S_15_F_in1[1]), .A2(S_15_F_in2[3]), 
        .ZN(S_15_F_Inst_12__CF_Inst_n3) );
  NOR2_X1 S_15_F_Inst_13__CF_Inst_U2 ( .A1(S_15_F_in2[3]), .A2(
        S_15_F_Inst_13__CF_Inst_n3), .ZN(S_15_F_CF_Out[13]) );
  INV_X1 S_15_F_Inst_13__CF_Inst_U1 ( .A(S_15_F_in2[1]), .ZN(
        S_15_F_Inst_13__CF_Inst_n3) );
  AND2_X1 S_15_F_Inst_14__CF_Inst_U1 ( .A1(S_15_F_in3[1]), .A2(S_15_F_in2[3]), 
        .ZN(S_15_F_CF_Out[14]) );
  XNOR2_X1 S_15_F_Inst_15__CF_Inst_U2 ( .A(S_15_F_Inst_15__CF_Inst_n7), .B(
        S_15_F_in3[0]), .ZN(S_15_F_CF_Out[15]) );
  NOR2_X1 S_15_F_Inst_15__CF_Inst_U1 ( .A1(S_15_F_in1[1]), .A2(S_15_F_in3[3]), 
        .ZN(S_15_F_Inst_15__CF_Inst_n7) );
  NOR2_X1 S_15_F_Inst_16__CF_Inst_U2 ( .A1(S_15_F_in3[3]), .A2(
        S_15_F_Inst_16__CF_Inst_n3), .ZN(S_15_F_CF_Out[16]) );
  INV_X1 S_15_F_Inst_16__CF_Inst_U1 ( .A(S_15_F_in2[1]), .ZN(
        S_15_F_Inst_16__CF_Inst_n3) );
  NOR2_X1 S_15_F_Inst_17__CF_Inst_U2 ( .A1(S_15_F_in3[1]), .A2(
        S_15_F_Inst_17__CF_Inst_n3), .ZN(S_15_F_CF_Out[17]) );
  INV_X1 S_15_F_Inst_17__CF_Inst_U1 ( .A(S_15_F_in3[3]), .ZN(
        S_15_F_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_15_F_InstXOR_0__Compression1_U2 ( .A(
        S_15_F_InstXOR_0__Compression1_n3), .B(S_15_F_CF_Reg[2]), .ZN(
        S_15_F_q1[2]) );
  XNOR2_X1 S_15_F_InstXOR_0__Compression1_U1 ( .A(S_15_F_CF_Reg[0]), .B(
        S_15_F_CF_Reg[1]), .ZN(S_15_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_15_F_InstXOR_0__Compression2_U2 ( .A(
        S_15_F_InstXOR_0__Compression2_n3), .B(S_15_F_CF_Reg[5]), .ZN(
        S_15_F_q2[2]) );
  XNOR2_X1 S_15_F_InstXOR_0__Compression2_U1 ( .A(S_15_F_CF_Reg[3]), .B(
        S_15_F_CF_Reg[4]), .ZN(S_15_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_15_F_InstXOR_0__Compression3_U2 ( .A(
        S_15_F_InstXOR_0__Compression3_n3), .B(S_15_F_CF_Reg[8]), .ZN(
        S_15_F_q3[2]) );
  XNOR2_X1 S_15_F_InstXOR_0__Compression3_U1 ( .A(S_15_F_CF_Reg[6]), .B(
        S_15_F_CF_Reg[7]), .ZN(S_15_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_15_F_InstXOR_1__Compression1_U2 ( .A(
        S_15_F_InstXOR_1__Compression1_n3), .B(S_15_F_CF_Reg[11]), .ZN(
        S_15_F_q1[3]) );
  XNOR2_X1 S_15_F_InstXOR_1__Compression1_U1 ( .A(S_15_F_CF_Reg[9]), .B(
        S_15_F_CF_Reg[10]), .ZN(S_15_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_15_F_InstXOR_1__Compression2_U2 ( .A(
        S_15_F_InstXOR_1__Compression2_n3), .B(S_15_F_CF_Reg[14]), .ZN(
        S_15_F_q2[3]) );
  XNOR2_X1 S_15_F_InstXOR_1__Compression2_U1 ( .A(S_15_F_CF_Reg[12]), .B(
        S_15_F_CF_Reg[13]), .ZN(S_15_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_15_F_InstXOR_1__Compression3_U2 ( .A(
        S_15_F_InstXOR_1__Compression3_n3), .B(S_15_F_CF_Reg[17]), .ZN(
        S_15_F_q3[3]) );
  XNOR2_X1 S_15_F_InstXOR_1__Compression3_U1 ( .A(S_15_F_CF_Reg[15]), .B(
        S_15_F_CF_Reg[16]), .ZN(S_15_F_InstXOR_1__Compression3_n3) );
  DFF_X1 S_15_G_CF_Reg_reg_0_ ( .D(S_15_G_CF_Out[0]), .CK(CLK), .Q(
        S_15_G_CF_Reg[0]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_1_ ( .D(S_15_G_CF_Out[1]), .CK(CLK), .Q(
        S_15_G_CF_Reg[1]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_2_ ( .D(S_15_G_CF_Out[2]), .CK(CLK), .Q(
        S_15_G_CF_Reg[2]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_3_ ( .D(S_15_G_CF_Out[3]), .CK(CLK), .Q(
        S_15_G_CF_Reg[3]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_4_ ( .D(S_15_G_CF_Out[4]), .CK(CLK), .Q(
        S_15_G_CF_Reg[4]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_5_ ( .D(S_15_G_CF_Out[5]), .CK(CLK), .Q(
        S_15_G_CF_Reg[5]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_6_ ( .D(S_15_G_CF_Out[6]), .CK(CLK), .Q(
        S_15_G_CF_Reg[6]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_7_ ( .D(S_15_G_CF_Out[7]), .CK(CLK), .Q(
        S_15_G_CF_Reg[7]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_8_ ( .D(S_15_G_CF_Out[8]), .CK(CLK), .Q(
        S_15_G_CF_Reg[8]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_9_ ( .D(S_15_G_CF_Out[9]), .CK(CLK), .Q(
        S_15_G_CF_Reg[9]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_10_ ( .D(S_15_G_CF_Out[10]), .CK(CLK), .Q(
        S_15_G_CF_Reg[10]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_11_ ( .D(S_15_G_CF_Out[11]), .CK(CLK), .Q(
        S_15_G_CF_Reg[11]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_12_ ( .D(S_15_G_CF_Out[12]), .CK(CLK), .Q(
        S_15_G_CF_Reg[12]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_13_ ( .D(S_15_G_CF_Out[13]), .CK(CLK), .Q(
        S_15_G_CF_Reg[13]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_14_ ( .D(S_15_G_CF_Out[14]), .CK(CLK), .Q(
        S_15_G_CF_Reg[14]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_15_ ( .D(S_15_G_CF_Out[15]), .CK(CLK), .Q(
        S_15_G_CF_Reg[15]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_16_ ( .D(S_15_G_CF_Out[16]), .CK(CLK), .Q(
        S_15_G_CF_Reg[16]), .QN() );
  DFF_X1 S_15_G_CF_Reg_reg_17_ ( .D(S_15_G_CF_Out[17]), .CK(CLK), .Q(
        S_15_G_CF_Reg[17]), .QN() );
  DFF_X1 S_15_G_out1_reg_2_ ( .D(S_15_Rq1[2]), .CK(CLK), .Q(S_15_G_out1[2]), 
        .QN() );
  DFF_X1 S_15_G_out1_reg_3_ ( .D(S_15_Rq1[3]), .CK(CLK), .Q(S_15_G_out1[3]), 
        .QN() );
  DFF_X1 S_15_G_out2_reg_2_ ( .D(S_15_Rq2[2]), .CK(CLK), .Q(SUB_OUT2[62]), 
        .QN() );
  DFF_X1 S_15_G_out2_reg_3_ ( .D(S_15_Rq2[3]), .CK(CLK), .Q(SUB_OUT2[63]), 
        .QN() );
  DFF_X1 S_15_G_out3_reg_2_ ( .D(S_15_Rq3[2]), .CK(CLK), .Q(SUB_OUT3[62]), 
        .QN() );
  DFF_X1 S_15_G_out3_reg_3_ ( .D(S_15_Rq3[3]), .CK(CLK), .Q(SUB_OUT3[63]), 
        .QN() );
  AND2_X1 S_15_G_Inst_0__CF_Inst_U1 ( .A1(S_15_Rq1[1]), .A2(S_15_Rq1[3]), .ZN(
        S_15_G_CF_Out[0]) );
  NOR2_X1 S_15_G_Inst_1__CF_Inst_U2 ( .A1(S_15_Rq1[3]), .A2(
        S_15_G_Inst_1__CF_Inst_n3), .ZN(S_15_G_CF_Out[1]) );
  INV_X1 S_15_G_Inst_1__CF_Inst_U1 ( .A(S_15_Rq2[1]), .ZN(
        S_15_G_Inst_1__CF_Inst_n3) );
  XNOR2_X1 S_15_G_Inst_2__CF_Inst_U2 ( .A(S_15_G_Inst_2__CF_Inst_n3), .B(
        S_15_Rq2[0]), .ZN(S_15_G_CF_Out[2]) );
  NAND2_X1 S_15_G_Inst_2__CF_Inst_U1 ( .A1(S_15_Rq1[1]), .A2(S_15_Rq2[3]), 
        .ZN(S_15_G_Inst_2__CF_Inst_n3) );
  XNOR2_X1 S_15_G_Inst_3__CF_Inst_U3 ( .A(S_15_Rq1[0]), .B(
        S_15_G_Inst_3__CF_Inst_n6), .ZN(S_15_G_CF_Out[3]) );
  NAND2_X1 S_15_G_Inst_3__CF_Inst_U2 ( .A1(S_15_Rq3[1]), .A2(
        S_15_G_Inst_3__CF_Inst_n5), .ZN(S_15_G_Inst_3__CF_Inst_n6) );
  INV_X1 S_15_G_Inst_3__CF_Inst_U1 ( .A(S_15_Rq1[3]), .ZN(
        S_15_G_Inst_3__CF_Inst_n5) );
  AND2_X1 S_15_G_Inst_4__CF_Inst_U1 ( .A1(S_15_Rq2[1]), .A2(S_15_Rq2[3]), .ZN(
        S_15_G_CF_Out[4]) );
  OR2_X1 S_15_G_Inst_5__CF_Inst_U1 ( .A1(S_15_Rq3[3]), .A2(S_15_Rq2[1]), .ZN(
        S_15_G_CF_Out[5]) );
  AND2_X1 S_15_G_Inst_6__CF_Inst_U1 ( .A1(S_15_Rq3[1]), .A2(S_15_Rq2[3]), .ZN(
        S_15_G_CF_Out[6]) );
  XNOR2_X1 S_15_G_Inst_7__CF_Inst_U2 ( .A(S_15_G_Inst_7__CF_Inst_n3), .B(
        S_15_Rq3[0]), .ZN(S_15_G_CF_Out[7]) );
  NAND2_X1 S_15_G_Inst_7__CF_Inst_U1 ( .A1(S_15_Rq1[1]), .A2(S_15_Rq3[3]), 
        .ZN(S_15_G_Inst_7__CF_Inst_n3) );
  OR2_X1 S_15_G_Inst_8__CF_Inst_U1 ( .A1(S_15_Rq3[3]), .A2(S_15_Rq3[1]), .ZN(
        S_15_G_CF_Out[8]) );
  NOR2_X1 S_15_G_Inst_9__CF_Inst_U2 ( .A1(S_15_Rq1[3]), .A2(
        S_15_G_Inst_9__CF_Inst_n3), .ZN(S_15_G_CF_Out[9]) );
  INV_X1 S_15_G_Inst_9__CF_Inst_U1 ( .A(S_15_Rq1[2]), .ZN(
        S_15_G_Inst_9__CF_Inst_n3) );
  NOR2_X1 S_15_G_Inst_10__CF_Inst_U2 ( .A1(S_15_Rq2[2]), .A2(
        S_15_G_Inst_10__CF_Inst_n3), .ZN(S_15_G_CF_Out[10]) );
  INV_X1 S_15_G_Inst_10__CF_Inst_U1 ( .A(S_15_Rq1[3]), .ZN(
        S_15_G_Inst_10__CF_Inst_n3) );
  XNOR2_X1 S_15_G_Inst_11__CF_Inst_U3 ( .A(S_15_Rq1[1]), .B(
        S_15_G_Inst_11__CF_Inst_n6), .ZN(S_15_G_CF_Out[11]) );
  NAND2_X1 S_15_G_Inst_11__CF_Inst_U2 ( .A1(S_15_Rq1[3]), .A2(
        S_15_G_Inst_11__CF_Inst_n5), .ZN(S_15_G_Inst_11__CF_Inst_n6) );
  INV_X1 S_15_G_Inst_11__CF_Inst_U1 ( .A(S_15_Rq3[2]), .ZN(
        S_15_G_Inst_11__CF_Inst_n5) );
  NOR2_X1 S_15_G_Inst_12__CF_Inst_U2 ( .A1(S_15_Rq2[3]), .A2(
        S_15_G_Inst_12__CF_Inst_n3), .ZN(S_15_G_CF_Out[12]) );
  INV_X1 S_15_G_Inst_12__CF_Inst_U1 ( .A(S_15_Rq1[2]), .ZN(
        S_15_G_Inst_12__CF_Inst_n3) );
  AND2_X1 S_15_G_Inst_13__CF_Inst_U1 ( .A1(S_15_Rq2[2]), .A2(S_15_Rq2[3]), 
        .ZN(S_15_G_CF_Out[13]) );
  XNOR2_X1 S_15_G_Inst_14__CF_Inst_U3 ( .A(S_15_Rq2[1]), .B(
        S_15_G_Inst_14__CF_Inst_n6), .ZN(S_15_G_CF_Out[14]) );
  NAND2_X1 S_15_G_Inst_14__CF_Inst_U2 ( .A1(S_15_Rq3[2]), .A2(
        S_15_G_Inst_14__CF_Inst_n5), .ZN(S_15_G_Inst_14__CF_Inst_n6) );
  INV_X1 S_15_G_Inst_14__CF_Inst_U1 ( .A(S_15_Rq2[3]), .ZN(
        S_15_G_Inst_14__CF_Inst_n5) );
  XNOR2_X1 S_15_G_Inst_15__CF_Inst_U2 ( .A(S_15_G_Inst_15__CF_Inst_n3), .B(
        S_15_Rq3[1]), .ZN(S_15_G_CF_Out[15]) );
  NAND2_X1 S_15_G_Inst_15__CF_Inst_U1 ( .A1(S_15_Rq1[2]), .A2(S_15_Rq3[3]), 
        .ZN(S_15_G_Inst_15__CF_Inst_n3) );
  AND2_X1 S_15_G_Inst_16__CF_Inst_U1 ( .A1(S_15_Rq2[2]), .A2(S_15_Rq3[3]), 
        .ZN(S_15_G_CF_Out[16]) );
  NOR2_X1 S_15_G_Inst_17__CF_Inst_U2 ( .A1(S_15_Rq3[3]), .A2(
        S_15_G_Inst_17__CF_Inst_n3), .ZN(S_15_G_CF_Out[17]) );
  INV_X1 S_15_G_Inst_17__CF_Inst_U1 ( .A(S_15_Rq3[2]), .ZN(
        S_15_G_Inst_17__CF_Inst_n3) );
  XNOR2_X1 S_15_G_InstXOR_0__Compression1_U2 ( .A(
        S_15_G_InstXOR_0__Compression1_n3), .B(S_15_G_CF_Reg[2]), .ZN(
        S_15_G_out1[0]) );
  XNOR2_X1 S_15_G_InstXOR_0__Compression1_U1 ( .A(S_15_G_CF_Reg[0]), .B(
        S_15_G_CF_Reg[1]), .ZN(S_15_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 S_15_G_InstXOR_0__Compression2_U2 ( .A(
        S_15_G_InstXOR_0__Compression2_n3), .B(S_15_G_CF_Reg[5]), .ZN(
        SUB_OUT2[61]) );
  XNOR2_X1 S_15_G_InstXOR_0__Compression2_U1 ( .A(S_15_G_CF_Reg[3]), .B(
        S_15_G_CF_Reg[4]), .ZN(S_15_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 S_15_G_InstXOR_0__Compression3_U2 ( .A(
        S_15_G_InstXOR_0__Compression3_n3), .B(S_15_G_CF_Reg[8]), .ZN(
        SUB_OUT3[61]) );
  XNOR2_X1 S_15_G_InstXOR_0__Compression3_U1 ( .A(S_15_G_CF_Reg[6]), .B(
        S_15_G_CF_Reg[7]), .ZN(S_15_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 S_15_G_InstXOR_1__Compression1_U2 ( .A(
        S_15_G_InstXOR_1__Compression1_n3), .B(S_15_G_CF_Reg[11]), .ZN(
        S_15_G_out1[1]) );
  XNOR2_X1 S_15_G_InstXOR_1__Compression1_U1 ( .A(S_15_G_CF_Reg[9]), .B(
        S_15_G_CF_Reg[10]), .ZN(S_15_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 S_15_G_InstXOR_1__Compression2_U2 ( .A(
        S_15_G_InstXOR_1__Compression2_n3), .B(S_15_G_CF_Reg[14]), .ZN(
        SUB_OUT2[60]) );
  XNOR2_X1 S_15_G_InstXOR_1__Compression2_U1 ( .A(S_15_G_CF_Reg[12]), .B(
        S_15_G_CF_Reg[13]), .ZN(S_15_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 S_15_G_InstXOR_1__Compression3_U2 ( .A(
        S_15_G_InstXOR_1__Compression3_n3), .B(S_15_G_CF_Reg[17]), .ZN(
        SUB_OUT3[60]) );
  XNOR2_X1 S_15_G_InstXOR_1__Compression3_U1 ( .A(S_15_G_CF_Reg[15]), .B(
        S_15_G_CF_Reg[16]), .ZN(S_15_G_InstXOR_1__Compression3_n3) );
  INV_X1 S_15_OutputAffine_U4 ( .A(S_15_G_out1[3]), .ZN(SUB_OUT1[63]) );
  INV_X1 S_15_OutputAffine_U3 ( .A(S_15_G_out1[2]), .ZN(SUB_OUT1[62]) );
  INV_X1 S_15_OutputAffine_U2 ( .A(S_15_G_out1[1]), .ZN(SUB_OUT1[60]) );
  INV_X1 S_15_OutputAffine_U1 ( .A(S_15_G_out1[0]), .ZN(SUB_OUT1[61]) );
  BUF_X1 KE1_RS_U6 ( .A(KEY_EN), .Z(KE1_RS_n7) );
  BUF_X1 KE1_RS_U5 ( .A(KEY_EN), .Z(KE1_RS_n12) );
  BUF_X1 KE1_RS_U4 ( .A(KEY_EN), .Z(KE1_RS_n11) );
  BUF_X1 KE1_RS_U3 ( .A(KEY_EN), .Z(KE1_RS_n10) );
  BUF_X1 KE1_RS_U2 ( .A(KEY_EN), .Z(KE1_RS_n9) );
  BUF_X1 KE1_RS_U1 ( .A(KEY_EN), .Z(KE1_RS_n8) );
  OAI21_X1 KE1_RS_SFF_0_U4 ( .B1(KEY_EN), .B2(KE1_RS_SFF_0_n7), .A(
        KE1_RS_SFF_0_n10), .ZN(KE1_RS_SFF_0_n6) );
  OAI221_X1 KE1_RS_SFF_0_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[0]), .C1(
        KE1_RS_SFF_0_n9), .C2(KEY1[0]), .A(KEY_EN), .ZN(KE1_RS_SFF_0_n10) );
  INV_X1 KE1_RS_SFF_0_U2 ( .A(RESET), .ZN(KE1_RS_SFF_0_n9) );
  DFF_X1 KE1_RS_SFF_0_Q_reg ( .D(KE1_RS_SFF_0_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[56]), .QN(KE1_RS_SFF_0_n7) );
  OAI21_X1 KE1_RS_SFF_1_U4 ( .B1(KEY_EN), .B2(KE1_RS_SFF_1_n8), .A(
        KE1_RS_SFF_1_n11), .ZN(KE1_RS_SFF_1_n7) );
  OAI221_X1 KE1_RS_SFF_1_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[1]), .C1(
        KE1_RS_SFF_1_n10), .C2(KEY1[1]), .A(KEY_EN), .ZN(KE1_RS_SFF_1_n11) );
  INV_X1 KE1_RS_SFF_1_U2 ( .A(RESET), .ZN(KE1_RS_SFF_1_n10) );
  DFF_X1 KE1_RS_SFF_1_Q_reg ( .D(KE1_RS_SFF_1_n7), .CK(CLK), .Q(
        KE1_KEY_PERM[57]), .QN(KE1_RS_SFF_1_n8) );
  OAI21_X1 KE1_RS_SFF_2_U4 ( .B1(KE1_RS_n10), .B2(KE1_RS_SFF_2_n8), .A(
        KE1_RS_SFF_2_n11), .ZN(KE1_RS_SFF_2_n7) );
  OAI221_X1 KE1_RS_SFF_2_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[2]), .C1(
        KE1_RS_SFF_2_n10), .C2(KEY1[2]), .A(KE1_RS_n10), .ZN(KE1_RS_SFF_2_n11)
         );
  INV_X1 KE1_RS_SFF_2_U2 ( .A(RESET), .ZN(KE1_RS_SFF_2_n10) );
  DFF_X1 KE1_RS_SFF_2_Q_reg ( .D(KE1_RS_SFF_2_n7), .CK(CLK), .Q(
        KE1_KEY_PERM[58]), .QN(KE1_RS_SFF_2_n8) );
  OAI21_X1 KE1_RS_SFF_3_U4 ( .B1(KE1_RS_n7), .B2(KE1_RS_SFF_3_n7), .A(
        KE1_RS_SFF_3_n10), .ZN(KE1_RS_SFF_3_n6) );
  OAI221_X1 KE1_RS_SFF_3_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[3]), .C1(
        KE1_RS_SFF_3_n9), .C2(KEY1[3]), .A(KE1_RS_n7), .ZN(KE1_RS_SFF_3_n10)
         );
  INV_X1 KE1_RS_SFF_3_U2 ( .A(RESET), .ZN(KE1_RS_SFF_3_n9) );
  DFF_X1 KE1_RS_SFF_3_Q_reg ( .D(KE1_RS_SFF_3_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[59]), .QN(KE1_RS_SFF_3_n7) );
  OAI21_X1 KE1_RS_SFF_4_U4 ( .B1(KE1_RS_n7), .B2(KE1_RS_SFF_4_n7), .A(
        KE1_RS_SFF_4_n10), .ZN(KE1_RS_SFF_4_n6) );
  OAI221_X1 KE1_RS_SFF_4_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[4]), .C1(
        KE1_RS_SFF_4_n9), .C2(KEY1[4]), .A(KE1_RS_n7), .ZN(KE1_RS_SFF_4_n10)
         );
  INV_X1 KE1_RS_SFF_4_U2 ( .A(RESET), .ZN(KE1_RS_SFF_4_n9) );
  DFF_X1 KE1_RS_SFF_4_Q_reg ( .D(KE1_RS_SFF_4_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[40]), .QN(KE1_RS_SFF_4_n7) );
  OAI21_X1 KE1_RS_SFF_5_U4 ( .B1(KE1_RS_n7), .B2(KE1_RS_SFF_5_n7), .A(
        KE1_RS_SFF_5_n10), .ZN(KE1_RS_SFF_5_n6) );
  OAI221_X1 KE1_RS_SFF_5_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[5]), .C1(
        KE1_RS_SFF_5_n9), .C2(KEY1[5]), .A(KE1_RS_n7), .ZN(KE1_RS_SFF_5_n10)
         );
  INV_X1 KE1_RS_SFF_5_U2 ( .A(RESET), .ZN(KE1_RS_SFF_5_n9) );
  DFF_X1 KE1_RS_SFF_5_Q_reg ( .D(KE1_RS_SFF_5_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[41]), .QN(KE1_RS_SFF_5_n7) );
  OAI21_X1 KE1_RS_SFF_6_U4 ( .B1(KE1_RS_n7), .B2(KE1_RS_SFF_6_n7), .A(
        KE1_RS_SFF_6_n10), .ZN(KE1_RS_SFF_6_n6) );
  OAI221_X1 KE1_RS_SFF_6_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[6]), .C1(
        KE1_RS_SFF_6_n9), .C2(KEY1[6]), .A(KE1_RS_n7), .ZN(KE1_RS_SFF_6_n10)
         );
  INV_X1 KE1_RS_SFF_6_U2 ( .A(RESET), .ZN(KE1_RS_SFF_6_n9) );
  DFF_X1 KE1_RS_SFF_6_Q_reg ( .D(KE1_RS_SFF_6_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[42]), .QN(KE1_RS_SFF_6_n7) );
  OAI21_X1 KE1_RS_SFF_7_U4 ( .B1(KE1_RS_n7), .B2(KE1_RS_SFF_7_n7), .A(
        KE1_RS_SFF_7_n10), .ZN(KE1_RS_SFF_7_n6) );
  OAI221_X1 KE1_RS_SFF_7_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[7]), .C1(
        KE1_RS_SFF_7_n9), .C2(KEY1[7]), .A(KE1_RS_n7), .ZN(KE1_RS_SFF_7_n10)
         );
  INV_X1 KE1_RS_SFF_7_U2 ( .A(RESET), .ZN(KE1_RS_SFF_7_n9) );
  DFF_X1 KE1_RS_SFF_7_Q_reg ( .D(KE1_RS_SFF_7_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[43]), .QN(KE1_RS_SFF_7_n7) );
  OAI21_X1 KE1_RS_SFF_8_U4 ( .B1(KE1_RS_n7), .B2(KE1_RS_SFF_8_n7), .A(
        KE1_RS_SFF_8_n10), .ZN(KE1_RS_SFF_8_n6) );
  OAI221_X1 KE1_RS_SFF_8_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[8]), .C1(
        KE1_RS_SFF_8_n9), .C2(KEY1[8]), .A(KE1_RS_n7), .ZN(KE1_RS_SFF_8_n10)
         );
  INV_X1 KE1_RS_SFF_8_U2 ( .A(RESET), .ZN(KE1_RS_SFF_8_n9) );
  DFF_X1 KE1_RS_SFF_8_Q_reg ( .D(KE1_RS_SFF_8_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[48]), .QN(KE1_RS_SFF_8_n7) );
  OAI21_X1 KE1_RS_SFF_9_U4 ( .B1(KE1_RS_n7), .B2(KE1_RS_SFF_9_n7), .A(
        KE1_RS_SFF_9_n10), .ZN(KE1_RS_SFF_9_n6) );
  OAI221_X1 KE1_RS_SFF_9_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[9]), .C1(
        KE1_RS_SFF_9_n9), .C2(KEY1[9]), .A(KE1_RS_n7), .ZN(KE1_RS_SFF_9_n10)
         );
  INV_X1 KE1_RS_SFF_9_U2 ( .A(RESET), .ZN(KE1_RS_SFF_9_n9) );
  DFF_X1 KE1_RS_SFF_9_Q_reg ( .D(KE1_RS_SFF_9_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[49]), .QN(KE1_RS_SFF_9_n7) );
  OAI21_X1 KE1_RS_SFF_10_U4 ( .B1(KE1_RS_n7), .B2(KE1_RS_SFF_10_n7), .A(
        KE1_RS_SFF_10_n10), .ZN(KE1_RS_SFF_10_n6) );
  OAI221_X1 KE1_RS_SFF_10_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[10]), .C1(
        KE1_RS_SFF_10_n9), .C2(KEY1[10]), .A(KE1_RS_n7), .ZN(KE1_RS_SFF_10_n10) );
  INV_X1 KE1_RS_SFF_10_U2 ( .A(RESET), .ZN(KE1_RS_SFF_10_n9) );
  DFF_X1 KE1_RS_SFF_10_Q_reg ( .D(KE1_RS_SFF_10_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[50]), .QN(KE1_RS_SFF_10_n7) );
  OAI21_X1 KE1_RS_SFF_11_U4 ( .B1(KE1_RS_n8), .B2(KE1_RS_SFF_11_n7), .A(
        KE1_RS_SFF_11_n10), .ZN(KE1_RS_SFF_11_n6) );
  OAI221_X1 KE1_RS_SFF_11_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[11]), .C1(
        KE1_RS_SFF_11_n9), .C2(KEY1[11]), .A(KE1_RS_n8), .ZN(KE1_RS_SFF_11_n10) );
  INV_X1 KE1_RS_SFF_11_U2 ( .A(RESET), .ZN(KE1_RS_SFF_11_n9) );
  DFF_X1 KE1_RS_SFF_11_Q_reg ( .D(KE1_RS_SFF_11_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[51]), .QN(KE1_RS_SFF_11_n7) );
  OAI21_X1 KE1_RS_SFF_12_U4 ( .B1(KE1_RS_n8), .B2(KE1_RS_SFF_12_n7), .A(
        KE1_RS_SFF_12_n10), .ZN(KE1_RS_SFF_12_n6) );
  OAI221_X1 KE1_RS_SFF_12_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[12]), .C1(
        KE1_RS_SFF_12_n9), .C2(KEY1[12]), .A(KE1_RS_n8), .ZN(KE1_RS_SFF_12_n10) );
  INV_X1 KE1_RS_SFF_12_U2 ( .A(RESET), .ZN(KE1_RS_SFF_12_n9) );
  DFF_X1 KE1_RS_SFF_12_Q_reg ( .D(KE1_RS_SFF_12_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[36]), .QN(KE1_RS_SFF_12_n7) );
  OAI21_X1 KE1_RS_SFF_13_U4 ( .B1(KE1_RS_n9), .B2(KE1_RS_SFF_13_n8), .A(
        KE1_RS_SFF_13_n11), .ZN(KE1_RS_SFF_13_n7) );
  OAI221_X1 KE1_RS_SFF_13_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[13]), .C1(
        KE1_RS_SFF_13_n10), .C2(KEY1[13]), .A(KE1_RS_n9), .ZN(
        KE1_RS_SFF_13_n11) );
  INV_X1 KE1_RS_SFF_13_U2 ( .A(RESET), .ZN(KE1_RS_SFF_13_n10) );
  DFF_X1 KE1_RS_SFF_13_Q_reg ( .D(KE1_RS_SFF_13_n7), .CK(CLK), .Q(
        KE1_KEY_PERM[37]), .QN(KE1_RS_SFF_13_n8) );
  OAI21_X1 KE1_RS_SFF_14_U4 ( .B1(KE1_RS_n8), .B2(KE1_RS_SFF_14_n8), .A(
        KE1_RS_SFF_14_n11), .ZN(KE1_RS_SFF_14_n7) );
  OAI221_X1 KE1_RS_SFF_14_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[14]), .C1(
        KE1_RS_SFF_14_n10), .C2(KEY1[14]), .A(KE1_RS_n8), .ZN(
        KE1_RS_SFF_14_n11) );
  INV_X1 KE1_RS_SFF_14_U2 ( .A(RESET), .ZN(KE1_RS_SFF_14_n10) );
  DFF_X1 KE1_RS_SFF_14_Q_reg ( .D(KE1_RS_SFF_14_n7), .CK(CLK), .Q(
        KE1_KEY_PERM[38]), .QN(KE1_RS_SFF_14_n8) );
  OAI21_X1 KE1_RS_SFF_15_U4 ( .B1(KE1_RS_n8), .B2(KE1_RS_SFF_15_n7), .A(
        KE1_RS_SFF_15_n10), .ZN(KE1_RS_SFF_15_n6) );
  OAI221_X1 KE1_RS_SFF_15_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[15]), .C1(
        KE1_RS_SFF_15_n9), .C2(KEY1[15]), .A(KE1_RS_n8), .ZN(KE1_RS_SFF_15_n10) );
  INV_X1 KE1_RS_SFF_15_U2 ( .A(RESET), .ZN(KE1_RS_SFF_15_n9) );
  DFF_X1 KE1_RS_SFF_15_Q_reg ( .D(KE1_RS_SFF_15_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[39]), .QN(KE1_RS_SFF_15_n7) );
  OAI21_X1 KE1_RS_SFF_16_U4 ( .B1(KE1_RS_n8), .B2(KE1_RS_SFF_16_n7), .A(
        KE1_RS_SFF_16_n10), .ZN(KE1_RS_SFF_16_n6) );
  OAI221_X1 KE1_RS_SFF_16_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[16]), .C1(
        KE1_RS_SFF_16_n9), .C2(KEY1[16]), .A(KE1_RS_n8), .ZN(KE1_RS_SFF_16_n10) );
  INV_X1 KE1_RS_SFF_16_U2 ( .A(RESET), .ZN(KE1_RS_SFF_16_n9) );
  DFF_X1 KE1_RS_SFF_16_Q_reg ( .D(KE1_RS_SFF_16_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[32]), .QN(KE1_RS_SFF_16_n7) );
  OAI21_X1 KE1_RS_SFF_17_U4 ( .B1(KE1_RS_n8), .B2(KE1_RS_SFF_17_n7), .A(
        KE1_RS_SFF_17_n10), .ZN(KE1_RS_SFF_17_n6) );
  OAI221_X1 KE1_RS_SFF_17_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[17]), .C1(
        KE1_RS_SFF_17_n9), .C2(KEY1[17]), .A(KE1_RS_n8), .ZN(KE1_RS_SFF_17_n10) );
  INV_X1 KE1_RS_SFF_17_U2 ( .A(RESET), .ZN(KE1_RS_SFF_17_n9) );
  DFF_X1 KE1_RS_SFF_17_Q_reg ( .D(KE1_RS_SFF_17_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[33]), .QN(KE1_RS_SFF_17_n7) );
  OAI21_X1 KE1_RS_SFF_18_U4 ( .B1(KE1_RS_n8), .B2(KE1_RS_SFF_18_n7), .A(
        KE1_RS_SFF_18_n10), .ZN(KE1_RS_SFF_18_n6) );
  OAI221_X1 KE1_RS_SFF_18_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[18]), .C1(
        KE1_RS_SFF_18_n9), .C2(KEY1[18]), .A(KE1_RS_n8), .ZN(KE1_RS_SFF_18_n10) );
  INV_X1 KE1_RS_SFF_18_U2 ( .A(RESET), .ZN(KE1_RS_SFF_18_n9) );
  DFF_X1 KE1_RS_SFF_18_Q_reg ( .D(KE1_RS_SFF_18_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[34]), .QN(KE1_RS_SFF_18_n7) );
  OAI21_X1 KE1_RS_SFF_19_U4 ( .B1(KE1_RS_n8), .B2(KE1_RS_SFF_19_n7), .A(
        KE1_RS_SFF_19_n10), .ZN(KE1_RS_SFF_19_n6) );
  OAI221_X1 KE1_RS_SFF_19_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[19]), .C1(
        KE1_RS_SFF_19_n9), .C2(KEY1[19]), .A(KE1_RS_n8), .ZN(KE1_RS_SFF_19_n10) );
  INV_X1 KE1_RS_SFF_19_U2 ( .A(RESET), .ZN(KE1_RS_SFF_19_n9) );
  DFF_X1 KE1_RS_SFF_19_Q_reg ( .D(KE1_RS_SFF_19_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[35]), .QN(KE1_RS_SFF_19_n7) );
  OAI21_X1 KE1_RS_SFF_20_U4 ( .B1(KE1_RS_n8), .B2(KE1_RS_SFF_20_n7), .A(
        KE1_RS_SFF_20_n10), .ZN(KE1_RS_SFF_20_n6) );
  OAI221_X1 KE1_RS_SFF_20_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[20]), .C1(
        KE1_RS_SFF_20_n9), .C2(KEY1[20]), .A(KE1_RS_n8), .ZN(KE1_RS_SFF_20_n10) );
  INV_X1 KE1_RS_SFF_20_U2 ( .A(RESET), .ZN(KE1_RS_SFF_20_n9) );
  DFF_X1 KE1_RS_SFF_20_Q_reg ( .D(KE1_RS_SFF_20_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[44]), .QN(KE1_RS_SFF_20_n7) );
  OAI21_X1 KE1_RS_SFF_21_U4 ( .B1(KE1_RS_n9), .B2(KE1_RS_SFF_21_n7), .A(
        KE1_RS_SFF_21_n10), .ZN(KE1_RS_SFF_21_n6) );
  OAI221_X1 KE1_RS_SFF_21_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[21]), .C1(
        KE1_RS_SFF_21_n9), .C2(KEY1[21]), .A(KE1_RS_n9), .ZN(KE1_RS_SFF_21_n10) );
  INV_X1 KE1_RS_SFF_21_U2 ( .A(RESET), .ZN(KE1_RS_SFF_21_n9) );
  DFF_X1 KE1_RS_SFF_21_Q_reg ( .D(KE1_RS_SFF_21_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[45]), .QN(KE1_RS_SFF_21_n7) );
  OAI21_X1 KE1_RS_SFF_22_U4 ( .B1(KE1_RS_n9), .B2(KE1_RS_SFF_22_n7), .A(
        KE1_RS_SFF_22_n10), .ZN(KE1_RS_SFF_22_n6) );
  OAI221_X1 KE1_RS_SFF_22_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[22]), .C1(
        KE1_RS_SFF_22_n9), .C2(KEY1[22]), .A(KE1_RS_n9), .ZN(KE1_RS_SFF_22_n10) );
  INV_X1 KE1_RS_SFF_22_U2 ( .A(RESET), .ZN(KE1_RS_SFF_22_n9) );
  DFF_X1 KE1_RS_SFF_22_Q_reg ( .D(KE1_RS_SFF_22_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[46]), .QN(KE1_RS_SFF_22_n7) );
  OAI21_X1 KE1_RS_SFF_23_U4 ( .B1(KE1_RS_n9), .B2(KE1_RS_SFF_23_n7), .A(
        KE1_RS_SFF_23_n10), .ZN(KE1_RS_SFF_23_n6) );
  OAI221_X1 KE1_RS_SFF_23_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[23]), .C1(
        KE1_RS_SFF_23_n9), .C2(KEY1[23]), .A(KE1_RS_n9), .ZN(KE1_RS_SFF_23_n10) );
  INV_X1 KE1_RS_SFF_23_U2 ( .A(RESET), .ZN(KE1_RS_SFF_23_n9) );
  DFF_X1 KE1_RS_SFF_23_Q_reg ( .D(KE1_RS_SFF_23_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[47]), .QN(KE1_RS_SFF_23_n7) );
  OAI21_X1 KE1_RS_SFF_24_U4 ( .B1(KE1_RS_n9), .B2(KE1_RS_SFF_24_n7), .A(
        KE1_RS_SFF_24_n10), .ZN(KE1_RS_SFF_24_n6) );
  OAI221_X1 KE1_RS_SFF_24_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[24]), .C1(
        KE1_RS_SFF_24_n9), .C2(KEY1[24]), .A(KE1_RS_n9), .ZN(KE1_RS_SFF_24_n10) );
  INV_X1 KE1_RS_SFF_24_U2 ( .A(RESET), .ZN(KE1_RS_SFF_24_n9) );
  DFF_X1 KE1_RS_SFF_24_Q_reg ( .D(KE1_RS_SFF_24_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[60]), .QN(KE1_RS_SFF_24_n7) );
  OAI21_X1 KE1_RS_SFF_25_U4 ( .B1(KEY_EN), .B2(KE1_RS_SFF_25_n8), .A(
        KE1_RS_SFF_25_n11), .ZN(KE1_RS_SFF_25_n7) );
  OAI221_X1 KE1_RS_SFF_25_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[25]), .C1(
        KE1_RS_SFF_25_n10), .C2(KEY1[25]), .A(KEY_EN), .ZN(KE1_RS_SFF_25_n11)
         );
  INV_X1 KE1_RS_SFF_25_U2 ( .A(RESET), .ZN(KE1_RS_SFF_25_n10) );
  DFF_X1 KE1_RS_SFF_25_Q_reg ( .D(KE1_RS_SFF_25_n7), .CK(CLK), .Q(
        KE1_KEY_PERM[61]), .QN(KE1_RS_SFF_25_n8) );
  OAI21_X1 KE1_RS_SFF_26_U4 ( .B1(KEY_EN), .B2(KE1_RS_SFF_26_n8), .A(
        KE1_RS_SFF_26_n11), .ZN(KE1_RS_SFF_26_n7) );
  OAI221_X1 KE1_RS_SFF_26_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[26]), .C1(
        KE1_RS_SFF_26_n10), .C2(KEY1[26]), .A(KEY_EN), .ZN(KE1_RS_SFF_26_n11)
         );
  INV_X1 KE1_RS_SFF_26_U2 ( .A(RESET), .ZN(KE1_RS_SFF_26_n10) );
  DFF_X1 KE1_RS_SFF_26_Q_reg ( .D(KE1_RS_SFF_26_n7), .CK(CLK), .Q(
        KE1_KEY_PERM[62]), .QN(KE1_RS_SFF_26_n8) );
  OAI21_X1 KE1_RS_SFF_27_U4 ( .B1(KE1_RS_n9), .B2(KE1_RS_SFF_27_n7), .A(
        KE1_RS_SFF_27_n10), .ZN(KE1_RS_SFF_27_n6) );
  OAI221_X1 KE1_RS_SFF_27_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[27]), .C1(
        KE1_RS_SFF_27_n9), .C2(KEY1[27]), .A(KE1_RS_n9), .ZN(KE1_RS_SFF_27_n10) );
  INV_X1 KE1_RS_SFF_27_U2 ( .A(RESET), .ZN(KE1_RS_SFF_27_n9) );
  DFF_X1 KE1_RS_SFF_27_Q_reg ( .D(KE1_RS_SFF_27_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[63]), .QN(KE1_RS_SFF_27_n7) );
  OAI21_X1 KE1_RS_SFF_28_U4 ( .B1(KE1_RS_n9), .B2(KE1_RS_SFF_28_n7), .A(
        KE1_RS_SFF_28_n10), .ZN(KE1_RS_SFF_28_n6) );
  OAI221_X1 KE1_RS_SFF_28_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[28]), .C1(
        KE1_RS_SFF_28_n9), .C2(KEY1[28]), .A(KE1_RS_n9), .ZN(KE1_RS_SFF_28_n10) );
  INV_X1 KE1_RS_SFF_28_U2 ( .A(RESET), .ZN(KE1_RS_SFF_28_n9) );
  DFF_X1 KE1_RS_SFF_28_Q_reg ( .D(KE1_RS_SFF_28_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[52]), .QN(KE1_RS_SFF_28_n7) );
  OAI21_X1 KE1_RS_SFF_29_U4 ( .B1(KE1_RS_n9), .B2(KE1_RS_SFF_29_n7), .A(
        KE1_RS_SFF_29_n10), .ZN(KE1_RS_SFF_29_n6) );
  OAI221_X1 KE1_RS_SFF_29_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[29]), .C1(
        KE1_RS_SFF_29_n9), .C2(KEY1[29]), .A(KE1_RS_n9), .ZN(KE1_RS_SFF_29_n10) );
  INV_X1 KE1_RS_SFF_29_U2 ( .A(RESET), .ZN(KE1_RS_SFF_29_n9) );
  DFF_X1 KE1_RS_SFF_29_Q_reg ( .D(KE1_RS_SFF_29_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[53]), .QN(KE1_RS_SFF_29_n7) );
  OAI21_X1 KE1_RS_SFF_30_U4 ( .B1(KE1_RS_n9), .B2(KE1_RS_SFF_30_n7), .A(
        KE1_RS_SFF_30_n10), .ZN(KE1_RS_SFF_30_n6) );
  OAI221_X1 KE1_RS_SFF_30_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[30]), .C1(
        KE1_RS_SFF_30_n9), .C2(KEY1[30]), .A(KE1_RS_n9), .ZN(KE1_RS_SFF_30_n10) );
  INV_X1 KE1_RS_SFF_30_U2 ( .A(RESET), .ZN(KE1_RS_SFF_30_n9) );
  DFF_X1 KE1_RS_SFF_30_Q_reg ( .D(KE1_RS_SFF_30_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[54]), .QN(KE1_RS_SFF_30_n7) );
  OAI21_X1 KE1_RS_SFF_31_U4 ( .B1(KE1_RS_n10), .B2(KE1_RS_SFF_31_n7), .A(
        KE1_RS_SFF_31_n10), .ZN(KE1_RS_SFF_31_n6) );
  OAI221_X1 KE1_RS_SFF_31_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[31]), .C1(
        KE1_RS_SFF_31_n9), .C2(KEY1[31]), .A(KE1_RS_n10), .ZN(
        KE1_RS_SFF_31_n10) );
  INV_X1 KE1_RS_SFF_31_U2 ( .A(RESET), .ZN(KE1_RS_SFF_31_n9) );
  DFF_X1 KE1_RS_SFF_31_Q_reg ( .D(KE1_RS_SFF_31_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[55]), .QN(KE1_RS_SFF_31_n7) );
  OAI21_X1 KE1_RS_SFF_32_U4 ( .B1(KE1_RS_n10), .B2(KE1_RS_SFF_32_n7), .A(
        KE1_RS_SFF_32_n10), .ZN(KE1_RS_SFF_32_n6) );
  OAI221_X1 KE1_RS_SFF_32_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[32]), .C1(
        KE1_RS_SFF_32_n9), .C2(KEY1[32]), .A(KE1_RS_n10), .ZN(
        KE1_RS_SFF_32_n10) );
  INV_X1 KE1_RS_SFF_32_U2 ( .A(RESET), .ZN(KE1_RS_SFF_32_n9) );
  DFF_X1 KE1_RS_SFF_32_Q_reg ( .D(KE1_RS_SFF_32_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[0]), .QN(KE1_RS_SFF_32_n7) );
  OAI21_X1 KE1_RS_SFF_33_U4 ( .B1(KE1_RS_n10), .B2(KE1_RS_SFF_33_n7), .A(
        KE1_RS_SFF_33_n10), .ZN(KE1_RS_SFF_33_n6) );
  OAI221_X1 KE1_RS_SFF_33_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[33]), .C1(
        KE1_RS_SFF_33_n9), .C2(KEY1[33]), .A(KE1_RS_n10), .ZN(
        KE1_RS_SFF_33_n10) );
  INV_X1 KE1_RS_SFF_33_U2 ( .A(RESET), .ZN(KE1_RS_SFF_33_n9) );
  DFF_X1 KE1_RS_SFF_33_Q_reg ( .D(KE1_RS_SFF_33_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[1]), .QN(KE1_RS_SFF_33_n7) );
  OAI21_X1 KE1_RS_SFF_34_U4 ( .B1(KE1_RS_n10), .B2(KE1_RS_SFF_34_n7), .A(
        KE1_RS_SFF_34_n10), .ZN(KE1_RS_SFF_34_n6) );
  OAI221_X1 KE1_RS_SFF_34_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[34]), .C1(
        KE1_RS_SFF_34_n9), .C2(KEY1[34]), .A(KE1_RS_n10), .ZN(
        KE1_RS_SFF_34_n10) );
  INV_X1 KE1_RS_SFF_34_U2 ( .A(RESET), .ZN(KE1_RS_SFF_34_n9) );
  DFF_X1 KE1_RS_SFF_34_Q_reg ( .D(KE1_RS_SFF_34_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[2]), .QN(KE1_RS_SFF_34_n7) );
  OAI21_X1 KE1_RS_SFF_35_U4 ( .B1(KE1_RS_n10), .B2(KE1_RS_SFF_35_n7), .A(
        KE1_RS_SFF_35_n10), .ZN(KE1_RS_SFF_35_n6) );
  OAI221_X1 KE1_RS_SFF_35_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[35]), .C1(
        KE1_RS_SFF_35_n9), .C2(KEY1[35]), .A(KE1_RS_n10), .ZN(
        KE1_RS_SFF_35_n10) );
  INV_X1 KE1_RS_SFF_35_U2 ( .A(RESET), .ZN(KE1_RS_SFF_35_n9) );
  DFF_X1 KE1_RS_SFF_35_Q_reg ( .D(KE1_RS_SFF_35_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[3]), .QN(KE1_RS_SFF_35_n7) );
  OAI21_X1 KE1_RS_SFF_36_U4 ( .B1(KE1_RS_n10), .B2(KE1_RS_SFF_36_n7), .A(
        KE1_RS_SFF_36_n10), .ZN(KE1_RS_SFF_36_n6) );
  OAI221_X1 KE1_RS_SFF_36_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[36]), .C1(
        KE1_RS_SFF_36_n9), .C2(KEY1[36]), .A(KE1_RS_n10), .ZN(
        KE1_RS_SFF_36_n10) );
  INV_X1 KE1_RS_SFF_36_U2 ( .A(RESET), .ZN(KE1_RS_SFF_36_n9) );
  DFF_X1 KE1_RS_SFF_36_Q_reg ( .D(KE1_RS_SFF_36_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[4]), .QN(KE1_RS_SFF_36_n7) );
  OAI21_X1 KE1_RS_SFF_37_U4 ( .B1(KEY_EN), .B2(KE1_RS_SFF_37_n8), .A(
        KE1_RS_SFF_37_n11), .ZN(KE1_RS_SFF_37_n7) );
  OAI221_X1 KE1_RS_SFF_37_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[37]), .C1(
        KE1_RS_SFF_37_n10), .C2(KEY1[37]), .A(KEY_EN), .ZN(KE1_RS_SFF_37_n11)
         );
  INV_X1 KE1_RS_SFF_37_U2 ( .A(RESET), .ZN(KE1_RS_SFF_37_n10) );
  DFF_X1 KE1_RS_SFF_37_Q_reg ( .D(KE1_RS_SFF_37_n7), .CK(CLK), .Q(
        KE1_KEY_PERM[5]), .QN(KE1_RS_SFF_37_n8) );
  OAI21_X1 KE1_RS_SFF_38_U4 ( .B1(KEY_EN), .B2(KE1_RS_SFF_38_n8), .A(
        KE1_RS_SFF_38_n11), .ZN(KE1_RS_SFF_38_n7) );
  OAI221_X1 KE1_RS_SFF_38_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[38]), .C1(
        KE1_RS_SFF_38_n10), .C2(KEY1[38]), .A(KEY_EN), .ZN(KE1_RS_SFF_38_n11)
         );
  INV_X1 KE1_RS_SFF_38_U2 ( .A(RESET), .ZN(KE1_RS_SFF_38_n10) );
  DFF_X1 KE1_RS_SFF_38_Q_reg ( .D(KE1_RS_SFF_38_n7), .CK(CLK), .Q(
        KE1_KEY_PERM[6]), .QN(KE1_RS_SFF_38_n8) );
  OAI21_X1 KE1_RS_SFF_39_U4 ( .B1(KE1_RS_n10), .B2(KE1_RS_SFF_39_n7), .A(
        KE1_RS_SFF_39_n10), .ZN(KE1_RS_SFF_39_n6) );
  OAI221_X1 KE1_RS_SFF_39_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[39]), .C1(
        KE1_RS_SFF_39_n9), .C2(KEY1[39]), .A(KE1_RS_n10), .ZN(
        KE1_RS_SFF_39_n10) );
  INV_X1 KE1_RS_SFF_39_U2 ( .A(RESET), .ZN(KE1_RS_SFF_39_n9) );
  DFF_X1 KE1_RS_SFF_39_Q_reg ( .D(KE1_RS_SFF_39_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[7]), .QN(KE1_RS_SFF_39_n7) );
  OAI21_X1 KE1_RS_SFF_40_U4 ( .B1(KE1_RS_n10), .B2(KE1_RS_SFF_40_n7), .A(
        KE1_RS_SFF_40_n10), .ZN(KE1_RS_SFF_40_n6) );
  OAI221_X1 KE1_RS_SFF_40_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[40]), .C1(
        KE1_RS_SFF_40_n9), .C2(KEY1[40]), .A(KE1_RS_n10), .ZN(
        KE1_RS_SFF_40_n10) );
  INV_X1 KE1_RS_SFF_40_U2 ( .A(RESET), .ZN(KE1_RS_SFF_40_n9) );
  DFF_X1 KE1_RS_SFF_40_Q_reg ( .D(KE1_RS_SFF_40_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[8]), .QN(KE1_RS_SFF_40_n7) );
  OAI21_X1 KE1_RS_SFF_41_U4 ( .B1(KE1_RS_n11), .B2(KE1_RS_SFF_41_n7), .A(
        KE1_RS_SFF_41_n10), .ZN(KE1_RS_SFF_41_n6) );
  OAI221_X1 KE1_RS_SFF_41_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[41]), .C1(
        KE1_RS_SFF_41_n9), .C2(KEY1[41]), .A(KE1_RS_n11), .ZN(
        KE1_RS_SFF_41_n10) );
  INV_X1 KE1_RS_SFF_41_U2 ( .A(RESET), .ZN(KE1_RS_SFF_41_n9) );
  DFF_X1 KE1_RS_SFF_41_Q_reg ( .D(KE1_RS_SFF_41_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[9]), .QN(KE1_RS_SFF_41_n7) );
  OAI21_X1 KE1_RS_SFF_42_U4 ( .B1(KE1_RS_n11), .B2(KE1_RS_SFF_42_n7), .A(
        KE1_RS_SFF_42_n10), .ZN(KE1_RS_SFF_42_n6) );
  OAI221_X1 KE1_RS_SFF_42_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[42]), .C1(
        KE1_RS_SFF_42_n9), .C2(KEY1[42]), .A(KE1_RS_n11), .ZN(
        KE1_RS_SFF_42_n10) );
  INV_X1 KE1_RS_SFF_42_U2 ( .A(RESET), .ZN(KE1_RS_SFF_42_n9) );
  DFF_X1 KE1_RS_SFF_42_Q_reg ( .D(KE1_RS_SFF_42_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[10]), .QN(KE1_RS_SFF_42_n7) );
  OAI21_X1 KE1_RS_SFF_43_U4 ( .B1(KE1_RS_n11), .B2(KE1_RS_SFF_43_n7), .A(
        KE1_RS_SFF_43_n10), .ZN(KE1_RS_SFF_43_n6) );
  OAI221_X1 KE1_RS_SFF_43_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[43]), .C1(
        KE1_RS_SFF_43_n9), .C2(KEY1[43]), .A(KE1_RS_n11), .ZN(
        KE1_RS_SFF_43_n10) );
  INV_X1 KE1_RS_SFF_43_U2 ( .A(RESET), .ZN(KE1_RS_SFF_43_n9) );
  DFF_X1 KE1_RS_SFF_43_Q_reg ( .D(KE1_RS_SFF_43_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[11]), .QN(KE1_RS_SFF_43_n7) );
  OAI21_X1 KE1_RS_SFF_44_U4 ( .B1(KE1_RS_n11), .B2(KE1_RS_SFF_44_n7), .A(
        KE1_RS_SFF_44_n10), .ZN(KE1_RS_SFF_44_n6) );
  OAI221_X1 KE1_RS_SFF_44_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[44]), .C1(
        KE1_RS_SFF_44_n9), .C2(KEY1[44]), .A(KE1_RS_n11), .ZN(
        KE1_RS_SFF_44_n10) );
  INV_X1 KE1_RS_SFF_44_U2 ( .A(RESET), .ZN(KE1_RS_SFF_44_n9) );
  DFF_X1 KE1_RS_SFF_44_Q_reg ( .D(KE1_RS_SFF_44_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[12]), .QN(KE1_RS_SFF_44_n7) );
  OAI21_X1 KE1_RS_SFF_45_U4 ( .B1(KE1_RS_n11), .B2(KE1_RS_SFF_45_n7), .A(
        KE1_RS_SFF_45_n10), .ZN(KE1_RS_SFF_45_n6) );
  OAI221_X1 KE1_RS_SFF_45_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[45]), .C1(
        KE1_RS_SFF_45_n9), .C2(KEY1[45]), .A(KE1_RS_n11), .ZN(
        KE1_RS_SFF_45_n10) );
  INV_X1 KE1_RS_SFF_45_U2 ( .A(RESET), .ZN(KE1_RS_SFF_45_n9) );
  DFF_X1 KE1_RS_SFF_45_Q_reg ( .D(KE1_RS_SFF_45_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[13]), .QN(KE1_RS_SFF_45_n7) );
  OAI21_X1 KE1_RS_SFF_46_U4 ( .B1(KE1_RS_n11), .B2(KE1_RS_SFF_46_n7), .A(
        KE1_RS_SFF_46_n10), .ZN(KE1_RS_SFF_46_n6) );
  OAI221_X1 KE1_RS_SFF_46_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[46]), .C1(
        KE1_RS_SFF_46_n9), .C2(KEY1[46]), .A(KE1_RS_n11), .ZN(
        KE1_RS_SFF_46_n10) );
  INV_X1 KE1_RS_SFF_46_U2 ( .A(RESET), .ZN(KE1_RS_SFF_46_n9) );
  DFF_X1 KE1_RS_SFF_46_Q_reg ( .D(KE1_RS_SFF_46_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[14]), .QN(KE1_RS_SFF_46_n7) );
  OAI21_X1 KE1_RS_SFF_47_U4 ( .B1(KE1_RS_n11), .B2(KE1_RS_SFF_47_n7), .A(
        KE1_RS_SFF_47_n10), .ZN(KE1_RS_SFF_47_n6) );
  OAI221_X1 KE1_RS_SFF_47_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[47]), .C1(
        KE1_RS_SFF_47_n9), .C2(KEY1[47]), .A(KE1_RS_n11), .ZN(
        KE1_RS_SFF_47_n10) );
  INV_X1 KE1_RS_SFF_47_U2 ( .A(RESET), .ZN(KE1_RS_SFF_47_n9) );
  DFF_X1 KE1_RS_SFF_47_Q_reg ( .D(KE1_RS_SFF_47_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[15]), .QN(KE1_RS_SFF_47_n7) );
  OAI21_X1 KE1_RS_SFF_48_U4 ( .B1(KE1_RS_n11), .B2(KE1_RS_SFF_48_n7), .A(
        KE1_RS_SFF_48_n10), .ZN(KE1_RS_SFF_48_n6) );
  OAI221_X1 KE1_RS_SFF_48_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[48]), .C1(
        KE1_RS_SFF_48_n9), .C2(KEY1[48]), .A(KE1_RS_n11), .ZN(
        KE1_RS_SFF_48_n10) );
  INV_X1 KE1_RS_SFF_48_U2 ( .A(RESET), .ZN(KE1_RS_SFF_48_n9) );
  DFF_X1 KE1_RS_SFF_48_Q_reg ( .D(KE1_RS_SFF_48_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[16]), .QN(KE1_RS_SFF_48_n7) );
  OAI21_X1 KE1_RS_SFF_49_U4 ( .B1(KEY_EN), .B2(KE1_RS_SFF_49_n8), .A(
        KE1_RS_SFF_49_n11), .ZN(KE1_RS_SFF_49_n7) );
  OAI221_X1 KE1_RS_SFF_49_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[49]), .C1(
        KE1_RS_SFF_49_n10), .C2(KEY1[49]), .A(KEY_EN), .ZN(KE1_RS_SFF_49_n11)
         );
  INV_X1 KE1_RS_SFF_49_U2 ( .A(RESET), .ZN(KE1_RS_SFF_49_n10) );
  DFF_X1 KE1_RS_SFF_49_Q_reg ( .D(KE1_RS_SFF_49_n7), .CK(CLK), .Q(
        KE1_KEY_PERM[17]), .QN(KE1_RS_SFF_49_n8) );
  OAI21_X1 KE1_RS_SFF_50_U4 ( .B1(KEY_EN), .B2(KE1_RS_SFF_50_n8), .A(
        KE1_RS_SFF_50_n11), .ZN(KE1_RS_SFF_50_n7) );
  OAI221_X1 KE1_RS_SFF_50_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[50]), .C1(
        KE1_RS_SFF_50_n10), .C2(KEY1[50]), .A(KEY_EN), .ZN(KE1_RS_SFF_50_n11)
         );
  INV_X1 KE1_RS_SFF_50_U2 ( .A(RESET), .ZN(KE1_RS_SFF_50_n10) );
  DFF_X1 KE1_RS_SFF_50_Q_reg ( .D(KE1_RS_SFF_50_n7), .CK(CLK), .Q(
        KE1_KEY_PERM[18]), .QN(KE1_RS_SFF_50_n8) );
  OAI21_X1 KE1_RS_SFF_51_U4 ( .B1(KE1_RS_n12), .B2(KE1_RS_SFF_51_n7), .A(
        KE1_RS_SFF_51_n10), .ZN(KE1_RS_SFF_51_n6) );
  OAI221_X1 KE1_RS_SFF_51_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[51]), .C1(
        KE1_RS_SFF_51_n9), .C2(KEY1[51]), .A(KE1_RS_n12), .ZN(
        KE1_RS_SFF_51_n10) );
  INV_X1 KE1_RS_SFF_51_U2 ( .A(RESET), .ZN(KE1_RS_SFF_51_n9) );
  DFF_X1 KE1_RS_SFF_51_Q_reg ( .D(KE1_RS_SFF_51_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[19]), .QN(KE1_RS_SFF_51_n7) );
  OAI21_X1 KE1_RS_SFF_52_U4 ( .B1(KE1_RS_n12), .B2(KE1_RS_SFF_52_n7), .A(
        KE1_RS_SFF_52_n10), .ZN(KE1_RS_SFF_52_n6) );
  OAI221_X1 KE1_RS_SFF_52_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[52]), .C1(
        KE1_RS_SFF_52_n9), .C2(KEY1[52]), .A(KE1_RS_n12), .ZN(
        KE1_RS_SFF_52_n10) );
  INV_X1 KE1_RS_SFF_52_U2 ( .A(RESET), .ZN(KE1_RS_SFF_52_n9) );
  DFF_X1 KE1_RS_SFF_52_Q_reg ( .D(KE1_RS_SFF_52_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[20]), .QN(KE1_RS_SFF_52_n7) );
  OAI21_X1 KE1_RS_SFF_53_U4 ( .B1(KE1_RS_n12), .B2(KE1_RS_SFF_53_n7), .A(
        KE1_RS_SFF_53_n10), .ZN(KE1_RS_SFF_53_n6) );
  OAI221_X1 KE1_RS_SFF_53_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[53]), .C1(
        KE1_RS_SFF_53_n9), .C2(KEY1[53]), .A(KE1_RS_n12), .ZN(
        KE1_RS_SFF_53_n10) );
  INV_X1 KE1_RS_SFF_53_U2 ( .A(RESET), .ZN(KE1_RS_SFF_53_n9) );
  DFF_X1 KE1_RS_SFF_53_Q_reg ( .D(KE1_RS_SFF_53_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[21]), .QN(KE1_RS_SFF_53_n7) );
  OAI21_X1 KE1_RS_SFF_54_U4 ( .B1(KE1_RS_n12), .B2(KE1_RS_SFF_54_n7), .A(
        KE1_RS_SFF_54_n10), .ZN(KE1_RS_SFF_54_n6) );
  OAI221_X1 KE1_RS_SFF_54_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[54]), .C1(
        KE1_RS_SFF_54_n9), .C2(KEY1[54]), .A(KE1_RS_n12), .ZN(
        KE1_RS_SFF_54_n10) );
  INV_X1 KE1_RS_SFF_54_U2 ( .A(RESET), .ZN(KE1_RS_SFF_54_n9) );
  DFF_X1 KE1_RS_SFF_54_Q_reg ( .D(KE1_RS_SFF_54_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[22]), .QN(KE1_RS_SFF_54_n7) );
  OAI21_X1 KE1_RS_SFF_55_U4 ( .B1(KE1_RS_n12), .B2(KE1_RS_SFF_55_n7), .A(
        KE1_RS_SFF_55_n10), .ZN(KE1_RS_SFF_55_n6) );
  OAI221_X1 KE1_RS_SFF_55_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[55]), .C1(
        KE1_RS_SFF_55_n9), .C2(KEY1[55]), .A(KE1_RS_n12), .ZN(
        KE1_RS_SFF_55_n10) );
  INV_X1 KE1_RS_SFF_55_U2 ( .A(RESET), .ZN(KE1_RS_SFF_55_n9) );
  DFF_X1 KE1_RS_SFF_55_Q_reg ( .D(KE1_RS_SFF_55_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[23]), .QN(KE1_RS_SFF_55_n7) );
  OAI21_X1 KE1_RS_SFF_56_U4 ( .B1(KE1_RS_n12), .B2(KE1_RS_SFF_56_n7), .A(
        KE1_RS_SFF_56_n10), .ZN(KE1_RS_SFF_56_n6) );
  OAI221_X1 KE1_RS_SFF_56_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[56]), .C1(
        KE1_RS_SFF_56_n9), .C2(KEY1[56]), .A(KE1_RS_n12), .ZN(
        KE1_RS_SFF_56_n10) );
  INV_X1 KE1_RS_SFF_56_U2 ( .A(RESET), .ZN(KE1_RS_SFF_56_n9) );
  DFF_X1 KE1_RS_SFF_56_Q_reg ( .D(KE1_RS_SFF_56_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[24]), .QN(KE1_RS_SFF_56_n7) );
  OAI21_X1 KE1_RS_SFF_57_U4 ( .B1(KE1_RS_n12), .B2(KE1_RS_SFF_57_n7), .A(
        KE1_RS_SFF_57_n10), .ZN(KE1_RS_SFF_57_n6) );
  OAI221_X1 KE1_RS_SFF_57_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[57]), .C1(
        KE1_RS_SFF_57_n9), .C2(KEY1[57]), .A(KE1_RS_n12), .ZN(
        KE1_RS_SFF_57_n10) );
  INV_X1 KE1_RS_SFF_57_U2 ( .A(RESET), .ZN(KE1_RS_SFF_57_n9) );
  DFF_X1 KE1_RS_SFF_57_Q_reg ( .D(KE1_RS_SFF_57_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[25]), .QN(KE1_RS_SFF_57_n7) );
  OAI21_X1 KE1_RS_SFF_58_U4 ( .B1(KE1_RS_n12), .B2(KE1_RS_SFF_58_n7), .A(
        KE1_RS_SFF_58_n10), .ZN(KE1_RS_SFF_58_n6) );
  OAI221_X1 KE1_RS_SFF_58_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[58]), .C1(
        KE1_RS_SFF_58_n9), .C2(KEY1[58]), .A(KE1_RS_n12), .ZN(
        KE1_RS_SFF_58_n10) );
  INV_X1 KE1_RS_SFF_58_U2 ( .A(RESET), .ZN(KE1_RS_SFF_58_n9) );
  DFF_X1 KE1_RS_SFF_58_Q_reg ( .D(KE1_RS_SFF_58_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[26]), .QN(KE1_RS_SFF_58_n7) );
  OAI21_X1 KE1_RS_SFF_59_U4 ( .B1(KE1_RS_n9), .B2(KE1_RS_SFF_59_n7), .A(
        KE1_RS_SFF_59_n10), .ZN(KE1_RS_SFF_59_n6) );
  OAI221_X1 KE1_RS_SFF_59_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[59]), .C1(
        KE1_RS_SFF_59_n9), .C2(KEY1[59]), .A(KE1_RS_n9), .ZN(KE1_RS_SFF_59_n10) );
  INV_X1 KE1_RS_SFF_59_U2 ( .A(RESET), .ZN(KE1_RS_SFF_59_n9) );
  DFF_X1 KE1_RS_SFF_59_Q_reg ( .D(KE1_RS_SFF_59_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[27]), .QN(KE1_RS_SFF_59_n7) );
  OAI21_X1 KE1_RS_SFF_60_U4 ( .B1(KE1_RS_n8), .B2(KE1_RS_SFF_60_n7), .A(
        KE1_RS_SFF_60_n10), .ZN(KE1_RS_SFF_60_n6) );
  OAI221_X1 KE1_RS_SFF_60_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[60]), .C1(
        KE1_RS_SFF_60_n9), .C2(KEY1[60]), .A(KE1_RS_n8), .ZN(KE1_RS_SFF_60_n10) );
  INV_X1 KE1_RS_SFF_60_U2 ( .A(RESET), .ZN(KE1_RS_SFF_60_n9) );
  DFF_X1 KE1_RS_SFF_60_Q_reg ( .D(KE1_RS_SFF_60_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[28]), .QN(KE1_RS_SFF_60_n7) );
  OAI21_X1 KE1_RS_SFF_61_U4 ( .B1(KE1_RS_n7), .B2(KE1_RS_SFF_61_n7), .A(
        KE1_RS_SFF_61_n10), .ZN(KE1_RS_SFF_61_n6) );
  OAI221_X1 KE1_RS_SFF_61_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[61]), .C1(
        KE1_RS_SFF_61_n9), .C2(KEY1[61]), .A(KE1_RS_n7), .ZN(KE1_RS_SFF_61_n10) );
  INV_X1 KE1_RS_SFF_61_U2 ( .A(RESET), .ZN(KE1_RS_SFF_61_n9) );
  DFF_X1 KE1_RS_SFF_61_Q_reg ( .D(KE1_RS_SFF_61_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[29]), .QN(KE1_RS_SFF_61_n7) );
  OAI21_X1 KE1_RS_SFF_62_U4 ( .B1(KE1_RS_n12), .B2(KE1_RS_SFF_62_n7), .A(
        KE1_RS_SFF_62_n10), .ZN(KE1_RS_SFF_62_n6) );
  OAI221_X1 KE1_RS_SFF_62_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[62]), .C1(
        KE1_RS_SFF_62_n9), .C2(KEY1[62]), .A(KE1_RS_n12), .ZN(
        KE1_RS_SFF_62_n10) );
  INV_X1 KE1_RS_SFF_62_U2 ( .A(RESET), .ZN(KE1_RS_SFF_62_n9) );
  DFF_X1 KE1_RS_SFF_62_Q_reg ( .D(KE1_RS_SFF_62_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[30]), .QN(KE1_RS_SFF_62_n7) );
  OAI21_X1 KE1_RS_SFF_63_U4 ( .B1(KE1_RS_n11), .B2(KE1_RS_SFF_63_n7), .A(
        KE1_RS_SFF_63_n10), .ZN(KE1_RS_SFF_63_n6) );
  OAI221_X1 KE1_RS_SFF_63_U3 ( .B1(RESET), .B2(KE1_KEY_PERM[63]), .C1(
        KE1_RS_SFF_63_n9), .C2(KEY1[63]), .A(KE1_RS_n11), .ZN(
        KE1_RS_SFF_63_n10) );
  INV_X1 KE1_RS_SFF_63_U2 ( .A(RESET), .ZN(KE1_RS_SFF_63_n9) );
  DFF_X1 KE1_RS_SFF_63_Q_reg ( .D(KE1_RS_SFF_63_n6), .CK(CLK), .Q(
        KE1_KEY_PERM[31]), .QN(KE1_RS_SFF_63_n7) );
  BUF_X1 KE2_RS_U6 ( .A(KEY_EN), .Z(KE2_RS_n11) );
  BUF_X1 KE2_RS_U5 ( .A(KEY_EN), .Z(KE2_RS_n10) );
  BUF_X1 KE2_RS_U4 ( .A(KEY_EN), .Z(KE2_RS_n9) );
  BUF_X1 KE2_RS_U3 ( .A(KEY_EN), .Z(KE2_RS_n8) );
  BUF_X1 KE2_RS_U2 ( .A(KEY_EN), .Z(KE2_RS_n7) );
  BUF_X1 KE2_RS_U1 ( .A(KEY_EN), .Z(KE2_RS_n6) );
  OAI21_X1 KE2_RS_SFF_0_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_0_n8), .A(
        KE2_RS_SFF_0_n11), .ZN(KE2_RS_SFF_0_n7) );
  OAI221_X1 KE2_RS_SFF_0_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[0]), .C1(
        KE2_RS_SFF_0_n10), .C2(KEY2[0]), .A(KE2_RS_n8), .ZN(KE2_RS_SFF_0_n11)
         );
  INV_X1 KE2_RS_SFF_0_U2 ( .A(RESET), .ZN(KE2_RS_SFF_0_n10) );
  DFF_X1 KE2_RS_SFF_0_Q_reg ( .D(KE2_RS_SFF_0_n7), .CK(CLK), .Q(
        KE2_KEY_PERM[56]), .QN(KE2_RS_SFF_0_n8) );
  OAI21_X1 KE2_RS_SFF_1_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_1_n8), .A(
        KE2_RS_SFF_1_n11), .ZN(KE2_RS_SFF_1_n7) );
  OAI221_X1 KE2_RS_SFF_1_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[1]), .C1(
        KE2_RS_SFF_1_n10), .C2(KEY2[1]), .A(KE2_RS_n7), .ZN(KE2_RS_SFF_1_n11)
         );
  INV_X1 KE2_RS_SFF_1_U2 ( .A(RESET), .ZN(KE2_RS_SFF_1_n10) );
  DFF_X1 KE2_RS_SFF_1_Q_reg ( .D(KE2_RS_SFF_1_n7), .CK(CLK), .Q(
        KE2_KEY_PERM[57]), .QN(KE2_RS_SFF_1_n8) );
  OAI21_X1 KE2_RS_SFF_2_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_2_n7), .A(
        KE2_RS_SFF_2_n10), .ZN(KE2_RS_SFF_2_n6) );
  OAI221_X1 KE2_RS_SFF_2_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[2]), .C1(
        KE2_RS_SFF_2_n9), .C2(KEY2[2]), .A(KE2_RS_n6), .ZN(KE2_RS_SFF_2_n10)
         );
  INV_X1 KE2_RS_SFF_2_U2 ( .A(RESET), .ZN(KE2_RS_SFF_2_n9) );
  DFF_X1 KE2_RS_SFF_2_Q_reg ( .D(KE2_RS_SFF_2_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[58]), .QN(KE2_RS_SFF_2_n7) );
  OAI21_X1 KE2_RS_SFF_3_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_3_n7), .A(
        KE2_RS_SFF_3_n10), .ZN(KE2_RS_SFF_3_n6) );
  OAI221_X1 KE2_RS_SFF_3_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[3]), .C1(
        KE2_RS_SFF_3_n9), .C2(KEY2[3]), .A(KE2_RS_n6), .ZN(KE2_RS_SFF_3_n10)
         );
  INV_X1 KE2_RS_SFF_3_U2 ( .A(RESET), .ZN(KE2_RS_SFF_3_n9) );
  DFF_X1 KE2_RS_SFF_3_Q_reg ( .D(KE2_RS_SFF_3_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[59]), .QN(KE2_RS_SFF_3_n7) );
  OAI21_X1 KE2_RS_SFF_4_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_4_n7), .A(
        KE2_RS_SFF_4_n10), .ZN(KE2_RS_SFF_4_n6) );
  OAI221_X1 KE2_RS_SFF_4_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[4]), .C1(
        KE2_RS_SFF_4_n9), .C2(KEY2[4]), .A(KE2_RS_n6), .ZN(KE2_RS_SFF_4_n10)
         );
  INV_X1 KE2_RS_SFF_4_U2 ( .A(RESET), .ZN(KE2_RS_SFF_4_n9) );
  DFF_X1 KE2_RS_SFF_4_Q_reg ( .D(KE2_RS_SFF_4_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[40]), .QN(KE2_RS_SFF_4_n7) );
  OAI21_X1 KE2_RS_SFF_5_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_5_n7), .A(
        KE2_RS_SFF_5_n10), .ZN(KE2_RS_SFF_5_n6) );
  OAI221_X1 KE2_RS_SFF_5_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[5]), .C1(
        KE2_RS_SFF_5_n9), .C2(KEY2[5]), .A(KE2_RS_n6), .ZN(KE2_RS_SFF_5_n10)
         );
  INV_X1 KE2_RS_SFF_5_U2 ( .A(RESET), .ZN(KE2_RS_SFF_5_n9) );
  DFF_X1 KE2_RS_SFF_5_Q_reg ( .D(KE2_RS_SFF_5_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[41]), .QN(KE2_RS_SFF_5_n7) );
  OAI21_X1 KE2_RS_SFF_6_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_6_n7), .A(
        KE2_RS_SFF_6_n10), .ZN(KE2_RS_SFF_6_n6) );
  OAI221_X1 KE2_RS_SFF_6_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[6]), .C1(
        KE2_RS_SFF_6_n9), .C2(KEY2[6]), .A(KE2_RS_n6), .ZN(KE2_RS_SFF_6_n10)
         );
  INV_X1 KE2_RS_SFF_6_U2 ( .A(RESET), .ZN(KE2_RS_SFF_6_n9) );
  DFF_X1 KE2_RS_SFF_6_Q_reg ( .D(KE2_RS_SFF_6_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[42]), .QN(KE2_RS_SFF_6_n7) );
  OAI21_X1 KE2_RS_SFF_7_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_7_n7), .A(
        KE2_RS_SFF_7_n10), .ZN(KE2_RS_SFF_7_n6) );
  OAI221_X1 KE2_RS_SFF_7_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[7]), .C1(
        KE2_RS_SFF_7_n9), .C2(KEY2[7]), .A(KE2_RS_n6), .ZN(KE2_RS_SFF_7_n10)
         );
  INV_X1 KE2_RS_SFF_7_U2 ( .A(RESET), .ZN(KE2_RS_SFF_7_n9) );
  DFF_X1 KE2_RS_SFF_7_Q_reg ( .D(KE2_RS_SFF_7_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[43]), .QN(KE2_RS_SFF_7_n7) );
  OAI21_X1 KE2_RS_SFF_8_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_8_n7), .A(
        KE2_RS_SFF_8_n10), .ZN(KE2_RS_SFF_8_n6) );
  OAI221_X1 KE2_RS_SFF_8_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[8]), .C1(
        KE2_RS_SFF_8_n9), .C2(KEY2[8]), .A(KE2_RS_n6), .ZN(KE2_RS_SFF_8_n10)
         );
  INV_X1 KE2_RS_SFF_8_U2 ( .A(RESET), .ZN(KE2_RS_SFF_8_n9) );
  DFF_X1 KE2_RS_SFF_8_Q_reg ( .D(KE2_RS_SFF_8_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[48]), .QN(KE2_RS_SFF_8_n7) );
  OAI21_X1 KE2_RS_SFF_9_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_9_n7), .A(
        KE2_RS_SFF_9_n10), .ZN(KE2_RS_SFF_9_n6) );
  OAI221_X1 KE2_RS_SFF_9_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[9]), .C1(
        KE2_RS_SFF_9_n9), .C2(KEY2[9]), .A(KE2_RS_n6), .ZN(KE2_RS_SFF_9_n10)
         );
  INV_X1 KE2_RS_SFF_9_U2 ( .A(RESET), .ZN(KE2_RS_SFF_9_n9) );
  DFF_X1 KE2_RS_SFF_9_Q_reg ( .D(KE2_RS_SFF_9_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[49]), .QN(KE2_RS_SFF_9_n7) );
  OAI21_X1 KE2_RS_SFF_10_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_10_n7), .A(
        KE2_RS_SFF_10_n10), .ZN(KE2_RS_SFF_10_n6) );
  OAI221_X1 KE2_RS_SFF_10_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[10]), .C1(
        KE2_RS_SFF_10_n9), .C2(KEY2[10]), .A(KE2_RS_n7), .ZN(KE2_RS_SFF_10_n10) );
  INV_X1 KE2_RS_SFF_10_U2 ( .A(RESET), .ZN(KE2_RS_SFF_10_n9) );
  DFF_X1 KE2_RS_SFF_10_Q_reg ( .D(KE2_RS_SFF_10_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[50]), .QN(KE2_RS_SFF_10_n7) );
  OAI21_X1 KE2_RS_SFF_11_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_11_n7), .A(
        KE2_RS_SFF_11_n10), .ZN(KE2_RS_SFF_11_n6) );
  OAI221_X1 KE2_RS_SFF_11_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[11]), .C1(
        KE2_RS_SFF_11_n9), .C2(KEY2[11]), .A(KE2_RS_n7), .ZN(KE2_RS_SFF_11_n10) );
  INV_X1 KE2_RS_SFF_11_U2 ( .A(RESET), .ZN(KE2_RS_SFF_11_n9) );
  DFF_X1 KE2_RS_SFF_11_Q_reg ( .D(KE2_RS_SFF_11_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[51]), .QN(KE2_RS_SFF_11_n7) );
  OAI21_X1 KE2_RS_SFF_12_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_12_n8), .A(
        KE2_RS_SFF_12_n11), .ZN(KE2_RS_SFF_12_n7) );
  OAI221_X1 KE2_RS_SFF_12_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[12]), .C1(
        KE2_RS_SFF_12_n10), .C2(KEY2[12]), .A(KE2_RS_n6), .ZN(
        KE2_RS_SFF_12_n11) );
  INV_X1 KE2_RS_SFF_12_U2 ( .A(RESET), .ZN(KE2_RS_SFF_12_n10) );
  DFF_X1 KE2_RS_SFF_12_Q_reg ( .D(KE2_RS_SFF_12_n7), .CK(CLK), .Q(
        KE2_KEY_PERM[36]), .QN(KE2_RS_SFF_12_n8) );
  OAI21_X1 KE2_RS_SFF_13_U4 ( .B1(KE2_RS_n11), .B2(KE2_RS_SFF_13_n8), .A(
        KE2_RS_SFF_13_n11), .ZN(KE2_RS_SFF_13_n7) );
  OAI221_X1 KE2_RS_SFF_13_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[13]), .C1(
        KE2_RS_SFF_13_n10), .C2(KEY2[13]), .A(KE2_RS_n11), .ZN(
        KE2_RS_SFF_13_n11) );
  INV_X1 KE2_RS_SFF_13_U2 ( .A(RESET), .ZN(KE2_RS_SFF_13_n10) );
  DFF_X1 KE2_RS_SFF_13_Q_reg ( .D(KE2_RS_SFF_13_n7), .CK(CLK), .Q(
        KE2_KEY_PERM[37]), .QN(KE2_RS_SFF_13_n8) );
  OAI21_X1 KE2_RS_SFF_14_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_14_n7), .A(
        KE2_RS_SFF_14_n10), .ZN(KE2_RS_SFF_14_n6) );
  OAI221_X1 KE2_RS_SFF_14_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[14]), .C1(
        KE2_RS_SFF_14_n9), .C2(KEY2[14]), .A(KE2_RS_n7), .ZN(KE2_RS_SFF_14_n10) );
  INV_X1 KE2_RS_SFF_14_U2 ( .A(RESET), .ZN(KE2_RS_SFF_14_n9) );
  DFF_X1 KE2_RS_SFF_14_Q_reg ( .D(KE2_RS_SFF_14_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[38]), .QN(KE2_RS_SFF_14_n7) );
  OAI21_X1 KE2_RS_SFF_15_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_15_n7), .A(
        KE2_RS_SFF_15_n10), .ZN(KE2_RS_SFF_15_n6) );
  OAI221_X1 KE2_RS_SFF_15_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[15]), .C1(
        KE2_RS_SFF_15_n9), .C2(KEY2[15]), .A(KE2_RS_n7), .ZN(KE2_RS_SFF_15_n10) );
  INV_X1 KE2_RS_SFF_15_U2 ( .A(RESET), .ZN(KE2_RS_SFF_15_n9) );
  DFF_X1 KE2_RS_SFF_15_Q_reg ( .D(KE2_RS_SFF_15_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[39]), .QN(KE2_RS_SFF_15_n7) );
  OAI21_X1 KE2_RS_SFF_16_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_16_n7), .A(
        KE2_RS_SFF_16_n10), .ZN(KE2_RS_SFF_16_n6) );
  OAI221_X1 KE2_RS_SFF_16_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[16]), .C1(
        KE2_RS_SFF_16_n9), .C2(KEY2[16]), .A(KE2_RS_n7), .ZN(KE2_RS_SFF_16_n10) );
  INV_X1 KE2_RS_SFF_16_U2 ( .A(RESET), .ZN(KE2_RS_SFF_16_n9) );
  DFF_X1 KE2_RS_SFF_16_Q_reg ( .D(KE2_RS_SFF_16_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[32]), .QN(KE2_RS_SFF_16_n7) );
  OAI21_X1 KE2_RS_SFF_17_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_17_n7), .A(
        KE2_RS_SFF_17_n10), .ZN(KE2_RS_SFF_17_n6) );
  OAI221_X1 KE2_RS_SFF_17_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[17]), .C1(
        KE2_RS_SFF_17_n9), .C2(KEY2[17]), .A(KE2_RS_n7), .ZN(KE2_RS_SFF_17_n10) );
  INV_X1 KE2_RS_SFF_17_U2 ( .A(RESET), .ZN(KE2_RS_SFF_17_n9) );
  DFF_X1 KE2_RS_SFF_17_Q_reg ( .D(KE2_RS_SFF_17_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[33]), .QN(KE2_RS_SFF_17_n7) );
  OAI21_X1 KE2_RS_SFF_18_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_18_n7), .A(
        KE2_RS_SFF_18_n10), .ZN(KE2_RS_SFF_18_n6) );
  OAI221_X1 KE2_RS_SFF_18_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[18]), .C1(
        KE2_RS_SFF_18_n9), .C2(KEY2[18]), .A(KE2_RS_n7), .ZN(KE2_RS_SFF_18_n10) );
  INV_X1 KE2_RS_SFF_18_U2 ( .A(RESET), .ZN(KE2_RS_SFF_18_n9) );
  DFF_X1 KE2_RS_SFF_18_Q_reg ( .D(KE2_RS_SFF_18_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[34]), .QN(KE2_RS_SFF_18_n7) );
  OAI21_X1 KE2_RS_SFF_19_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_19_n7), .A(
        KE2_RS_SFF_19_n10), .ZN(KE2_RS_SFF_19_n6) );
  OAI221_X1 KE2_RS_SFF_19_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[19]), .C1(
        KE2_RS_SFF_19_n9), .C2(KEY2[19]), .A(KE2_RS_n7), .ZN(KE2_RS_SFF_19_n10) );
  INV_X1 KE2_RS_SFF_19_U2 ( .A(RESET), .ZN(KE2_RS_SFF_19_n9) );
  DFF_X1 KE2_RS_SFF_19_Q_reg ( .D(KE2_RS_SFF_19_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[35]), .QN(KE2_RS_SFF_19_n7) );
  OAI21_X1 KE2_RS_SFF_20_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_20_n7), .A(
        KE2_RS_SFF_20_n10), .ZN(KE2_RS_SFF_20_n6) );
  OAI221_X1 KE2_RS_SFF_20_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[20]), .C1(
        KE2_RS_SFF_20_n9), .C2(KEY2[20]), .A(KE2_RS_n8), .ZN(KE2_RS_SFF_20_n10) );
  INV_X1 KE2_RS_SFF_20_U2 ( .A(RESET), .ZN(KE2_RS_SFF_20_n9) );
  DFF_X1 KE2_RS_SFF_20_Q_reg ( .D(KE2_RS_SFF_20_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[44]), .QN(KE2_RS_SFF_20_n7) );
  OAI21_X1 KE2_RS_SFF_21_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_21_n7), .A(
        KE2_RS_SFF_21_n10), .ZN(KE2_RS_SFF_21_n6) );
  OAI221_X1 KE2_RS_SFF_21_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[21]), .C1(
        KE2_RS_SFF_21_n9), .C2(KEY2[21]), .A(KE2_RS_n8), .ZN(KE2_RS_SFF_21_n10) );
  INV_X1 KE2_RS_SFF_21_U2 ( .A(RESET), .ZN(KE2_RS_SFF_21_n9) );
  DFF_X1 KE2_RS_SFF_21_Q_reg ( .D(KE2_RS_SFF_21_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[45]), .QN(KE2_RS_SFF_21_n7) );
  OAI21_X1 KE2_RS_SFF_22_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_22_n7), .A(
        KE2_RS_SFF_22_n10), .ZN(KE2_RS_SFF_22_n6) );
  OAI221_X1 KE2_RS_SFF_22_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[22]), .C1(
        KE2_RS_SFF_22_n9), .C2(KEY2[22]), .A(KE2_RS_n8), .ZN(KE2_RS_SFF_22_n10) );
  INV_X1 KE2_RS_SFF_22_U2 ( .A(RESET), .ZN(KE2_RS_SFF_22_n9) );
  DFF_X1 KE2_RS_SFF_22_Q_reg ( .D(KE2_RS_SFF_22_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[46]), .QN(KE2_RS_SFF_22_n7) );
  OAI21_X1 KE2_RS_SFF_23_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_23_n7), .A(
        KE2_RS_SFF_23_n10), .ZN(KE2_RS_SFF_23_n6) );
  OAI221_X1 KE2_RS_SFF_23_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[23]), .C1(
        KE2_RS_SFF_23_n9), .C2(KEY2[23]), .A(KE2_RS_n8), .ZN(KE2_RS_SFF_23_n10) );
  INV_X1 KE2_RS_SFF_23_U2 ( .A(RESET), .ZN(KE2_RS_SFF_23_n9) );
  DFF_X1 KE2_RS_SFF_23_Q_reg ( .D(KE2_RS_SFF_23_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[47]), .QN(KE2_RS_SFF_23_n7) );
  OAI21_X1 KE2_RS_SFF_24_U4 ( .B1(KE2_RS_n10), .B2(KE2_RS_SFF_24_n8), .A(
        KE2_RS_SFF_24_n11), .ZN(KE2_RS_SFF_24_n7) );
  OAI221_X1 KE2_RS_SFF_24_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[24]), .C1(
        KE2_RS_SFF_24_n10), .C2(KEY2[24]), .A(KE2_RS_n10), .ZN(
        KE2_RS_SFF_24_n11) );
  INV_X1 KE2_RS_SFF_24_U2 ( .A(RESET), .ZN(KE2_RS_SFF_24_n10) );
  DFF_X1 KE2_RS_SFF_24_Q_reg ( .D(KE2_RS_SFF_24_n7), .CK(CLK), .Q(
        KE2_KEY_PERM[60]), .QN(KE2_RS_SFF_24_n8) );
  OAI21_X1 KE2_RS_SFF_25_U4 ( .B1(KE2_RS_n9), .B2(KE2_RS_SFF_25_n8), .A(
        KE2_RS_SFF_25_n11), .ZN(KE2_RS_SFF_25_n7) );
  OAI221_X1 KE2_RS_SFF_25_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[25]), .C1(
        KE2_RS_SFF_25_n10), .C2(KEY2[25]), .A(KE2_RS_n9), .ZN(
        KE2_RS_SFF_25_n11) );
  INV_X1 KE2_RS_SFF_25_U2 ( .A(RESET), .ZN(KE2_RS_SFF_25_n10) );
  DFF_X1 KE2_RS_SFF_25_Q_reg ( .D(KE2_RS_SFF_25_n7), .CK(CLK), .Q(
        KE2_KEY_PERM[61]), .QN(KE2_RS_SFF_25_n8) );
  OAI21_X1 KE2_RS_SFF_26_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_26_n7), .A(
        KE2_RS_SFF_26_n10), .ZN(KE2_RS_SFF_26_n6) );
  OAI221_X1 KE2_RS_SFF_26_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[26]), .C1(
        KE2_RS_SFF_26_n9), .C2(KEY2[26]), .A(KE2_RS_n8), .ZN(KE2_RS_SFF_26_n10) );
  INV_X1 KE2_RS_SFF_26_U2 ( .A(RESET), .ZN(KE2_RS_SFF_26_n9) );
  DFF_X1 KE2_RS_SFF_26_Q_reg ( .D(KE2_RS_SFF_26_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[62]), .QN(KE2_RS_SFF_26_n7) );
  OAI21_X1 KE2_RS_SFF_27_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_27_n7), .A(
        KE2_RS_SFF_27_n10), .ZN(KE2_RS_SFF_27_n6) );
  OAI221_X1 KE2_RS_SFF_27_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[27]), .C1(
        KE2_RS_SFF_27_n9), .C2(KEY2[27]), .A(KE2_RS_n8), .ZN(KE2_RS_SFF_27_n10) );
  INV_X1 KE2_RS_SFF_27_U2 ( .A(RESET), .ZN(KE2_RS_SFF_27_n9) );
  DFF_X1 KE2_RS_SFF_27_Q_reg ( .D(KE2_RS_SFF_27_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[63]), .QN(KE2_RS_SFF_27_n7) );
  OAI21_X1 KE2_RS_SFF_28_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_28_n7), .A(
        KE2_RS_SFF_28_n10), .ZN(KE2_RS_SFF_28_n6) );
  OAI221_X1 KE2_RS_SFF_28_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[28]), .C1(
        KE2_RS_SFF_28_n9), .C2(KEY2[28]), .A(KE2_RS_n8), .ZN(KE2_RS_SFF_28_n10) );
  INV_X1 KE2_RS_SFF_28_U2 ( .A(RESET), .ZN(KE2_RS_SFF_28_n9) );
  DFF_X1 KE2_RS_SFF_28_Q_reg ( .D(KE2_RS_SFF_28_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[52]), .QN(KE2_RS_SFF_28_n7) );
  OAI21_X1 KE2_RS_SFF_29_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_29_n7), .A(
        KE2_RS_SFF_29_n10), .ZN(KE2_RS_SFF_29_n6) );
  OAI221_X1 KE2_RS_SFF_29_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[29]), .C1(
        KE2_RS_SFF_29_n9), .C2(KEY2[29]), .A(KE2_RS_n8), .ZN(KE2_RS_SFF_29_n10) );
  INV_X1 KE2_RS_SFF_29_U2 ( .A(RESET), .ZN(KE2_RS_SFF_29_n9) );
  DFF_X1 KE2_RS_SFF_29_Q_reg ( .D(KE2_RS_SFF_29_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[53]), .QN(KE2_RS_SFF_29_n7) );
  OAI21_X1 KE2_RS_SFF_30_U4 ( .B1(KE2_RS_n9), .B2(KE2_RS_SFF_30_n7), .A(
        KE2_RS_SFF_30_n10), .ZN(KE2_RS_SFF_30_n6) );
  OAI221_X1 KE2_RS_SFF_30_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[30]), .C1(
        KE2_RS_SFF_30_n9), .C2(KEY2[30]), .A(KE2_RS_n9), .ZN(KE2_RS_SFF_30_n10) );
  INV_X1 KE2_RS_SFF_30_U2 ( .A(RESET), .ZN(KE2_RS_SFF_30_n9) );
  DFF_X1 KE2_RS_SFF_30_Q_reg ( .D(KE2_RS_SFF_30_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[54]), .QN(KE2_RS_SFF_30_n7) );
  OAI21_X1 KE2_RS_SFF_31_U4 ( .B1(KE2_RS_n9), .B2(KE2_RS_SFF_31_n7), .A(
        KE2_RS_SFF_31_n10), .ZN(KE2_RS_SFF_31_n6) );
  OAI221_X1 KE2_RS_SFF_31_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[31]), .C1(
        KE2_RS_SFF_31_n9), .C2(KEY2[31]), .A(KE2_RS_n9), .ZN(KE2_RS_SFF_31_n10) );
  INV_X1 KE2_RS_SFF_31_U2 ( .A(RESET), .ZN(KE2_RS_SFF_31_n9) );
  DFF_X1 KE2_RS_SFF_31_Q_reg ( .D(KE2_RS_SFF_31_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[55]), .QN(KE2_RS_SFF_31_n7) );
  OAI21_X1 KE2_RS_SFF_32_U4 ( .B1(KE2_RS_n9), .B2(KE2_RS_SFF_32_n7), .A(
        KE2_RS_SFF_32_n10), .ZN(KE2_RS_SFF_32_n6) );
  OAI221_X1 KE2_RS_SFF_32_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[32]), .C1(
        KE2_RS_SFF_32_n9), .C2(KEY2[32]), .A(KE2_RS_n9), .ZN(KE2_RS_SFF_32_n10) );
  INV_X1 KE2_RS_SFF_32_U2 ( .A(RESET), .ZN(KE2_RS_SFF_32_n9) );
  DFF_X1 KE2_RS_SFF_32_Q_reg ( .D(KE2_RS_SFF_32_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[0]), .QN(KE2_RS_SFF_32_n7) );
  OAI21_X1 KE2_RS_SFF_33_U4 ( .B1(KE2_RS_n9), .B2(KE2_RS_SFF_33_n7), .A(
        KE2_RS_SFF_33_n10), .ZN(KE2_RS_SFF_33_n6) );
  OAI221_X1 KE2_RS_SFF_33_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[33]), .C1(
        KE2_RS_SFF_33_n9), .C2(KEY2[33]), .A(KE2_RS_n9), .ZN(KE2_RS_SFF_33_n10) );
  INV_X1 KE2_RS_SFF_33_U2 ( .A(RESET), .ZN(KE2_RS_SFF_33_n9) );
  DFF_X1 KE2_RS_SFF_33_Q_reg ( .D(KE2_RS_SFF_33_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[1]), .QN(KE2_RS_SFF_33_n7) );
  OAI21_X1 KE2_RS_SFF_34_U4 ( .B1(KE2_RS_n9), .B2(KE2_RS_SFF_34_n7), .A(
        KE2_RS_SFF_34_n10), .ZN(KE2_RS_SFF_34_n6) );
  OAI221_X1 KE2_RS_SFF_34_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[34]), .C1(
        KE2_RS_SFF_34_n9), .C2(KEY2[34]), .A(KE2_RS_n9), .ZN(KE2_RS_SFF_34_n10) );
  INV_X1 KE2_RS_SFF_34_U2 ( .A(RESET), .ZN(KE2_RS_SFF_34_n9) );
  DFF_X1 KE2_RS_SFF_34_Q_reg ( .D(KE2_RS_SFF_34_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[2]), .QN(KE2_RS_SFF_34_n7) );
  OAI21_X1 KE2_RS_SFF_35_U4 ( .B1(KE2_RS_n9), .B2(KE2_RS_SFF_35_n7), .A(
        KE2_RS_SFF_35_n10), .ZN(KE2_RS_SFF_35_n6) );
  OAI221_X1 KE2_RS_SFF_35_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[35]), .C1(
        KE2_RS_SFF_35_n9), .C2(KEY2[35]), .A(KE2_RS_n9), .ZN(KE2_RS_SFF_35_n10) );
  INV_X1 KE2_RS_SFF_35_U2 ( .A(RESET), .ZN(KE2_RS_SFF_35_n9) );
  DFF_X1 KE2_RS_SFF_35_Q_reg ( .D(KE2_RS_SFF_35_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[3]), .QN(KE2_RS_SFF_35_n7) );
  OAI21_X1 KE2_RS_SFF_36_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_36_n8), .A(
        KE2_RS_SFF_36_n11), .ZN(KE2_RS_SFF_36_n7) );
  OAI221_X1 KE2_RS_SFF_36_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[36]), .C1(
        KE2_RS_SFF_36_n10), .C2(KEY2[36]), .A(KE2_RS_n8), .ZN(
        KE2_RS_SFF_36_n11) );
  INV_X1 KE2_RS_SFF_36_U2 ( .A(RESET), .ZN(KE2_RS_SFF_36_n10) );
  DFF_X1 KE2_RS_SFF_36_Q_reg ( .D(KE2_RS_SFF_36_n7), .CK(CLK), .Q(
        KE2_KEY_PERM[4]), .QN(KE2_RS_SFF_36_n8) );
  OAI21_X1 KE2_RS_SFF_37_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_37_n8), .A(
        KE2_RS_SFF_37_n11), .ZN(KE2_RS_SFF_37_n7) );
  OAI221_X1 KE2_RS_SFF_37_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[37]), .C1(
        KE2_RS_SFF_37_n10), .C2(KEY2[37]), .A(KE2_RS_n7), .ZN(
        KE2_RS_SFF_37_n11) );
  INV_X1 KE2_RS_SFF_37_U2 ( .A(RESET), .ZN(KE2_RS_SFF_37_n10) );
  DFF_X1 KE2_RS_SFF_37_Q_reg ( .D(KE2_RS_SFF_37_n7), .CK(CLK), .Q(
        KE2_KEY_PERM[5]), .QN(KE2_RS_SFF_37_n8) );
  OAI21_X1 KE2_RS_SFF_38_U4 ( .B1(KE2_RS_n9), .B2(KE2_RS_SFF_38_n7), .A(
        KE2_RS_SFF_38_n10), .ZN(KE2_RS_SFF_38_n6) );
  OAI221_X1 KE2_RS_SFF_38_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[38]), .C1(
        KE2_RS_SFF_38_n9), .C2(KEY2[38]), .A(KE2_RS_n9), .ZN(KE2_RS_SFF_38_n10) );
  INV_X1 KE2_RS_SFF_38_U2 ( .A(RESET), .ZN(KE2_RS_SFF_38_n9) );
  DFF_X1 KE2_RS_SFF_38_Q_reg ( .D(KE2_RS_SFF_38_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[6]), .QN(KE2_RS_SFF_38_n7) );
  OAI21_X1 KE2_RS_SFF_39_U4 ( .B1(KE2_RS_n9), .B2(KE2_RS_SFF_39_n7), .A(
        KE2_RS_SFF_39_n10), .ZN(KE2_RS_SFF_39_n6) );
  OAI221_X1 KE2_RS_SFF_39_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[39]), .C1(
        KE2_RS_SFF_39_n9), .C2(KEY2[39]), .A(KE2_RS_n9), .ZN(KE2_RS_SFF_39_n10) );
  INV_X1 KE2_RS_SFF_39_U2 ( .A(RESET), .ZN(KE2_RS_SFF_39_n9) );
  DFF_X1 KE2_RS_SFF_39_Q_reg ( .D(KE2_RS_SFF_39_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[7]), .QN(KE2_RS_SFF_39_n7) );
  OAI21_X1 KE2_RS_SFF_40_U4 ( .B1(KE2_RS_n10), .B2(KE2_RS_SFF_40_n7), .A(
        KE2_RS_SFF_40_n10), .ZN(KE2_RS_SFF_40_n6) );
  OAI221_X1 KE2_RS_SFF_40_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[40]), .C1(
        KE2_RS_SFF_40_n9), .C2(KEY2[40]), .A(KE2_RS_n10), .ZN(
        KE2_RS_SFF_40_n10) );
  INV_X1 KE2_RS_SFF_40_U2 ( .A(RESET), .ZN(KE2_RS_SFF_40_n9) );
  DFF_X1 KE2_RS_SFF_40_Q_reg ( .D(KE2_RS_SFF_40_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[8]), .QN(KE2_RS_SFF_40_n7) );
  OAI21_X1 KE2_RS_SFF_41_U4 ( .B1(KE2_RS_n10), .B2(KE2_RS_SFF_41_n7), .A(
        KE2_RS_SFF_41_n10), .ZN(KE2_RS_SFF_41_n6) );
  OAI221_X1 KE2_RS_SFF_41_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[41]), .C1(
        KE2_RS_SFF_41_n9), .C2(KEY2[41]), .A(KE2_RS_n10), .ZN(
        KE2_RS_SFF_41_n10) );
  INV_X1 KE2_RS_SFF_41_U2 ( .A(RESET), .ZN(KE2_RS_SFF_41_n9) );
  DFF_X1 KE2_RS_SFF_41_Q_reg ( .D(KE2_RS_SFF_41_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[9]), .QN(KE2_RS_SFF_41_n7) );
  OAI21_X1 KE2_RS_SFF_42_U4 ( .B1(KE2_RS_n10), .B2(KE2_RS_SFF_42_n7), .A(
        KE2_RS_SFF_42_n10), .ZN(KE2_RS_SFF_42_n6) );
  OAI221_X1 KE2_RS_SFF_42_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[42]), .C1(
        KE2_RS_SFF_42_n9), .C2(KEY2[42]), .A(KE2_RS_n10), .ZN(
        KE2_RS_SFF_42_n10) );
  INV_X1 KE2_RS_SFF_42_U2 ( .A(RESET), .ZN(KE2_RS_SFF_42_n9) );
  DFF_X1 KE2_RS_SFF_42_Q_reg ( .D(KE2_RS_SFF_42_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[10]), .QN(KE2_RS_SFF_42_n7) );
  OAI21_X1 KE2_RS_SFF_43_U4 ( .B1(KE2_RS_n10), .B2(KE2_RS_SFF_43_n7), .A(
        KE2_RS_SFF_43_n10), .ZN(KE2_RS_SFF_43_n6) );
  OAI221_X1 KE2_RS_SFF_43_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[43]), .C1(
        KE2_RS_SFF_43_n9), .C2(KEY2[43]), .A(KE2_RS_n10), .ZN(
        KE2_RS_SFF_43_n10) );
  INV_X1 KE2_RS_SFF_43_U2 ( .A(RESET), .ZN(KE2_RS_SFF_43_n9) );
  DFF_X1 KE2_RS_SFF_43_Q_reg ( .D(KE2_RS_SFF_43_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[11]), .QN(KE2_RS_SFF_43_n7) );
  OAI21_X1 KE2_RS_SFF_44_U4 ( .B1(KE2_RS_n10), .B2(KE2_RS_SFF_44_n7), .A(
        KE2_RS_SFF_44_n10), .ZN(KE2_RS_SFF_44_n6) );
  OAI221_X1 KE2_RS_SFF_44_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[44]), .C1(
        KE2_RS_SFF_44_n9), .C2(KEY2[44]), .A(KE2_RS_n10), .ZN(
        KE2_RS_SFF_44_n10) );
  INV_X1 KE2_RS_SFF_44_U2 ( .A(RESET), .ZN(KE2_RS_SFF_44_n9) );
  DFF_X1 KE2_RS_SFF_44_Q_reg ( .D(KE2_RS_SFF_44_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[12]), .QN(KE2_RS_SFF_44_n7) );
  OAI21_X1 KE2_RS_SFF_45_U4 ( .B1(KE2_RS_n10), .B2(KE2_RS_SFF_45_n7), .A(
        KE2_RS_SFF_45_n10), .ZN(KE2_RS_SFF_45_n6) );
  OAI221_X1 KE2_RS_SFF_45_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[45]), .C1(
        KE2_RS_SFF_45_n9), .C2(KEY2[45]), .A(KE2_RS_n10), .ZN(
        KE2_RS_SFF_45_n10) );
  INV_X1 KE2_RS_SFF_45_U2 ( .A(RESET), .ZN(KE2_RS_SFF_45_n9) );
  DFF_X1 KE2_RS_SFF_45_Q_reg ( .D(KE2_RS_SFF_45_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[13]), .QN(KE2_RS_SFF_45_n7) );
  OAI21_X1 KE2_RS_SFF_46_U4 ( .B1(KE2_RS_n10), .B2(KE2_RS_SFF_46_n7), .A(
        KE2_RS_SFF_46_n10), .ZN(KE2_RS_SFF_46_n6) );
  OAI221_X1 KE2_RS_SFF_46_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[46]), .C1(
        KE2_RS_SFF_46_n9), .C2(KEY2[46]), .A(KE2_RS_n10), .ZN(
        KE2_RS_SFF_46_n10) );
  INV_X1 KE2_RS_SFF_46_U2 ( .A(RESET), .ZN(KE2_RS_SFF_46_n9) );
  DFF_X1 KE2_RS_SFF_46_Q_reg ( .D(KE2_RS_SFF_46_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[14]), .QN(KE2_RS_SFF_46_n7) );
  OAI21_X1 KE2_RS_SFF_47_U4 ( .B1(KE2_RS_n10), .B2(KE2_RS_SFF_47_n7), .A(
        KE2_RS_SFF_47_n10), .ZN(KE2_RS_SFF_47_n6) );
  OAI221_X1 KE2_RS_SFF_47_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[47]), .C1(
        KE2_RS_SFF_47_n9), .C2(KEY2[47]), .A(KE2_RS_n10), .ZN(
        KE2_RS_SFF_47_n10) );
  INV_X1 KE2_RS_SFF_47_U2 ( .A(RESET), .ZN(KE2_RS_SFF_47_n9) );
  DFF_X1 KE2_RS_SFF_47_Q_reg ( .D(KE2_RS_SFF_47_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[15]), .QN(KE2_RS_SFF_47_n7) );
  OAI21_X1 KE2_RS_SFF_48_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_48_n8), .A(
        KE2_RS_SFF_48_n11), .ZN(KE2_RS_SFF_48_n7) );
  OAI221_X1 KE2_RS_SFF_48_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[48]), .C1(
        KE2_RS_SFF_48_n10), .C2(KEY2[48]), .A(KE2_RS_n6), .ZN(
        KE2_RS_SFF_48_n11) );
  INV_X1 KE2_RS_SFF_48_U2 ( .A(RESET), .ZN(KE2_RS_SFF_48_n10) );
  DFF_X1 KE2_RS_SFF_48_Q_reg ( .D(KE2_RS_SFF_48_n7), .CK(CLK), .Q(
        KE2_KEY_PERM[16]), .QN(KE2_RS_SFF_48_n8) );
  OAI21_X1 KE2_RS_SFF_49_U4 ( .B1(KEY_EN), .B2(KE2_RS_SFF_49_n8), .A(
        KE2_RS_SFF_49_n11), .ZN(KE2_RS_SFF_49_n7) );
  OAI221_X1 KE2_RS_SFF_49_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[49]), .C1(
        KE2_RS_SFF_49_n10), .C2(KEY2[49]), .A(KEY_EN), .ZN(KE2_RS_SFF_49_n11)
         );
  INV_X1 KE2_RS_SFF_49_U2 ( .A(RESET), .ZN(KE2_RS_SFF_49_n10) );
  DFF_X1 KE2_RS_SFF_49_Q_reg ( .D(KE2_RS_SFF_49_n7), .CK(CLK), .Q(
        KE2_KEY_PERM[17]), .QN(KE2_RS_SFF_49_n8) );
  OAI21_X1 KE2_RS_SFF_50_U4 ( .B1(KE2_RS_n11), .B2(KE2_RS_SFF_50_n7), .A(
        KE2_RS_SFF_50_n10), .ZN(KE2_RS_SFF_50_n6) );
  OAI221_X1 KE2_RS_SFF_50_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[50]), .C1(
        KE2_RS_SFF_50_n9), .C2(KEY2[50]), .A(KE2_RS_n11), .ZN(
        KE2_RS_SFF_50_n10) );
  INV_X1 KE2_RS_SFF_50_U2 ( .A(RESET), .ZN(KE2_RS_SFF_50_n9) );
  DFF_X1 KE2_RS_SFF_50_Q_reg ( .D(KE2_RS_SFF_50_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[18]), .QN(KE2_RS_SFF_50_n7) );
  OAI21_X1 KE2_RS_SFF_51_U4 ( .B1(KE2_RS_n11), .B2(KE2_RS_SFF_51_n7), .A(
        KE2_RS_SFF_51_n10), .ZN(KE2_RS_SFF_51_n6) );
  OAI221_X1 KE2_RS_SFF_51_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[51]), .C1(
        KE2_RS_SFF_51_n9), .C2(KEY2[51]), .A(KE2_RS_n11), .ZN(
        KE2_RS_SFF_51_n10) );
  INV_X1 KE2_RS_SFF_51_U2 ( .A(RESET), .ZN(KE2_RS_SFF_51_n9) );
  DFF_X1 KE2_RS_SFF_51_Q_reg ( .D(KE2_RS_SFF_51_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[19]), .QN(KE2_RS_SFF_51_n7) );
  OAI21_X1 KE2_RS_SFF_52_U4 ( .B1(KE2_RS_n11), .B2(KE2_RS_SFF_52_n7), .A(
        KE2_RS_SFF_52_n10), .ZN(KE2_RS_SFF_52_n6) );
  OAI221_X1 KE2_RS_SFF_52_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[52]), .C1(
        KE2_RS_SFF_52_n9), .C2(KEY2[52]), .A(KE2_RS_n11), .ZN(
        KE2_RS_SFF_52_n10) );
  INV_X1 KE2_RS_SFF_52_U2 ( .A(RESET), .ZN(KE2_RS_SFF_52_n9) );
  DFF_X1 KE2_RS_SFF_52_Q_reg ( .D(KE2_RS_SFF_52_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[20]), .QN(KE2_RS_SFF_52_n7) );
  OAI21_X1 KE2_RS_SFF_53_U4 ( .B1(KE2_RS_n11), .B2(KE2_RS_SFF_53_n7), .A(
        KE2_RS_SFF_53_n10), .ZN(KE2_RS_SFF_53_n6) );
  OAI221_X1 KE2_RS_SFF_53_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[53]), .C1(
        KE2_RS_SFF_53_n9), .C2(KEY2[53]), .A(KE2_RS_n11), .ZN(
        KE2_RS_SFF_53_n10) );
  INV_X1 KE2_RS_SFF_53_U2 ( .A(RESET), .ZN(KE2_RS_SFF_53_n9) );
  DFF_X1 KE2_RS_SFF_53_Q_reg ( .D(KE2_RS_SFF_53_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[21]), .QN(KE2_RS_SFF_53_n7) );
  OAI21_X1 KE2_RS_SFF_54_U4 ( .B1(KE2_RS_n11), .B2(KE2_RS_SFF_54_n7), .A(
        KE2_RS_SFF_54_n10), .ZN(KE2_RS_SFF_54_n6) );
  OAI221_X1 KE2_RS_SFF_54_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[54]), .C1(
        KE2_RS_SFF_54_n9), .C2(KEY2[54]), .A(KE2_RS_n11), .ZN(
        KE2_RS_SFF_54_n10) );
  INV_X1 KE2_RS_SFF_54_U2 ( .A(RESET), .ZN(KE2_RS_SFF_54_n9) );
  DFF_X1 KE2_RS_SFF_54_Q_reg ( .D(KE2_RS_SFF_54_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[22]), .QN(KE2_RS_SFF_54_n7) );
  OAI21_X1 KE2_RS_SFF_55_U4 ( .B1(KE2_RS_n11), .B2(KE2_RS_SFF_55_n7), .A(
        KE2_RS_SFF_55_n10), .ZN(KE2_RS_SFF_55_n6) );
  OAI221_X1 KE2_RS_SFF_55_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[55]), .C1(
        KE2_RS_SFF_55_n9), .C2(KEY2[55]), .A(KE2_RS_n11), .ZN(
        KE2_RS_SFF_55_n10) );
  INV_X1 KE2_RS_SFF_55_U2 ( .A(RESET), .ZN(KE2_RS_SFF_55_n9) );
  DFF_X1 KE2_RS_SFF_55_Q_reg ( .D(KE2_RS_SFF_55_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[23]), .QN(KE2_RS_SFF_55_n7) );
  OAI21_X1 KE2_RS_SFF_56_U4 ( .B1(KE2_RS_n11), .B2(KE2_RS_SFF_56_n7), .A(
        KE2_RS_SFF_56_n10), .ZN(KE2_RS_SFF_56_n6) );
  OAI221_X1 KE2_RS_SFF_56_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[56]), .C1(
        KE2_RS_SFF_56_n9), .C2(KEY2[56]), .A(KE2_RS_n11), .ZN(
        KE2_RS_SFF_56_n10) );
  INV_X1 KE2_RS_SFF_56_U2 ( .A(RESET), .ZN(KE2_RS_SFF_56_n9) );
  DFF_X1 KE2_RS_SFF_56_Q_reg ( .D(KE2_RS_SFF_56_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[24]), .QN(KE2_RS_SFF_56_n7) );
  OAI21_X1 KE2_RS_SFF_57_U4 ( .B1(KE2_RS_n11), .B2(KE2_RS_SFF_57_n7), .A(
        KE2_RS_SFF_57_n10), .ZN(KE2_RS_SFF_57_n6) );
  OAI221_X1 KE2_RS_SFF_57_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[57]), .C1(
        KE2_RS_SFF_57_n9), .C2(KEY2[57]), .A(KE2_RS_n11), .ZN(
        KE2_RS_SFF_57_n10) );
  INV_X1 KE2_RS_SFF_57_U2 ( .A(RESET), .ZN(KE2_RS_SFF_57_n9) );
  DFF_X1 KE2_RS_SFF_57_Q_reg ( .D(KE2_RS_SFF_57_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[25]), .QN(KE2_RS_SFF_57_n7) );
  OAI21_X1 KE2_RS_SFF_58_U4 ( .B1(KE2_RS_n8), .B2(KE2_RS_SFF_58_n7), .A(
        KE2_RS_SFF_58_n10), .ZN(KE2_RS_SFF_58_n6) );
  OAI221_X1 KE2_RS_SFF_58_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[58]), .C1(
        KE2_RS_SFF_58_n9), .C2(KEY2[58]), .A(KE2_RS_n8), .ZN(KE2_RS_SFF_58_n10) );
  INV_X1 KE2_RS_SFF_58_U2 ( .A(RESET), .ZN(KE2_RS_SFF_58_n9) );
  DFF_X1 KE2_RS_SFF_58_Q_reg ( .D(KE2_RS_SFF_58_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[26]), .QN(KE2_RS_SFF_58_n7) );
  OAI21_X1 KE2_RS_SFF_59_U4 ( .B1(KE2_RS_n7), .B2(KE2_RS_SFF_59_n7), .A(
        KE2_RS_SFF_59_n10), .ZN(KE2_RS_SFF_59_n6) );
  OAI221_X1 KE2_RS_SFF_59_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[59]), .C1(
        KE2_RS_SFF_59_n9), .C2(KEY2[59]), .A(KE2_RS_n7), .ZN(KE2_RS_SFF_59_n10) );
  INV_X1 KE2_RS_SFF_59_U2 ( .A(RESET), .ZN(KE2_RS_SFF_59_n9) );
  DFF_X1 KE2_RS_SFF_59_Q_reg ( .D(KE2_RS_SFF_59_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[27]), .QN(KE2_RS_SFF_59_n7) );
  OAI21_X1 KE2_RS_SFF_60_U4 ( .B1(KE2_RS_n6), .B2(KE2_RS_SFF_60_n7), .A(
        KE2_RS_SFF_60_n10), .ZN(KE2_RS_SFF_60_n6) );
  OAI221_X1 KE2_RS_SFF_60_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[60]), .C1(
        KE2_RS_SFF_60_n9), .C2(KEY2[60]), .A(KE2_RS_n6), .ZN(KE2_RS_SFF_60_n10) );
  INV_X1 KE2_RS_SFF_60_U2 ( .A(RESET), .ZN(KE2_RS_SFF_60_n9) );
  DFF_X1 KE2_RS_SFF_60_Q_reg ( .D(KE2_RS_SFF_60_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[28]), .QN(KE2_RS_SFF_60_n7) );
  OAI21_X1 KE2_RS_SFF_61_U4 ( .B1(KE2_RS_n11), .B2(KE2_RS_SFF_61_n7), .A(
        KE2_RS_SFF_61_n10), .ZN(KE2_RS_SFF_61_n6) );
  OAI221_X1 KE2_RS_SFF_61_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[61]), .C1(
        KE2_RS_SFF_61_n9), .C2(KEY2[61]), .A(KE2_RS_n11), .ZN(
        KE2_RS_SFF_61_n10) );
  INV_X1 KE2_RS_SFF_61_U2 ( .A(RESET), .ZN(KE2_RS_SFF_61_n9) );
  DFF_X1 KE2_RS_SFF_61_Q_reg ( .D(KE2_RS_SFF_61_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[29]), .QN(KE2_RS_SFF_61_n7) );
  OAI21_X1 KE2_RS_SFF_62_U4 ( .B1(KE2_RS_n10), .B2(KE2_RS_SFF_62_n7), .A(
        KE2_RS_SFF_62_n10), .ZN(KE2_RS_SFF_62_n6) );
  OAI221_X1 KE2_RS_SFF_62_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[62]), .C1(
        KE2_RS_SFF_62_n9), .C2(KEY2[62]), .A(KE2_RS_n10), .ZN(
        KE2_RS_SFF_62_n10) );
  INV_X1 KE2_RS_SFF_62_U2 ( .A(RESET), .ZN(KE2_RS_SFF_62_n9) );
  DFF_X1 KE2_RS_SFF_62_Q_reg ( .D(KE2_RS_SFF_62_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[30]), .QN(KE2_RS_SFF_62_n7) );
  OAI21_X1 KE2_RS_SFF_63_U4 ( .B1(KE2_RS_n9), .B2(KE2_RS_SFF_63_n7), .A(
        KE2_RS_SFF_63_n10), .ZN(KE2_RS_SFF_63_n6) );
  OAI221_X1 KE2_RS_SFF_63_U3 ( .B1(RESET), .B2(KE2_KEY_PERM[63]), .C1(
        KE2_RS_SFF_63_n9), .C2(KEY2[63]), .A(KE2_RS_n9), .ZN(KE2_RS_SFF_63_n10) );
  INV_X1 KE2_RS_SFF_63_U2 ( .A(RESET), .ZN(KE2_RS_SFF_63_n9) );
  DFF_X1 KE2_RS_SFF_63_Q_reg ( .D(KE2_RS_SFF_63_n6), .CK(CLK), .Q(
        KE2_KEY_PERM[31]), .QN(KE2_RS_SFF_63_n7) );
  BUF_X1 KE3_RS_U6 ( .A(KEY_EN), .Z(KE3_RS_n11) );
  BUF_X1 KE3_RS_U5 ( .A(KEY_EN), .Z(KE3_RS_n12) );
  BUF_X1 KE3_RS_U4 ( .A(KEY_EN), .Z(KE3_RS_n10) );
  BUF_X1 KE3_RS_U3 ( .A(KEY_EN), .Z(KE3_RS_n8) );
  BUF_X1 KE3_RS_U2 ( .A(KEY_EN), .Z(KE3_RS_n7) );
  BUF_X1 KE3_RS_U1 ( .A(KEY_EN), .Z(KE3_RS_n9) );
  OAI21_X1 KE3_RS_SFF_0_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_0_n8), .A(
        KE3_RS_SFF_0_n11), .ZN(KE3_RS_SFF_0_n7) );
  OAI221_X1 KE3_RS_SFF_0_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[0]), .C1(
        KE3_RS_SFF_0_n10), .C2(KEY3[0]), .A(KE3_RS_n9), .ZN(KE3_RS_SFF_0_n11)
         );
  INV_X1 KE3_RS_SFF_0_U2 ( .A(RESET), .ZN(KE3_RS_SFF_0_n10) );
  DFF_X1 KE3_RS_SFF_0_Q_reg ( .D(KE3_RS_SFF_0_n7), .CK(CLK), .Q(
        KE3_KEY_PERM[56]), .QN(KE3_RS_SFF_0_n8) );
  OAI21_X1 KE3_RS_SFF_1_U4 ( .B1(KE3_RS_n11), .B2(KE3_RS_SFF_1_n8), .A(
        KE3_RS_SFF_1_n11), .ZN(KE3_RS_SFF_1_n7) );
  OAI221_X1 KE3_RS_SFF_1_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[1]), .C1(
        KE3_RS_SFF_1_n10), .C2(KEY3[1]), .A(KE3_RS_n11), .ZN(KE3_RS_SFF_1_n11)
         );
  INV_X1 KE3_RS_SFF_1_U2 ( .A(RESET), .ZN(KE3_RS_SFF_1_n10) );
  DFF_X1 KE3_RS_SFF_1_Q_reg ( .D(KE3_RS_SFF_1_n7), .CK(CLK), .Q(
        KE3_KEY_PERM[57]), .QN(KE3_RS_SFF_1_n8) );
  OAI21_X1 KE3_RS_SFF_2_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_2_n7), .A(
        KE3_RS_SFF_2_n10), .ZN(KE3_RS_SFF_2_n6) );
  OAI221_X1 KE3_RS_SFF_2_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[2]), .C1(
        KE3_RS_SFF_2_n9), .C2(KEY3[2]), .A(KE3_RS_n7), .ZN(KE3_RS_SFF_2_n10)
         );
  INV_X1 KE3_RS_SFF_2_U2 ( .A(RESET), .ZN(KE3_RS_SFF_2_n9) );
  DFF_X1 KE3_RS_SFF_2_Q_reg ( .D(KE3_RS_SFF_2_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[58]), .QN(KE3_RS_SFF_2_n7) );
  OAI21_X1 KE3_RS_SFF_3_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_3_n7), .A(
        KE3_RS_SFF_3_n10), .ZN(KE3_RS_SFF_3_n6) );
  OAI221_X1 KE3_RS_SFF_3_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[3]), .C1(
        KE3_RS_SFF_3_n9), .C2(KEY3[3]), .A(KE3_RS_n7), .ZN(KE3_RS_SFF_3_n10)
         );
  INV_X1 KE3_RS_SFF_3_U2 ( .A(RESET), .ZN(KE3_RS_SFF_3_n9) );
  DFF_X1 KE3_RS_SFF_3_Q_reg ( .D(KE3_RS_SFF_3_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[59]), .QN(KE3_RS_SFF_3_n7) );
  OAI21_X1 KE3_RS_SFF_4_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_4_n7), .A(
        KE3_RS_SFF_4_n10), .ZN(KE3_RS_SFF_4_n6) );
  OAI221_X1 KE3_RS_SFF_4_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[4]), .C1(
        KE3_RS_SFF_4_n9), .C2(KEY3[4]), .A(KE3_RS_n7), .ZN(KE3_RS_SFF_4_n10)
         );
  INV_X1 KE3_RS_SFF_4_U2 ( .A(RESET), .ZN(KE3_RS_SFF_4_n9) );
  DFF_X1 KE3_RS_SFF_4_Q_reg ( .D(KE3_RS_SFF_4_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[40]), .QN(KE3_RS_SFF_4_n7) );
  OAI21_X1 KE3_RS_SFF_5_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_5_n7), .A(
        KE3_RS_SFF_5_n10), .ZN(KE3_RS_SFF_5_n6) );
  OAI221_X1 KE3_RS_SFF_5_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[5]), .C1(
        KE3_RS_SFF_5_n9), .C2(KEY3[5]), .A(KE3_RS_n7), .ZN(KE3_RS_SFF_5_n10)
         );
  INV_X1 KE3_RS_SFF_5_U2 ( .A(RESET), .ZN(KE3_RS_SFF_5_n9) );
  DFF_X1 KE3_RS_SFF_5_Q_reg ( .D(KE3_RS_SFF_5_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[41]), .QN(KE3_RS_SFF_5_n7) );
  OAI21_X1 KE3_RS_SFF_6_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_6_n7), .A(
        KE3_RS_SFF_6_n10), .ZN(KE3_RS_SFF_6_n6) );
  OAI221_X1 KE3_RS_SFF_6_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[6]), .C1(
        KE3_RS_SFF_6_n9), .C2(KEY3[6]), .A(KE3_RS_n7), .ZN(KE3_RS_SFF_6_n10)
         );
  INV_X1 KE3_RS_SFF_6_U2 ( .A(RESET), .ZN(KE3_RS_SFF_6_n9) );
  DFF_X1 KE3_RS_SFF_6_Q_reg ( .D(KE3_RS_SFF_6_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[42]), .QN(KE3_RS_SFF_6_n7) );
  OAI21_X1 KE3_RS_SFF_7_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_7_n7), .A(
        KE3_RS_SFF_7_n10), .ZN(KE3_RS_SFF_7_n6) );
  OAI221_X1 KE3_RS_SFF_7_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[7]), .C1(
        KE3_RS_SFF_7_n9), .C2(KEY3[7]), .A(KE3_RS_n7), .ZN(KE3_RS_SFF_7_n10)
         );
  INV_X1 KE3_RS_SFF_7_U2 ( .A(RESET), .ZN(KE3_RS_SFF_7_n9) );
  DFF_X1 KE3_RS_SFF_7_Q_reg ( .D(KE3_RS_SFF_7_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[43]), .QN(KE3_RS_SFF_7_n7) );
  OAI21_X1 KE3_RS_SFF_8_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_8_n7), .A(
        KE3_RS_SFF_8_n10), .ZN(KE3_RS_SFF_8_n6) );
  OAI221_X1 KE3_RS_SFF_8_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[8]), .C1(
        KE3_RS_SFF_8_n9), .C2(KEY3[8]), .A(KE3_RS_n7), .ZN(KE3_RS_SFF_8_n10)
         );
  INV_X1 KE3_RS_SFF_8_U2 ( .A(RESET), .ZN(KE3_RS_SFF_8_n9) );
  DFF_X1 KE3_RS_SFF_8_Q_reg ( .D(KE3_RS_SFF_8_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[48]), .QN(KE3_RS_SFF_8_n7) );
  OAI21_X1 KE3_RS_SFF_9_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_9_n7), .A(
        KE3_RS_SFF_9_n10), .ZN(KE3_RS_SFF_9_n6) );
  OAI221_X1 KE3_RS_SFF_9_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[9]), .C1(
        KE3_RS_SFF_9_n9), .C2(KEY3[9]), .A(KE3_RS_n7), .ZN(KE3_RS_SFF_9_n10)
         );
  INV_X1 KE3_RS_SFF_9_U2 ( .A(RESET), .ZN(KE3_RS_SFF_9_n9) );
  DFF_X1 KE3_RS_SFF_9_Q_reg ( .D(KE3_RS_SFF_9_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[49]), .QN(KE3_RS_SFF_9_n7) );
  OAI21_X1 KE3_RS_SFF_10_U4 ( .B1(KE3_RS_n8), .B2(KE3_RS_SFF_10_n7), .A(
        KE3_RS_SFF_10_n10), .ZN(KE3_RS_SFF_10_n6) );
  OAI221_X1 KE3_RS_SFF_10_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[10]), .C1(
        KE3_RS_SFF_10_n9), .C2(KEY3[10]), .A(KE3_RS_n8), .ZN(KE3_RS_SFF_10_n10) );
  INV_X1 KE3_RS_SFF_10_U2 ( .A(RESET), .ZN(KE3_RS_SFF_10_n9) );
  DFF_X1 KE3_RS_SFF_10_Q_reg ( .D(KE3_RS_SFF_10_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[50]), .QN(KE3_RS_SFF_10_n7) );
  OAI21_X1 KE3_RS_SFF_11_U4 ( .B1(KE3_RS_n8), .B2(KE3_RS_SFF_11_n7), .A(
        KE3_RS_SFF_11_n10), .ZN(KE3_RS_SFF_11_n6) );
  OAI221_X1 KE3_RS_SFF_11_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[11]), .C1(
        KE3_RS_SFF_11_n9), .C2(KEY3[11]), .A(KE3_RS_n8), .ZN(KE3_RS_SFF_11_n10) );
  INV_X1 KE3_RS_SFF_11_U2 ( .A(RESET), .ZN(KE3_RS_SFF_11_n9) );
  DFF_X1 KE3_RS_SFF_11_Q_reg ( .D(KE3_RS_SFF_11_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[51]), .QN(KE3_RS_SFF_11_n7) );
  OAI21_X1 KE3_RS_SFF_12_U4 ( .B1(KEY_EN), .B2(KE3_RS_SFF_12_n8), .A(
        KE3_RS_SFF_12_n11), .ZN(KE3_RS_SFF_12_n7) );
  OAI221_X1 KE3_RS_SFF_12_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[12]), .C1(
        KE3_RS_SFF_12_n10), .C2(KEY3[12]), .A(KEY_EN), .ZN(KE3_RS_SFF_12_n11)
         );
  INV_X1 KE3_RS_SFF_12_U2 ( .A(RESET), .ZN(KE3_RS_SFF_12_n10) );
  DFF_X1 KE3_RS_SFF_12_Q_reg ( .D(KE3_RS_SFF_12_n7), .CK(CLK), .Q(
        KE3_KEY_PERM[36]), .QN(KE3_RS_SFF_12_n8) );
  OAI21_X1 KE3_RS_SFF_13_U4 ( .B1(KE3_RS_n12), .B2(KE3_RS_SFF_13_n8), .A(
        KE3_RS_SFF_13_n11), .ZN(KE3_RS_SFF_13_n7) );
  OAI221_X1 KE3_RS_SFF_13_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[13]), .C1(
        KE3_RS_SFF_13_n10), .C2(KEY3[13]), .A(KE3_RS_n12), .ZN(
        KE3_RS_SFF_13_n11) );
  INV_X1 KE3_RS_SFF_13_U2 ( .A(RESET), .ZN(KE3_RS_SFF_13_n10) );
  DFF_X1 KE3_RS_SFF_13_Q_reg ( .D(KE3_RS_SFF_13_n7), .CK(CLK), .Q(
        KE3_KEY_PERM[37]), .QN(KE3_RS_SFF_13_n8) );
  OAI21_X1 KE3_RS_SFF_14_U4 ( .B1(KE3_RS_n8), .B2(KE3_RS_SFF_14_n7), .A(
        KE3_RS_SFF_14_n10), .ZN(KE3_RS_SFF_14_n6) );
  OAI221_X1 KE3_RS_SFF_14_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[14]), .C1(
        KE3_RS_SFF_14_n9), .C2(KEY3[14]), .A(KE3_RS_n8), .ZN(KE3_RS_SFF_14_n10) );
  INV_X1 KE3_RS_SFF_14_U2 ( .A(RESET), .ZN(KE3_RS_SFF_14_n9) );
  DFF_X1 KE3_RS_SFF_14_Q_reg ( .D(KE3_RS_SFF_14_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[38]), .QN(KE3_RS_SFF_14_n7) );
  OAI21_X1 KE3_RS_SFF_15_U4 ( .B1(KE3_RS_n8), .B2(KE3_RS_SFF_15_n7), .A(
        KE3_RS_SFF_15_n10), .ZN(KE3_RS_SFF_15_n6) );
  OAI221_X1 KE3_RS_SFF_15_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[15]), .C1(
        KE3_RS_SFF_15_n9), .C2(KEY3[15]), .A(KE3_RS_n8), .ZN(KE3_RS_SFF_15_n10) );
  INV_X1 KE3_RS_SFF_15_U2 ( .A(RESET), .ZN(KE3_RS_SFF_15_n9) );
  DFF_X1 KE3_RS_SFF_15_Q_reg ( .D(KE3_RS_SFF_15_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[39]), .QN(KE3_RS_SFF_15_n7) );
  OAI21_X1 KE3_RS_SFF_16_U4 ( .B1(KE3_RS_n8), .B2(KE3_RS_SFF_16_n7), .A(
        KE3_RS_SFF_16_n10), .ZN(KE3_RS_SFF_16_n6) );
  OAI221_X1 KE3_RS_SFF_16_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[16]), .C1(
        KE3_RS_SFF_16_n9), .C2(KEY3[16]), .A(KE3_RS_n8), .ZN(KE3_RS_SFF_16_n10) );
  INV_X1 KE3_RS_SFF_16_U2 ( .A(RESET), .ZN(KE3_RS_SFF_16_n9) );
  DFF_X1 KE3_RS_SFF_16_Q_reg ( .D(KE3_RS_SFF_16_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[32]), .QN(KE3_RS_SFF_16_n7) );
  OAI21_X1 KE3_RS_SFF_17_U4 ( .B1(KE3_RS_n8), .B2(KE3_RS_SFF_17_n7), .A(
        KE3_RS_SFF_17_n10), .ZN(KE3_RS_SFF_17_n6) );
  OAI221_X1 KE3_RS_SFF_17_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[17]), .C1(
        KE3_RS_SFF_17_n9), .C2(KEY3[17]), .A(KE3_RS_n8), .ZN(KE3_RS_SFF_17_n10) );
  INV_X1 KE3_RS_SFF_17_U2 ( .A(RESET), .ZN(KE3_RS_SFF_17_n9) );
  DFF_X1 KE3_RS_SFF_17_Q_reg ( .D(KE3_RS_SFF_17_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[33]), .QN(KE3_RS_SFF_17_n7) );
  OAI21_X1 KE3_RS_SFF_18_U4 ( .B1(KE3_RS_n8), .B2(KE3_RS_SFF_18_n7), .A(
        KE3_RS_SFF_18_n10), .ZN(KE3_RS_SFF_18_n6) );
  OAI221_X1 KE3_RS_SFF_18_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[18]), .C1(
        KE3_RS_SFF_18_n9), .C2(KEY3[18]), .A(KE3_RS_n8), .ZN(KE3_RS_SFF_18_n10) );
  INV_X1 KE3_RS_SFF_18_U2 ( .A(RESET), .ZN(KE3_RS_SFF_18_n9) );
  DFF_X1 KE3_RS_SFF_18_Q_reg ( .D(KE3_RS_SFF_18_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[34]), .QN(KE3_RS_SFF_18_n7) );
  OAI21_X1 KE3_RS_SFF_19_U4 ( .B1(KE3_RS_n8), .B2(KE3_RS_SFF_19_n7), .A(
        KE3_RS_SFF_19_n10), .ZN(KE3_RS_SFF_19_n6) );
  OAI221_X1 KE3_RS_SFF_19_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[19]), .C1(
        KE3_RS_SFF_19_n9), .C2(KEY3[19]), .A(KE3_RS_n8), .ZN(KE3_RS_SFF_19_n10) );
  INV_X1 KE3_RS_SFF_19_U2 ( .A(RESET), .ZN(KE3_RS_SFF_19_n9) );
  DFF_X1 KE3_RS_SFF_19_Q_reg ( .D(KE3_RS_SFF_19_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[35]), .QN(KE3_RS_SFF_19_n7) );
  OAI21_X1 KE3_RS_SFF_20_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_20_n7), .A(
        KE3_RS_SFF_20_n10), .ZN(KE3_RS_SFF_20_n6) );
  OAI221_X1 KE3_RS_SFF_20_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[20]), .C1(
        KE3_RS_SFF_20_n9), .C2(KEY3[20]), .A(KE3_RS_n9), .ZN(KE3_RS_SFF_20_n10) );
  INV_X1 KE3_RS_SFF_20_U2 ( .A(RESET), .ZN(KE3_RS_SFF_20_n9) );
  DFF_X1 KE3_RS_SFF_20_Q_reg ( .D(KE3_RS_SFF_20_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[44]), .QN(KE3_RS_SFF_20_n7) );
  OAI21_X1 KE3_RS_SFF_21_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_21_n7), .A(
        KE3_RS_SFF_21_n10), .ZN(KE3_RS_SFF_21_n6) );
  OAI221_X1 KE3_RS_SFF_21_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[21]), .C1(
        KE3_RS_SFF_21_n9), .C2(KEY3[21]), .A(KE3_RS_n9), .ZN(KE3_RS_SFF_21_n10) );
  INV_X1 KE3_RS_SFF_21_U2 ( .A(RESET), .ZN(KE3_RS_SFF_21_n9) );
  DFF_X1 KE3_RS_SFF_21_Q_reg ( .D(KE3_RS_SFF_21_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[45]), .QN(KE3_RS_SFF_21_n7) );
  OAI21_X1 KE3_RS_SFF_22_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_22_n7), .A(
        KE3_RS_SFF_22_n10), .ZN(KE3_RS_SFF_22_n6) );
  OAI221_X1 KE3_RS_SFF_22_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[22]), .C1(
        KE3_RS_SFF_22_n9), .C2(KEY3[22]), .A(KE3_RS_n9), .ZN(KE3_RS_SFF_22_n10) );
  INV_X1 KE3_RS_SFF_22_U2 ( .A(RESET), .ZN(KE3_RS_SFF_22_n9) );
  DFF_X1 KE3_RS_SFF_22_Q_reg ( .D(KE3_RS_SFF_22_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[46]), .QN(KE3_RS_SFF_22_n7) );
  OAI21_X1 KE3_RS_SFF_23_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_23_n7), .A(
        KE3_RS_SFF_23_n10), .ZN(KE3_RS_SFF_23_n6) );
  OAI221_X1 KE3_RS_SFF_23_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[23]), .C1(
        KE3_RS_SFF_23_n9), .C2(KEY3[23]), .A(KE3_RS_n9), .ZN(KE3_RS_SFF_23_n10) );
  INV_X1 KE3_RS_SFF_23_U2 ( .A(RESET), .ZN(KE3_RS_SFF_23_n9) );
  DFF_X1 KE3_RS_SFF_23_Q_reg ( .D(KE3_RS_SFF_23_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[47]), .QN(KE3_RS_SFF_23_n7) );
  OAI21_X1 KE3_RS_SFF_24_U4 ( .B1(KE3_RS_n10), .B2(KE3_RS_SFF_24_n8), .A(
        KE3_RS_SFF_24_n11), .ZN(KE3_RS_SFF_24_n7) );
  OAI221_X1 KE3_RS_SFF_24_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[24]), .C1(
        KE3_RS_SFF_24_n10), .C2(KEY3[24]), .A(KE3_RS_n10), .ZN(
        KE3_RS_SFF_24_n11) );
  INV_X1 KE3_RS_SFF_24_U2 ( .A(RESET), .ZN(KE3_RS_SFF_24_n10) );
  DFF_X1 KE3_RS_SFF_24_Q_reg ( .D(KE3_RS_SFF_24_n7), .CK(CLK), .Q(
        KE3_KEY_PERM[60]), .QN(KE3_RS_SFF_24_n8) );
  OAI21_X1 KE3_RS_SFF_25_U4 ( .B1(KE3_RS_n8), .B2(KE3_RS_SFF_25_n8), .A(
        KE3_RS_SFF_25_n11), .ZN(KE3_RS_SFF_25_n7) );
  OAI221_X1 KE3_RS_SFF_25_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[25]), .C1(
        KE3_RS_SFF_25_n10), .C2(KEY3[25]), .A(KE3_RS_n8), .ZN(
        KE3_RS_SFF_25_n11) );
  INV_X1 KE3_RS_SFF_25_U2 ( .A(RESET), .ZN(KE3_RS_SFF_25_n10) );
  DFF_X1 KE3_RS_SFF_25_Q_reg ( .D(KE3_RS_SFF_25_n7), .CK(CLK), .Q(
        KE3_KEY_PERM[61]), .QN(KE3_RS_SFF_25_n8) );
  OAI21_X1 KE3_RS_SFF_26_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_26_n7), .A(
        KE3_RS_SFF_26_n10), .ZN(KE3_RS_SFF_26_n6) );
  OAI221_X1 KE3_RS_SFF_26_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[26]), .C1(
        KE3_RS_SFF_26_n9), .C2(KEY3[26]), .A(KE3_RS_n9), .ZN(KE3_RS_SFF_26_n10) );
  INV_X1 KE3_RS_SFF_26_U2 ( .A(RESET), .ZN(KE3_RS_SFF_26_n9) );
  DFF_X1 KE3_RS_SFF_26_Q_reg ( .D(KE3_RS_SFF_26_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[62]), .QN(KE3_RS_SFF_26_n7) );
  OAI21_X1 KE3_RS_SFF_27_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_27_n7), .A(
        KE3_RS_SFF_27_n10), .ZN(KE3_RS_SFF_27_n6) );
  OAI221_X1 KE3_RS_SFF_27_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[27]), .C1(
        KE3_RS_SFF_27_n9), .C2(KEY3[27]), .A(KE3_RS_n9), .ZN(KE3_RS_SFF_27_n10) );
  INV_X1 KE3_RS_SFF_27_U2 ( .A(RESET), .ZN(KE3_RS_SFF_27_n9) );
  DFF_X1 KE3_RS_SFF_27_Q_reg ( .D(KE3_RS_SFF_27_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[63]), .QN(KE3_RS_SFF_27_n7) );
  OAI21_X1 KE3_RS_SFF_28_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_28_n7), .A(
        KE3_RS_SFF_28_n10), .ZN(KE3_RS_SFF_28_n6) );
  OAI221_X1 KE3_RS_SFF_28_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[28]), .C1(
        KE3_RS_SFF_28_n9), .C2(KEY3[28]), .A(KE3_RS_n9), .ZN(KE3_RS_SFF_28_n10) );
  INV_X1 KE3_RS_SFF_28_U2 ( .A(RESET), .ZN(KE3_RS_SFF_28_n9) );
  DFF_X1 KE3_RS_SFF_28_Q_reg ( .D(KE3_RS_SFF_28_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[52]), .QN(KE3_RS_SFF_28_n7) );
  OAI21_X1 KE3_RS_SFF_29_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_29_n7), .A(
        KE3_RS_SFF_29_n10), .ZN(KE3_RS_SFF_29_n6) );
  OAI221_X1 KE3_RS_SFF_29_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[29]), .C1(
        KE3_RS_SFF_29_n9), .C2(KEY3[29]), .A(KE3_RS_n9), .ZN(KE3_RS_SFF_29_n10) );
  INV_X1 KE3_RS_SFF_29_U2 ( .A(RESET), .ZN(KE3_RS_SFF_29_n9) );
  DFF_X1 KE3_RS_SFF_29_Q_reg ( .D(KE3_RS_SFF_29_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[53]), .QN(KE3_RS_SFF_29_n7) );
  OAI21_X1 KE3_RS_SFF_30_U4 ( .B1(KE3_RS_n10), .B2(KE3_RS_SFF_30_n7), .A(
        KE3_RS_SFF_30_n10), .ZN(KE3_RS_SFF_30_n6) );
  OAI221_X1 KE3_RS_SFF_30_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[30]), .C1(
        KE3_RS_SFF_30_n9), .C2(KEY3[30]), .A(KE3_RS_n10), .ZN(
        KE3_RS_SFF_30_n10) );
  INV_X1 KE3_RS_SFF_30_U2 ( .A(RESET), .ZN(KE3_RS_SFF_30_n9) );
  DFF_X1 KE3_RS_SFF_30_Q_reg ( .D(KE3_RS_SFF_30_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[54]), .QN(KE3_RS_SFF_30_n7) );
  OAI21_X1 KE3_RS_SFF_31_U4 ( .B1(KE3_RS_n10), .B2(KE3_RS_SFF_31_n7), .A(
        KE3_RS_SFF_31_n10), .ZN(KE3_RS_SFF_31_n6) );
  OAI221_X1 KE3_RS_SFF_31_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[31]), .C1(
        KE3_RS_SFF_31_n9), .C2(KEY3[31]), .A(KE3_RS_n10), .ZN(
        KE3_RS_SFF_31_n10) );
  INV_X1 KE3_RS_SFF_31_U2 ( .A(RESET), .ZN(KE3_RS_SFF_31_n9) );
  DFF_X1 KE3_RS_SFF_31_Q_reg ( .D(KE3_RS_SFF_31_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[55]), .QN(KE3_RS_SFF_31_n7) );
  OAI21_X1 KE3_RS_SFF_32_U4 ( .B1(KE3_RS_n10), .B2(KE3_RS_SFF_32_n7), .A(
        KE3_RS_SFF_32_n10), .ZN(KE3_RS_SFF_32_n6) );
  OAI221_X1 KE3_RS_SFF_32_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[32]), .C1(
        KE3_RS_SFF_32_n9), .C2(KEY3[32]), .A(KE3_RS_n10), .ZN(
        KE3_RS_SFF_32_n10) );
  INV_X1 KE3_RS_SFF_32_U2 ( .A(RESET), .ZN(KE3_RS_SFF_32_n9) );
  DFF_X1 KE3_RS_SFF_32_Q_reg ( .D(KE3_RS_SFF_32_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[0]), .QN(KE3_RS_SFF_32_n7) );
  OAI21_X1 KE3_RS_SFF_33_U4 ( .B1(KE3_RS_n10), .B2(KE3_RS_SFF_33_n7), .A(
        KE3_RS_SFF_33_n10), .ZN(KE3_RS_SFF_33_n6) );
  OAI221_X1 KE3_RS_SFF_33_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[33]), .C1(
        KE3_RS_SFF_33_n9), .C2(KEY3[33]), .A(KE3_RS_n10), .ZN(
        KE3_RS_SFF_33_n10) );
  INV_X1 KE3_RS_SFF_33_U2 ( .A(RESET), .ZN(KE3_RS_SFF_33_n9) );
  DFF_X1 KE3_RS_SFF_33_Q_reg ( .D(KE3_RS_SFF_33_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[1]), .QN(KE3_RS_SFF_33_n7) );
  OAI21_X1 KE3_RS_SFF_34_U4 ( .B1(KE3_RS_n10), .B2(KE3_RS_SFF_34_n7), .A(
        KE3_RS_SFF_34_n10), .ZN(KE3_RS_SFF_34_n6) );
  OAI221_X1 KE3_RS_SFF_34_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[34]), .C1(
        KE3_RS_SFF_34_n9), .C2(KEY3[34]), .A(KE3_RS_n10), .ZN(
        KE3_RS_SFF_34_n10) );
  INV_X1 KE3_RS_SFF_34_U2 ( .A(RESET), .ZN(KE3_RS_SFF_34_n9) );
  DFF_X1 KE3_RS_SFF_34_Q_reg ( .D(KE3_RS_SFF_34_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[2]), .QN(KE3_RS_SFF_34_n7) );
  OAI21_X1 KE3_RS_SFF_35_U4 ( .B1(KE3_RS_n10), .B2(KE3_RS_SFF_35_n7), .A(
        KE3_RS_SFF_35_n10), .ZN(KE3_RS_SFF_35_n6) );
  OAI221_X1 KE3_RS_SFF_35_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[35]), .C1(
        KE3_RS_SFF_35_n9), .C2(KEY3[35]), .A(KE3_RS_n10), .ZN(
        KE3_RS_SFF_35_n10) );
  INV_X1 KE3_RS_SFF_35_U2 ( .A(RESET), .ZN(KE3_RS_SFF_35_n9) );
  DFF_X1 KE3_RS_SFF_35_Q_reg ( .D(KE3_RS_SFF_35_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[3]), .QN(KE3_RS_SFF_35_n7) );
  OAI21_X1 KE3_RS_SFF_36_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_36_n8), .A(
        KE3_RS_SFF_36_n11), .ZN(KE3_RS_SFF_36_n7) );
  OAI221_X1 KE3_RS_SFF_36_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[36]), .C1(
        KE3_RS_SFF_36_n10), .C2(KEY3[36]), .A(KE3_RS_n7), .ZN(
        KE3_RS_SFF_36_n11) );
  INV_X1 KE3_RS_SFF_36_U2 ( .A(RESET), .ZN(KE3_RS_SFF_36_n10) );
  DFF_X1 KE3_RS_SFF_36_Q_reg ( .D(KE3_RS_SFF_36_n7), .CK(CLK), .Q(
        KE3_KEY_PERM[4]), .QN(KE3_RS_SFF_36_n8) );
  OAI21_X1 KE3_RS_SFF_37_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_37_n8), .A(
        KE3_RS_SFF_37_n11), .ZN(KE3_RS_SFF_37_n7) );
  OAI221_X1 KE3_RS_SFF_37_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[37]), .C1(
        KE3_RS_SFF_37_n10), .C2(KEY3[37]), .A(KE3_RS_n9), .ZN(
        KE3_RS_SFF_37_n11) );
  INV_X1 KE3_RS_SFF_37_U2 ( .A(RESET), .ZN(KE3_RS_SFF_37_n10) );
  DFF_X1 KE3_RS_SFF_37_Q_reg ( .D(KE3_RS_SFF_37_n7), .CK(CLK), .Q(
        KE3_KEY_PERM[5]), .QN(KE3_RS_SFF_37_n8) );
  OAI21_X1 KE3_RS_SFF_38_U4 ( .B1(KE3_RS_n10), .B2(KE3_RS_SFF_38_n7), .A(
        KE3_RS_SFF_38_n10), .ZN(KE3_RS_SFF_38_n6) );
  OAI221_X1 KE3_RS_SFF_38_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[38]), .C1(
        KE3_RS_SFF_38_n9), .C2(KEY3[38]), .A(KE3_RS_n10), .ZN(
        KE3_RS_SFF_38_n10) );
  INV_X1 KE3_RS_SFF_38_U2 ( .A(RESET), .ZN(KE3_RS_SFF_38_n9) );
  DFF_X1 KE3_RS_SFF_38_Q_reg ( .D(KE3_RS_SFF_38_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[6]), .QN(KE3_RS_SFF_38_n7) );
  OAI21_X1 KE3_RS_SFF_39_U4 ( .B1(KE3_RS_n10), .B2(KE3_RS_SFF_39_n7), .A(
        KE3_RS_SFF_39_n10), .ZN(KE3_RS_SFF_39_n6) );
  OAI221_X1 KE3_RS_SFF_39_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[39]), .C1(
        KE3_RS_SFF_39_n9), .C2(KEY3[39]), .A(KE3_RS_n10), .ZN(
        KE3_RS_SFF_39_n10) );
  INV_X1 KE3_RS_SFF_39_U2 ( .A(RESET), .ZN(KE3_RS_SFF_39_n9) );
  DFF_X1 KE3_RS_SFF_39_Q_reg ( .D(KE3_RS_SFF_39_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[7]), .QN(KE3_RS_SFF_39_n7) );
  OAI21_X1 KE3_RS_SFF_40_U4 ( .B1(KE3_RS_n11), .B2(KE3_RS_SFF_40_n7), .A(
        KE3_RS_SFF_40_n10), .ZN(KE3_RS_SFF_40_n6) );
  OAI221_X1 KE3_RS_SFF_40_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[40]), .C1(
        KE3_RS_SFF_40_n9), .C2(KEY3[40]), .A(KE3_RS_n11), .ZN(
        KE3_RS_SFF_40_n10) );
  INV_X1 KE3_RS_SFF_40_U2 ( .A(RESET), .ZN(KE3_RS_SFF_40_n9) );
  DFF_X1 KE3_RS_SFF_40_Q_reg ( .D(KE3_RS_SFF_40_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[8]), .QN(KE3_RS_SFF_40_n7) );
  OAI21_X1 KE3_RS_SFF_41_U4 ( .B1(KE3_RS_n11), .B2(KE3_RS_SFF_41_n7), .A(
        KE3_RS_SFF_41_n10), .ZN(KE3_RS_SFF_41_n6) );
  OAI221_X1 KE3_RS_SFF_41_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[41]), .C1(
        KE3_RS_SFF_41_n9), .C2(KEY3[41]), .A(KE3_RS_n11), .ZN(
        KE3_RS_SFF_41_n10) );
  INV_X1 KE3_RS_SFF_41_U2 ( .A(RESET), .ZN(KE3_RS_SFF_41_n9) );
  DFF_X1 KE3_RS_SFF_41_Q_reg ( .D(KE3_RS_SFF_41_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[9]), .QN(KE3_RS_SFF_41_n7) );
  OAI21_X1 KE3_RS_SFF_42_U4 ( .B1(KE3_RS_n11), .B2(KE3_RS_SFF_42_n7), .A(
        KE3_RS_SFF_42_n10), .ZN(KE3_RS_SFF_42_n6) );
  OAI221_X1 KE3_RS_SFF_42_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[42]), .C1(
        KE3_RS_SFF_42_n9), .C2(KEY3[42]), .A(KE3_RS_n11), .ZN(
        KE3_RS_SFF_42_n10) );
  INV_X1 KE3_RS_SFF_42_U2 ( .A(RESET), .ZN(KE3_RS_SFF_42_n9) );
  DFF_X1 KE3_RS_SFF_42_Q_reg ( .D(KE3_RS_SFF_42_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[10]), .QN(KE3_RS_SFF_42_n7) );
  OAI21_X1 KE3_RS_SFF_43_U4 ( .B1(KE3_RS_n11), .B2(KE3_RS_SFF_43_n7), .A(
        KE3_RS_SFF_43_n10), .ZN(KE3_RS_SFF_43_n6) );
  OAI221_X1 KE3_RS_SFF_43_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[43]), .C1(
        KE3_RS_SFF_43_n9), .C2(KEY3[43]), .A(KE3_RS_n11), .ZN(
        KE3_RS_SFF_43_n10) );
  INV_X1 KE3_RS_SFF_43_U2 ( .A(RESET), .ZN(KE3_RS_SFF_43_n9) );
  DFF_X1 KE3_RS_SFF_43_Q_reg ( .D(KE3_RS_SFF_43_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[11]), .QN(KE3_RS_SFF_43_n7) );
  OAI21_X1 KE3_RS_SFF_44_U4 ( .B1(KE3_RS_n11), .B2(KE3_RS_SFF_44_n7), .A(
        KE3_RS_SFF_44_n10), .ZN(KE3_RS_SFF_44_n6) );
  OAI221_X1 KE3_RS_SFF_44_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[44]), .C1(
        KE3_RS_SFF_44_n9), .C2(KEY3[44]), .A(KE3_RS_n11), .ZN(
        KE3_RS_SFF_44_n10) );
  INV_X1 KE3_RS_SFF_44_U2 ( .A(RESET), .ZN(KE3_RS_SFF_44_n9) );
  DFF_X1 KE3_RS_SFF_44_Q_reg ( .D(KE3_RS_SFF_44_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[12]), .QN(KE3_RS_SFF_44_n7) );
  OAI21_X1 KE3_RS_SFF_45_U4 ( .B1(KE3_RS_n11), .B2(KE3_RS_SFF_45_n7), .A(
        KE3_RS_SFF_45_n10), .ZN(KE3_RS_SFF_45_n6) );
  OAI221_X1 KE3_RS_SFF_45_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[45]), .C1(
        KE3_RS_SFF_45_n9), .C2(KEY3[45]), .A(KE3_RS_n11), .ZN(
        KE3_RS_SFF_45_n10) );
  INV_X1 KE3_RS_SFF_45_U2 ( .A(RESET), .ZN(KE3_RS_SFF_45_n9) );
  DFF_X1 KE3_RS_SFF_45_Q_reg ( .D(KE3_RS_SFF_45_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[13]), .QN(KE3_RS_SFF_45_n7) );
  OAI21_X1 KE3_RS_SFF_46_U4 ( .B1(KE3_RS_n11), .B2(KE3_RS_SFF_46_n7), .A(
        KE3_RS_SFF_46_n10), .ZN(KE3_RS_SFF_46_n6) );
  OAI221_X1 KE3_RS_SFF_46_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[46]), .C1(
        KE3_RS_SFF_46_n9), .C2(KEY3[46]), .A(KE3_RS_n11), .ZN(
        KE3_RS_SFF_46_n10) );
  INV_X1 KE3_RS_SFF_46_U2 ( .A(RESET), .ZN(KE3_RS_SFF_46_n9) );
  DFF_X1 KE3_RS_SFF_46_Q_reg ( .D(KE3_RS_SFF_46_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[14]), .QN(KE3_RS_SFF_46_n7) );
  OAI21_X1 KE3_RS_SFF_47_U4 ( .B1(KE3_RS_n11), .B2(KE3_RS_SFF_47_n7), .A(
        KE3_RS_SFF_47_n10), .ZN(KE3_RS_SFF_47_n6) );
  OAI221_X1 KE3_RS_SFF_47_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[47]), .C1(
        KE3_RS_SFF_47_n9), .C2(KEY3[47]), .A(KE3_RS_n11), .ZN(
        KE3_RS_SFF_47_n10) );
  INV_X1 KE3_RS_SFF_47_U2 ( .A(RESET), .ZN(KE3_RS_SFF_47_n9) );
  DFF_X1 KE3_RS_SFF_47_Q_reg ( .D(KE3_RS_SFF_47_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[15]), .QN(KE3_RS_SFF_47_n7) );
  OAI21_X1 KE3_RS_SFF_48_U4 ( .B1(KEY_EN), .B2(KE3_RS_SFF_48_n8), .A(
        KE3_RS_SFF_48_n11), .ZN(KE3_RS_SFF_48_n7) );
  OAI221_X1 KE3_RS_SFF_48_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[48]), .C1(
        KE3_RS_SFF_48_n10), .C2(KEY3[48]), .A(KEY_EN), .ZN(KE3_RS_SFF_48_n11)
         );
  INV_X1 KE3_RS_SFF_48_U2 ( .A(RESET), .ZN(KE3_RS_SFF_48_n10) );
  DFF_X1 KE3_RS_SFF_48_Q_reg ( .D(KE3_RS_SFF_48_n7), .CK(CLK), .Q(
        KE3_KEY_PERM[16]), .QN(KE3_RS_SFF_48_n8) );
  OAI21_X1 KE3_RS_SFF_49_U4 ( .B1(KEY_EN), .B2(KE3_RS_SFF_49_n8), .A(
        KE3_RS_SFF_49_n11), .ZN(KE3_RS_SFF_49_n7) );
  OAI221_X1 KE3_RS_SFF_49_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[49]), .C1(
        KE3_RS_SFF_49_n10), .C2(KEY3[49]), .A(KEY_EN), .ZN(KE3_RS_SFF_49_n11)
         );
  INV_X1 KE3_RS_SFF_49_U2 ( .A(RESET), .ZN(KE3_RS_SFF_49_n10) );
  DFF_X1 KE3_RS_SFF_49_Q_reg ( .D(KE3_RS_SFF_49_n7), .CK(CLK), .Q(
        KE3_KEY_PERM[17]), .QN(KE3_RS_SFF_49_n8) );
  OAI21_X1 KE3_RS_SFF_50_U4 ( .B1(KE3_RS_n12), .B2(KE3_RS_SFF_50_n7), .A(
        KE3_RS_SFF_50_n10), .ZN(KE3_RS_SFF_50_n6) );
  OAI221_X1 KE3_RS_SFF_50_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[50]), .C1(
        KE3_RS_SFF_50_n9), .C2(KEY3[50]), .A(KE3_RS_n12), .ZN(
        KE3_RS_SFF_50_n10) );
  INV_X1 KE3_RS_SFF_50_U2 ( .A(RESET), .ZN(KE3_RS_SFF_50_n9) );
  DFF_X1 KE3_RS_SFF_50_Q_reg ( .D(KE3_RS_SFF_50_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[18]), .QN(KE3_RS_SFF_50_n7) );
  OAI21_X1 KE3_RS_SFF_51_U4 ( .B1(KE3_RS_n12), .B2(KE3_RS_SFF_51_n7), .A(
        KE3_RS_SFF_51_n10), .ZN(KE3_RS_SFF_51_n6) );
  OAI221_X1 KE3_RS_SFF_51_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[51]), .C1(
        KE3_RS_SFF_51_n9), .C2(KEY3[51]), .A(KE3_RS_n12), .ZN(
        KE3_RS_SFF_51_n10) );
  INV_X1 KE3_RS_SFF_51_U2 ( .A(RESET), .ZN(KE3_RS_SFF_51_n9) );
  DFF_X1 KE3_RS_SFF_51_Q_reg ( .D(KE3_RS_SFF_51_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[19]), .QN(KE3_RS_SFF_51_n7) );
  OAI21_X1 KE3_RS_SFF_52_U4 ( .B1(KE3_RS_n12), .B2(KE3_RS_SFF_52_n7), .A(
        KE3_RS_SFF_52_n10), .ZN(KE3_RS_SFF_52_n6) );
  OAI221_X1 KE3_RS_SFF_52_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[52]), .C1(
        KE3_RS_SFF_52_n9), .C2(KEY3[52]), .A(KE3_RS_n12), .ZN(
        KE3_RS_SFF_52_n10) );
  INV_X1 KE3_RS_SFF_52_U2 ( .A(RESET), .ZN(KE3_RS_SFF_52_n9) );
  DFF_X1 KE3_RS_SFF_52_Q_reg ( .D(KE3_RS_SFF_52_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[20]), .QN(KE3_RS_SFF_52_n7) );
  OAI21_X1 KE3_RS_SFF_53_U4 ( .B1(KE3_RS_n12), .B2(KE3_RS_SFF_53_n7), .A(
        KE3_RS_SFF_53_n10), .ZN(KE3_RS_SFF_53_n6) );
  OAI221_X1 KE3_RS_SFF_53_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[53]), .C1(
        KE3_RS_SFF_53_n9), .C2(KEY3[53]), .A(KE3_RS_n12), .ZN(
        KE3_RS_SFF_53_n10) );
  INV_X1 KE3_RS_SFF_53_U2 ( .A(RESET), .ZN(KE3_RS_SFF_53_n9) );
  DFF_X1 KE3_RS_SFF_53_Q_reg ( .D(KE3_RS_SFF_53_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[21]), .QN(KE3_RS_SFF_53_n7) );
  OAI21_X1 KE3_RS_SFF_54_U4 ( .B1(KE3_RS_n12), .B2(KE3_RS_SFF_54_n7), .A(
        KE3_RS_SFF_54_n10), .ZN(KE3_RS_SFF_54_n6) );
  OAI221_X1 KE3_RS_SFF_54_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[54]), .C1(
        KE3_RS_SFF_54_n9), .C2(KEY3[54]), .A(KE3_RS_n12), .ZN(
        KE3_RS_SFF_54_n10) );
  INV_X1 KE3_RS_SFF_54_U2 ( .A(RESET), .ZN(KE3_RS_SFF_54_n9) );
  DFF_X1 KE3_RS_SFF_54_Q_reg ( .D(KE3_RS_SFF_54_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[22]), .QN(KE3_RS_SFF_54_n7) );
  OAI21_X1 KE3_RS_SFF_55_U4 ( .B1(KE3_RS_n12), .B2(KE3_RS_SFF_55_n7), .A(
        KE3_RS_SFF_55_n10), .ZN(KE3_RS_SFF_55_n6) );
  OAI221_X1 KE3_RS_SFF_55_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[55]), .C1(
        KE3_RS_SFF_55_n9), .C2(KEY3[55]), .A(KE3_RS_n12), .ZN(
        KE3_RS_SFF_55_n10) );
  INV_X1 KE3_RS_SFF_55_U2 ( .A(RESET), .ZN(KE3_RS_SFF_55_n9) );
  DFF_X1 KE3_RS_SFF_55_Q_reg ( .D(KE3_RS_SFF_55_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[23]), .QN(KE3_RS_SFF_55_n7) );
  OAI21_X1 KE3_RS_SFF_56_U4 ( .B1(KE3_RS_n12), .B2(KE3_RS_SFF_56_n7), .A(
        KE3_RS_SFF_56_n10), .ZN(KE3_RS_SFF_56_n6) );
  OAI221_X1 KE3_RS_SFF_56_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[56]), .C1(
        KE3_RS_SFF_56_n9), .C2(KEY3[56]), .A(KE3_RS_n12), .ZN(
        KE3_RS_SFF_56_n10) );
  INV_X1 KE3_RS_SFF_56_U2 ( .A(RESET), .ZN(KE3_RS_SFF_56_n9) );
  DFF_X1 KE3_RS_SFF_56_Q_reg ( .D(KE3_RS_SFF_56_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[24]), .QN(KE3_RS_SFF_56_n7) );
  OAI21_X1 KE3_RS_SFF_57_U4 ( .B1(KE3_RS_n12), .B2(KE3_RS_SFF_57_n7), .A(
        KE3_RS_SFF_57_n10), .ZN(KE3_RS_SFF_57_n6) );
  OAI221_X1 KE3_RS_SFF_57_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[57]), .C1(
        KE3_RS_SFF_57_n9), .C2(KEY3[57]), .A(KE3_RS_n12), .ZN(
        KE3_RS_SFF_57_n10) );
  INV_X1 KE3_RS_SFF_57_U2 ( .A(RESET), .ZN(KE3_RS_SFF_57_n9) );
  DFF_X1 KE3_RS_SFF_57_Q_reg ( .D(KE3_RS_SFF_57_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[25]), .QN(KE3_RS_SFF_57_n7) );
  OAI21_X1 KE3_RS_SFF_58_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_58_n7), .A(
        KE3_RS_SFF_58_n10), .ZN(KE3_RS_SFF_58_n6) );
  OAI221_X1 KE3_RS_SFF_58_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[58]), .C1(
        KE3_RS_SFF_58_n9), .C2(KEY3[58]), .A(KE3_RS_n7), .ZN(KE3_RS_SFF_58_n10) );
  INV_X1 KE3_RS_SFF_58_U2 ( .A(RESET), .ZN(KE3_RS_SFF_58_n9) );
  DFF_X1 KE3_RS_SFF_58_Q_reg ( .D(KE3_RS_SFF_58_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[26]), .QN(KE3_RS_SFF_58_n7) );
  OAI21_X1 KE3_RS_SFF_59_U4 ( .B1(KE3_RS_n9), .B2(KE3_RS_SFF_59_n7), .A(
        KE3_RS_SFF_59_n10), .ZN(KE3_RS_SFF_59_n6) );
  OAI221_X1 KE3_RS_SFF_59_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[59]), .C1(
        KE3_RS_SFF_59_n9), .C2(KEY3[59]), .A(KE3_RS_n9), .ZN(KE3_RS_SFF_59_n10) );
  INV_X1 KE3_RS_SFF_59_U2 ( .A(RESET), .ZN(KE3_RS_SFF_59_n9) );
  DFF_X1 KE3_RS_SFF_59_Q_reg ( .D(KE3_RS_SFF_59_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[27]), .QN(KE3_RS_SFF_59_n7) );
  OAI21_X1 KE3_RS_SFF_60_U4 ( .B1(KE3_RS_n12), .B2(KE3_RS_SFF_60_n7), .A(
        KE3_RS_SFF_60_n10), .ZN(KE3_RS_SFF_60_n6) );
  OAI221_X1 KE3_RS_SFF_60_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[60]), .C1(
        KE3_RS_SFF_60_n9), .C2(KEY3[60]), .A(KE3_RS_n12), .ZN(
        KE3_RS_SFF_60_n10) );
  INV_X1 KE3_RS_SFF_60_U2 ( .A(RESET), .ZN(KE3_RS_SFF_60_n9) );
  DFF_X1 KE3_RS_SFF_60_Q_reg ( .D(KE3_RS_SFF_60_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[28]), .QN(KE3_RS_SFF_60_n7) );
  OAI21_X1 KE3_RS_SFF_61_U4 ( .B1(KE3_RS_n10), .B2(KE3_RS_SFF_61_n7), .A(
        KE3_RS_SFF_61_n10), .ZN(KE3_RS_SFF_61_n6) );
  OAI221_X1 KE3_RS_SFF_61_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[61]), .C1(
        KE3_RS_SFF_61_n9), .C2(KEY3[61]), .A(KE3_RS_n10), .ZN(
        KE3_RS_SFF_61_n10) );
  INV_X1 KE3_RS_SFF_61_U2 ( .A(RESET), .ZN(KE3_RS_SFF_61_n9) );
  DFF_X1 KE3_RS_SFF_61_Q_reg ( .D(KE3_RS_SFF_61_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[29]), .QN(KE3_RS_SFF_61_n7) );
  OAI21_X1 KE3_RS_SFF_62_U4 ( .B1(KE3_RS_n8), .B2(KE3_RS_SFF_62_n7), .A(
        KE3_RS_SFF_62_n10), .ZN(KE3_RS_SFF_62_n6) );
  OAI221_X1 KE3_RS_SFF_62_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[62]), .C1(
        KE3_RS_SFF_62_n9), .C2(KEY3[62]), .A(KE3_RS_n8), .ZN(KE3_RS_SFF_62_n10) );
  INV_X1 KE3_RS_SFF_62_U2 ( .A(RESET), .ZN(KE3_RS_SFF_62_n9) );
  DFF_X1 KE3_RS_SFF_62_Q_reg ( .D(KE3_RS_SFF_62_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[30]), .QN(KE3_RS_SFF_62_n7) );
  OAI21_X1 KE3_RS_SFF_63_U4 ( .B1(KE3_RS_n7), .B2(KE3_RS_SFF_63_n7), .A(
        KE3_RS_SFF_63_n10), .ZN(KE3_RS_SFF_63_n6) );
  OAI221_X1 KE3_RS_SFF_63_U3 ( .B1(RESET), .B2(KE3_KEY_PERM[63]), .C1(
        KE3_RS_SFF_63_n9), .C2(KEY3[63]), .A(KE3_RS_n7), .ZN(KE3_RS_SFF_63_n10) );
  INV_X1 KE3_RS_SFF_63_U2 ( .A(RESET), .ZN(KE3_RS_SFF_63_n9) );
  DFF_X1 KE3_RS_SFF_63_Q_reg ( .D(KE3_RS_SFF_63_n6), .CK(CLK), .Q(
        KE3_KEY_PERM[31]), .QN(KE3_RS_SFF_63_n7) );
  NOR2_X1 CL_U19 ( .A1(RESET), .A2(CL_n23), .ZN(CL_n3) );
  NOR2_X1 CL_U18 ( .A1(RESET), .A2(CL_n22), .ZN(CL_n2) );
  AOI221_X1 CL_U17 ( .B1(CL_n9), .B2(CL_n24), .C1(CL_n26), .C2(CL_n11), .A(
        RESET), .ZN(CL_n19) );
  OAI22_X1 CL_U16 ( .A1(CL_n8), .A2(KEY_EN), .B1(CL_n9), .B2(CL_n25), .ZN(
        CL_n18) );
  OAI22_X1 CL_U15 ( .A1(CL_n7), .A2(KEY_EN), .B1(CL_n8), .B2(CL_n25), .ZN(
        CL_n17) );
  OAI22_X1 CL_U14 ( .A1(CL_n6), .A2(KEY_EN), .B1(CL_n7), .B2(CL_n25), .ZN(
        CL_n16) );
  OAI22_X1 CL_U13 ( .A1(CL_n5), .A2(KEY_EN), .B1(CL_n6), .B2(CL_n25), .ZN(
        CL_n15) );
  OAI22_X1 CL_U12 ( .A1(CL_n5), .A2(CL_n25), .B1(CL_n4), .B2(KEY_EN), .ZN(
        CL_n14) );
  NAND2_X1 CL_U11 ( .A1(CL_n13), .A2(KEY_EN), .ZN(CL_n25) );
  NOR2_X1 CL_U10 ( .A1(RESET), .A2(CL_n21), .ZN(CL_n1) );
  INV_X1 CL_U9 ( .A(CL_n26), .ZN(ROUND_CST[0]) );
  XOR2_X1 CL_U8 ( .A(CL_n5), .B(CL_n4), .Z(CL_n26) );
  NOR3_X1 CL_U7 ( .A1(CL_n6), .A2(CL_n7), .A3(CL_n20), .ZN(DONE) );
  NAND4_X1 CL_U6 ( .A1(CL_n4), .A2(CL_n8), .A3(CL_n9), .A4(ROUND_CST[5]), .ZN(
        CL_n20) );
  INV_X1 CL_U5 ( .A(RESET), .ZN(CL_n13) );
  NAND2_X1 CL_U4 ( .A1(CL_n24), .A2(CL_n13), .ZN(CL_N11) );
  BUF_X2 CL_U3 ( .A(CL_N11), .Z(KEY_EN) );
  DFF_X1 CL_SHIFT_reg_1_ ( .D(CL_n1), .CK(CLK), .Q(), .QN(CL_n22) );
  DFF_X1 CL_SHIFT_reg_2_ ( .D(CL_n2), .CK(CLK), .Q(), .QN(CL_n23) );
  DFF_X1 CL_SHIFT_reg_3_ ( .D(CL_n3), .CK(CLK), .Q(CL_n11), .QN(CL_n24) );
  DFF_X1 CL_STATE_reg_5_ ( .D(CL_n14), .CK(CLK), .Q(), .QN(CL_n4) );
  DFF_X1 CL_STATE_reg_4_ ( .D(CL_n15), .CK(CLK), .Q(ROUND_CST[5]), .QN(CL_n5)
         );
  DFF_X1 CL_STATE_reg_3_ ( .D(CL_n16), .CK(CLK), .Q(ROUND_CST[4]), .QN(CL_n6)
         );
  DFF_X1 CL_STATE_reg_2_ ( .D(CL_n17), .CK(CLK), .Q(ROUND_CST[3]), .QN(CL_n7)
         );
  DFF_X1 CL_STATE_reg_1_ ( .D(CL_n18), .CK(CLK), .Q(ROUND_CST[2]), .QN(CL_n8)
         );
  DFF_X1 CL_STATE_reg_0_ ( .D(CL_n19), .CK(CLK), .Q(ROUND_CST[1]), .QN(CL_n9)
         );
  DFF_X1 CL_SHIFT_reg_0_ ( .D(KEY_EN), .CK(CLK), .Q(), .QN(CL_n21) );
endmodule

