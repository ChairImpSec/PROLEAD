module circuit ( sboxIn, randomS2, randomS3, randomS4, randomS5, clk, sboxOut );
  input [23:0] sboxIn;
  input [35:0] randomS2;
  input [17:0] randomS3;
  input [35:0] randomS4;
  input [71:0] randomS5;
  output [23:0] sboxOut;
  input clk;
  wire   s1_linMapOut_0__0_, s1_linMapOut_0__1_, s1_linMapOut_0__3_,
         s1_linMapOut_0__4_, s1_linMapOut_0__5_, s1_linMapOut_0__6_,
         s1_linMapOut_0__7_, s1_linMapOut_1__0_, s1_linMapOut_1__1_,
         s1_linMapOut_1__3_, s1_linMapOut_1__4_, s1_linMapOut_1__5_,
         s1_linMapOut_1__6_, s1_linMapOut_1__7_, s1_linMapOut_2__0_,
         s1_linMapOut_2__1_, s1_linMapOut_2__3_, s1_linMapOut_2__4_,
         s1_linMapOut_2__5_, s1_linMapOut_2__6_, s1_linMapOut_2__7_,
         s1_input_mapping_2_n23, s1_input_mapping_2_n22,
         s1_input_mapping_2_n21, s1_input_mapping_2_n20,
         s1_input_mapping_2_n19, s1_input_mapping_2_n18,
         s1_input_mapping_2_n17, s1_input_mapping_1_n23,
         s1_input_mapping_1_n22, s1_input_mapping_1_n21,
         s1_input_mapping_1_n20, s1_input_mapping_1_n19,
         s1_input_mapping_1_n18, s1_input_mapping_1_n17,
         s1_input_mapping_0_n23, s1_input_mapping_0_n22,
         s1_input_mapping_0_n21, s1_input_mapping_0_n20,
         s1_input_mapping_0_n19, s1_input_mapping_0_n18,
         s1_input_mapping_0_n17, s2_n48, s2_n47, s2_n46, s2_n45, s2_n44,
         s2_n43, s2_n42, s2_n41, s2_n40, s2_n39, s2_n38, s2_n37, s2_n36,
         s2_n35, s2_n34, s2_n33, s2_n32, s2_n31, s2_n30, s2_n29, s2_n28,
         s2_n27, s2_n26, s2_n25, s2_n24, s2_n23, s2_n22, s2_n21, s2_n20,
         s2_n19, s2_n18, s2_n17, s2_n16, s2_n15, s2_n14, s2_n13, s2_n12,
         s2_n11, s2_n10, s2_n9, s2_n8, s2_n7, s2_n6, s2_n5, s2_n4, s2_n3,
         s2_n2, s2_n1, s2_chain_0__1__0_, s2_chain_0__1__1_, s2_chain_0__1__2_,
         s2_chain_0__1__3_, s2_chain_1__1__0_, s2_chain_1__1__1_,
         s2_chain_1__1__2_, s2_chain_1__1__3_, s2_chain_2__1__0_,
         s2_chain_2__1__1_, s2_chain_2__1__2_, s2_chain_2__1__3_,
         s2_regOut_0__1__0_, s2_regOut_0__1__1_, s2_regOut_0__1__2_,
         s2_regOut_0__1__3_, s2_regOut_0__2__0_, s2_regOut_0__2__1_,
         s2_regOut_0__2__2_, s2_regOut_0__2__3_, s2_regOut_0__3__0_,
         s2_regOut_0__3__1_, s2_regOut_0__3__2_, s2_regOut_0__3__3_,
         s2_regOut_1__1__0_, s2_regOut_1__1__1_, s2_regOut_1__1__2_,
         s2_regOut_1__1__3_, s2_regOut_1__2__0_, s2_regOut_1__2__1_,
         s2_regOut_1__2__2_, s2_regOut_1__2__3_, s2_regOut_1__3__0_,
         s2_regOut_1__3__1_, s2_regOut_1__3__2_, s2_regOut_1__3__3_,
         s2_regOut_2__1__0_, s2_regOut_2__1__1_, s2_regOut_2__1__2_,
         s2_regOut_2__1__3_, s2_regOut_2__2__0_, s2_regOut_2__2__1_,
         s2_regOut_2__2__2_, s2_regOut_2__2__3_, s2_regOut_2__3__0_,
         s2_regOut_2__3__1_, s2_regOut_2__3__2_, s2_regOut_2__3__3_,
         s2_gf2_mul_out_0__0__0_, s2_gf2_mul_out_0__0__1_,
         s2_gf2_mul_out_0__0__2_, s2_gf2_mul_out_0__0__3_,
         s2_gf2_mul_out_1__1__0_, s2_gf2_mul_out_1__1__1_,
         s2_gf2_mul_out_1__1__2_, s2_gf2_mul_out_1__1__3_,
         s2_gf2_mul_out_2__2__0_, s2_gf2_mul_out_2__2__1_,
         s2_gf2_mul_out_2__2__2_, s2_gf2_mul_out_2__2__3_, s2_mul1_2_2_n76,
         s2_mul1_2_2_n75, s2_mul1_2_2_n74, s2_mul1_2_2_n73, s2_mul1_2_2_n72,
         s2_mul1_2_2_n71, s2_mul1_2_2_n70, s2_mul1_2_2_n69, s2_mul1_2_2_n68,
         s2_mul1_2_2_n67, s2_mul1_2_2_n66, s2_mul1_2_2_n65, s2_mul1_2_2_n64,
         s2_mul1_2_2_n63, s2_mul1_2_2_n62, s2_mul1_2_2_n61, s2_mul1_2_2_n60,
         s2_mul1_2_2_n59, s2_mul1_2_2_n58, s2_mul1_2_2_n57, s2_mul1_2_2_n56,
         s2_mul1_2_2_n55, s2_mul1_2_2_n54, s2_mul1_2_2_n53, s2_mul1_2_1_n76,
         s2_mul1_2_1_n75, s2_mul1_2_1_n74, s2_mul1_2_1_n73, s2_mul1_2_1_n72,
         s2_mul1_2_1_n71, s2_mul1_2_1_n70, s2_mul1_2_1_n69, s2_mul1_2_1_n68,
         s2_mul1_2_1_n67, s2_mul1_2_1_n66, s2_mul1_2_1_n65, s2_mul1_2_1_n64,
         s2_mul1_2_1_n63, s2_mul1_2_1_n62, s2_mul1_2_1_n61, s2_mul1_2_1_n60,
         s2_mul1_2_1_n59, s2_mul1_2_1_n58, s2_mul1_2_1_n57, s2_mul1_2_1_n56,
         s2_mul1_2_1_n55, s2_mul1_2_1_n54, s2_mul1_2_1_n53, s2_mul1_2_0_n76,
         s2_mul1_2_0_n75, s2_mul1_2_0_n74, s2_mul1_2_0_n73, s2_mul1_2_0_n72,
         s2_mul1_2_0_n71, s2_mul1_2_0_n70, s2_mul1_2_0_n69, s2_mul1_2_0_n68,
         s2_mul1_2_0_n67, s2_mul1_2_0_n66, s2_mul1_2_0_n65, s2_mul1_2_0_n64,
         s2_mul1_2_0_n63, s2_mul1_2_0_n62, s2_mul1_2_0_n61, s2_mul1_2_0_n60,
         s2_mul1_2_0_n59, s2_mul1_2_0_n58, s2_mul1_2_0_n57, s2_mul1_2_0_n56,
         s2_mul1_2_0_n55, s2_mul1_2_0_n54, s2_mul1_2_0_n53, s2_mul1_1_2_n76,
         s2_mul1_1_2_n75, s2_mul1_1_2_n74, s2_mul1_1_2_n73, s2_mul1_1_2_n72,
         s2_mul1_1_2_n71, s2_mul1_1_2_n70, s2_mul1_1_2_n69, s2_mul1_1_2_n68,
         s2_mul1_1_2_n67, s2_mul1_1_2_n66, s2_mul1_1_2_n65, s2_mul1_1_2_n64,
         s2_mul1_1_2_n63, s2_mul1_1_2_n62, s2_mul1_1_2_n61, s2_mul1_1_2_n60,
         s2_mul1_1_2_n59, s2_mul1_1_2_n58, s2_mul1_1_2_n57, s2_mul1_1_2_n56,
         s2_mul1_1_2_n55, s2_mul1_1_2_n54, s2_mul1_1_2_n53, s2_mul1_1_1_n76,
         s2_mul1_1_1_n75, s2_mul1_1_1_n74, s2_mul1_1_1_n73, s2_mul1_1_1_n72,
         s2_mul1_1_1_n71, s2_mul1_1_1_n70, s2_mul1_1_1_n69, s2_mul1_1_1_n68,
         s2_mul1_1_1_n67, s2_mul1_1_1_n66, s2_mul1_1_1_n65, s2_mul1_1_1_n64,
         s2_mul1_1_1_n63, s2_mul1_1_1_n62, s2_mul1_1_1_n61, s2_mul1_1_1_n60,
         s2_mul1_1_1_n59, s2_mul1_1_1_n58, s2_mul1_1_1_n57, s2_mul1_1_1_n56,
         s2_mul1_1_1_n55, s2_mul1_1_1_n54, s2_mul1_1_1_n53, s2_mul1_1_0_n76,
         s2_mul1_1_0_n75, s2_mul1_1_0_n74, s2_mul1_1_0_n73, s2_mul1_1_0_n72,
         s2_mul1_1_0_n71, s2_mul1_1_0_n70, s2_mul1_1_0_n69, s2_mul1_1_0_n68,
         s2_mul1_1_0_n67, s2_mul1_1_0_n66, s2_mul1_1_0_n65, s2_mul1_1_0_n64,
         s2_mul1_1_0_n63, s2_mul1_1_0_n62, s2_mul1_1_0_n61, s2_mul1_1_0_n60,
         s2_mul1_1_0_n59, s2_mul1_1_0_n58, s2_mul1_1_0_n57, s2_mul1_1_0_n56,
         s2_mul1_1_0_n55, s2_mul1_1_0_n54, s2_mul1_1_0_n53, s2_mul1_0_2_n76,
         s2_mul1_0_2_n75, s2_mul1_0_2_n74, s2_mul1_0_2_n73, s2_mul1_0_2_n72,
         s2_mul1_0_2_n71, s2_mul1_0_2_n70, s2_mul1_0_2_n69, s2_mul1_0_2_n68,
         s2_mul1_0_2_n67, s2_mul1_0_2_n66, s2_mul1_0_2_n65, s2_mul1_0_2_n64,
         s2_mul1_0_2_n63, s2_mul1_0_2_n62, s2_mul1_0_2_n61, s2_mul1_0_2_n60,
         s2_mul1_0_2_n59, s2_mul1_0_2_n58, s2_mul1_0_2_n57, s2_mul1_0_2_n56,
         s2_mul1_0_2_n55, s2_mul1_0_2_n54, s2_mul1_0_2_n53, s2_mul1_0_1_n76,
         s2_mul1_0_1_n75, s2_mul1_0_1_n74, s2_mul1_0_1_n73, s2_mul1_0_1_n72,
         s2_mul1_0_1_n71, s2_mul1_0_1_n70, s2_mul1_0_1_n69, s2_mul1_0_1_n68,
         s2_mul1_0_1_n67, s2_mul1_0_1_n66, s2_mul1_0_1_n65, s2_mul1_0_1_n64,
         s2_mul1_0_1_n63, s2_mul1_0_1_n62, s2_mul1_0_1_n61, s2_mul1_0_1_n60,
         s2_mul1_0_1_n59, s2_mul1_0_1_n58, s2_mul1_0_1_n57, s2_mul1_0_1_n56,
         s2_mul1_0_1_n55, s2_mul1_0_1_n54, s2_mul1_0_1_n53, s2_mul1_0_0_n76,
         s2_mul1_0_0_n75, s2_mul1_0_0_n74, s2_mul1_0_0_n73, s2_mul1_0_0_n72,
         s2_mul1_0_0_n71, s2_mul1_0_0_n70, s2_mul1_0_0_n69, s2_mul1_0_0_n68,
         s2_mul1_0_0_n67, s2_mul1_0_0_n66, s2_mul1_0_0_n65, s2_mul1_0_0_n64,
         s2_mul1_0_0_n63, s2_mul1_0_0_n62, s2_mul1_0_0_n61, s2_mul1_0_0_n60,
         s2_mul1_0_0_n59, s2_mul1_0_0_n58, s2_mul1_0_0_n57, s2_mul1_0_0_n56,
         s2_mul1_0_0_n55, s2_mul1_0_0_n54, s2_mul1_0_0_n53, s3_n24, s3_n23,
         s3_n22, s3_n21, s3_n20, s3_n19, s3_n18, s3_n17, s3_n16, s3_n15,
         s3_n14, s3_n13, s3_n12, s3_n11, s3_n10, s3_n9, s3_n8, s3_n7, s3_n6,
         s3_n5, s3_n4, s3_n3, s3_n2, s3_n1, s3_chain_0__1__0_,
         s3_chain_0__1__1_, s3_chain_1__1__0_, s3_chain_1__1__1_,
         s3_chain_2__1__0_, s3_chain_2__1__1_, s3_regOut_0__3__0_,
         s3_regOut_0__3__1_, s3_regOut_0__4__0_, s3_regOut_0__4__1_,
         s3_regOut_0__5__0_, s3_regOut_0__5__1_, s3_regOut_1__3__0_,
         s3_regOut_1__3__1_, s3_regOut_1__4__0_, s3_regOut_1__4__1_,
         s3_regOut_1__5__0_, s3_regOut_1__5__1_, s3_regOut_2__3__0_,
         s3_regOut_2__3__1_, s3_regOut_2__4__0_, s3_regOut_2__4__1_,
         s3_regOut_2__5__0_, s3_regOut_2__5__1_, s3_gf2_mul_out_0__0__0_,
         s3_gf2_mul_out_0__0__1_, s3_gf2_mul_out_1__1__0_,
         s3_gf2_mul_out_1__1__1_, s3_gf2_mul_out_2__2__0_,
         s3_gf2_mul_out_2__2__1_, s3_mul1_2_2_n14, s3_mul1_2_2_n13,
         s3_mul1_2_2_n12, s3_mul1_2_2_n11, s3_mul1_2_1_n14, s3_mul1_2_1_n13,
         s3_mul1_2_1_n12, s3_mul1_2_1_n11, s3_mul1_2_0_n14, s3_mul1_2_0_n13,
         s3_mul1_2_0_n12, s3_mul1_2_0_n11, s3_mul1_1_2_n14, s3_mul1_1_2_n13,
         s3_mul1_1_2_n12, s3_mul1_1_2_n11, s3_mul1_1_1_n14, s3_mul1_1_1_n13,
         s3_mul1_1_1_n12, s3_mul1_1_1_n11, s3_mul1_1_0_n14, s3_mul1_1_0_n13,
         s3_mul1_1_0_n12, s3_mul1_1_0_n11, s3_mul1_0_2_n14, s3_mul1_0_2_n13,
         s3_mul1_0_2_n12, s3_mul1_0_2_n11, s3_mul1_0_1_n14, s3_mul1_0_1_n13,
         s3_mul1_0_1_n12, s3_mul1_0_1_n11, s3_mul1_0_0_n14, s3_mul1_0_0_n13,
         s3_mul1_0_0_n12, s3_mul1_0_0_n11, s4_n36, s4_n35, s4_n34, s4_n33,
         s4_n32, s4_n31, s4_n30, s4_n29, s4_n28, s4_n27, s4_n26, s4_n25,
         s4_n24, s4_n23, s4_n22, s4_n21, s4_n20, s4_n19, s4_n18, s4_n17,
         s4_n16, s4_n15, s4_n14, s4_n13, s4_n12, s4_n11, s4_n10, s4_n9, s4_n8,
         s4_n7, s4_n6, s4_n5, s4_n4, s4_n3, s4_n2, s4_n1, s4_chain_0__1__0_,
         s4_chain_0__1__1_, s4_chain_0__1__2_, s4_chain_0__1__3_,
         s4_chain_1__1__0_, s4_chain_1__1__1_, s4_chain_1__1__2_,
         s4_chain_1__1__3_, s4_chain_2__1__0_, s4_chain_2__1__1_,
         s4_chain_2__1__2_, s4_chain_2__1__3_, s4_regOut_0__1__0_,
         s4_regOut_0__1__1_, s4_regOut_0__1__2_, s4_regOut_0__1__3_,
         s4_regOut_0__2__0_, s4_regOut_0__2__1_, s4_regOut_0__2__2_,
         s4_regOut_0__2__3_, s4_regOut_0__3__0_, s4_regOut_0__3__1_,
         s4_regOut_0__3__2_, s4_regOut_0__3__3_, s4_regOut_1__1__0_,
         s4_regOut_1__1__1_, s4_regOut_1__1__2_, s4_regOut_1__1__3_,
         s4_regOut_1__2__0_, s4_regOut_1__2__1_, s4_regOut_1__2__2_,
         s4_regOut_1__2__3_, s4_regOut_1__3__0_, s4_regOut_1__3__1_,
         s4_regOut_1__3__2_, s4_regOut_1__3__3_, s4_regOut_2__1__0_,
         s4_regOut_2__1__1_, s4_regOut_2__1__2_, s4_regOut_2__1__3_,
         s4_regOut_2__2__0_, s4_regOut_2__2__1_, s4_regOut_2__2__2_,
         s4_regOut_2__2__3_, s4_regOut_2__3__0_, s4_regOut_2__3__1_,
         s4_regOut_2__3__2_, s4_regOut_2__3__3_, s4_inv_out_0__0_,
         s4_inv_out_0__1_, s4_inv_out_1__0_, s4_inv_out_1__1_,
         s4_inv_out_2__0_, s4_inv_out_2__1_, s4_mul1_2_2_n14, s4_mul1_2_2_n13,
         s4_mul1_2_2_n12, s4_mul1_2_2_n11, s4_mul1_2_1_n14, s4_mul1_2_1_n13,
         s4_mul1_2_1_n12, s4_mul1_2_1_n11, s4_mul1_2_0_n14, s4_mul1_2_0_n13,
         s4_mul1_2_0_n12, s4_mul1_2_0_n11, s4_mul1_1_2_n14, s4_mul1_1_2_n13,
         s4_mul1_1_2_n12, s4_mul1_1_2_n11, s4_mul1_1_1_n14, s4_mul1_1_1_n13,
         s4_mul1_1_1_n12, s4_mul1_1_1_n11, s4_mul1_1_0_n14, s4_mul1_1_0_n13,
         s4_mul1_1_0_n12, s4_mul1_1_0_n11, s4_mul1_0_2_n14, s4_mul1_0_2_n13,
         s4_mul1_0_2_n12, s4_mul1_0_2_n11, s4_mul1_0_1_n14, s4_mul1_0_1_n13,
         s4_mul1_0_1_n12, s4_mul1_0_1_n11, s4_mul1_0_0_n14, s4_mul1_0_0_n13,
         s4_mul1_0_0_n12, s4_mul1_0_0_n11, s4_mul2_2_2_n14, s4_mul2_2_2_n13,
         s4_mul2_2_2_n12, s4_mul2_2_2_n11, s4_mul2_2_1_n14, s4_mul2_2_1_n13,
         s4_mul2_2_1_n12, s4_mul2_2_1_n11, s4_mul2_2_0_n14, s4_mul2_2_0_n13,
         s4_mul2_2_0_n12, s4_mul2_2_0_n11, s4_mul2_1_2_n14, s4_mul2_1_2_n13,
         s4_mul2_1_2_n12, s4_mul2_1_2_n11, s4_mul2_1_1_n14, s4_mul2_1_1_n13,
         s4_mul2_1_1_n12, s4_mul2_1_1_n11, s4_mul2_1_0_n14, s4_mul2_1_0_n13,
         s4_mul2_1_0_n12, s4_mul2_1_0_n11, s4_mul2_0_2_n14, s4_mul2_0_2_n13,
         s4_mul2_0_2_n12, s4_mul2_0_2_n11, s4_mul2_0_1_n14, s4_mul2_0_1_n13,
         s4_mul2_0_1_n12, s4_mul2_0_1_n11, s4_mul2_0_0_n14, s4_mul2_0_0_n13,
         s4_mul2_0_0_n12, s4_mul2_0_0_n11, s5_n84, s5_n83, s5_n82, s5_n81,
         s5_n80, s5_n79, s5_n78, s5_n77, s5_n76, s5_n75, s5_n74, s5_n73,
         s5_n72, s5_n71, s5_n70, s5_n69, s5_n68, s5_n67, s5_n66, s5_n65,
         s5_n64, s5_n63, s5_n62, s5_n61, s5_n60, s5_n59, s5_n58, s5_n57,
         s5_n56, s5_n55, s5_n54, s5_n53, s5_n52, s5_n51, s5_n50, s5_n49,
         s5_n48, s5_n47, s5_n46, s5_n45, s5_n44, s5_n43, s5_n42, s5_n41,
         s5_n40, s5_n39, s5_n38, s5_n37, s5_n36, s5_n35, s5_n34, s5_n33,
         s5_n32, s5_n31, s5_n30, s5_n29, s5_n28, s5_n27, s5_n26, s5_n25,
         s5_n24, s5_n23, s5_n22, s5_n21, s5_n20, s5_n19, s5_n18, s5_n17,
         s5_n16, s5_n15, s5_n14, s5_n13, s5_n12, s5_n11, s5_n10, s5_n9, s5_n8,
         s5_n7, s5_n6, s5_n5, s5_n4, s5_n3, s5_n2, s5_n1, s5_chain_0__1__0_,
         s5_chain_0__1__1_, s5_chain_0__1__2_, s5_chain_0__1__3_,
         s5_chain_0__1__4_, s5_chain_0__1__5_, s5_chain_0__1__6_,
         s5_chain_0__1__7_, s5_chain_1__1__0_, s5_chain_1__1__1_,
         s5_chain_1__1__2_, s5_chain_1__1__3_, s5_chain_1__1__4_,
         s5_chain_1__1__5_, s5_chain_1__1__6_, s5_chain_1__1__7_,
         s5_chain_2__1__0_, s5_chain_2__1__1_, s5_chain_2__1__2_,
         s5_chain_2__1__3_, s5_chain_2__1__4_, s5_chain_2__1__5_,
         s5_chain_2__1__6_, s5_chain_2__1__7_, s5_mul1_2_2_n76,
         s5_mul1_2_2_n75, s5_mul1_2_2_n74, s5_mul1_2_2_n73, s5_mul1_2_2_n72,
         s5_mul1_2_2_n71, s5_mul1_2_2_n70, s5_mul1_2_2_n69, s5_mul1_2_2_n68,
         s5_mul1_2_2_n67, s5_mul1_2_2_n66, s5_mul1_2_2_n65, s5_mul1_2_2_n64,
         s5_mul1_2_2_n63, s5_mul1_2_2_n62, s5_mul1_2_2_n61, s5_mul1_2_2_n60,
         s5_mul1_2_2_n59, s5_mul1_2_2_n58, s5_mul1_2_2_n57, s5_mul1_2_2_n56,
         s5_mul1_2_2_n55, s5_mul1_2_2_n54, s5_mul1_2_2_n53, s5_mul1_2_1_n76,
         s5_mul1_2_1_n75, s5_mul1_2_1_n74, s5_mul1_2_1_n73, s5_mul1_2_1_n72,
         s5_mul1_2_1_n71, s5_mul1_2_1_n70, s5_mul1_2_1_n69, s5_mul1_2_1_n68,
         s5_mul1_2_1_n67, s5_mul1_2_1_n66, s5_mul1_2_1_n65, s5_mul1_2_1_n64,
         s5_mul1_2_1_n63, s5_mul1_2_1_n62, s5_mul1_2_1_n61, s5_mul1_2_1_n60,
         s5_mul1_2_1_n59, s5_mul1_2_1_n58, s5_mul1_2_1_n57, s5_mul1_2_1_n56,
         s5_mul1_2_1_n55, s5_mul1_2_1_n54, s5_mul1_2_1_n53, s5_mul1_2_0_n76,
         s5_mul1_2_0_n75, s5_mul1_2_0_n74, s5_mul1_2_0_n73, s5_mul1_2_0_n72,
         s5_mul1_2_0_n71, s5_mul1_2_0_n70, s5_mul1_2_0_n69, s5_mul1_2_0_n68,
         s5_mul1_2_0_n67, s5_mul1_2_0_n66, s5_mul1_2_0_n65, s5_mul1_2_0_n64,
         s5_mul1_2_0_n63, s5_mul1_2_0_n62, s5_mul1_2_0_n61, s5_mul1_2_0_n60,
         s5_mul1_2_0_n59, s5_mul1_2_0_n58, s5_mul1_2_0_n57, s5_mul1_2_0_n56,
         s5_mul1_2_0_n55, s5_mul1_2_0_n54, s5_mul1_2_0_n53, s5_mul1_1_2_n76,
         s5_mul1_1_2_n75, s5_mul1_1_2_n74, s5_mul1_1_2_n73, s5_mul1_1_2_n72,
         s5_mul1_1_2_n71, s5_mul1_1_2_n70, s5_mul1_1_2_n69, s5_mul1_1_2_n68,
         s5_mul1_1_2_n67, s5_mul1_1_2_n66, s5_mul1_1_2_n65, s5_mul1_1_2_n64,
         s5_mul1_1_2_n63, s5_mul1_1_2_n62, s5_mul1_1_2_n61, s5_mul1_1_2_n60,
         s5_mul1_1_2_n59, s5_mul1_1_2_n58, s5_mul1_1_2_n57, s5_mul1_1_2_n56,
         s5_mul1_1_2_n55, s5_mul1_1_2_n54, s5_mul1_1_2_n53, s5_mul1_1_1_n76,
         s5_mul1_1_1_n75, s5_mul1_1_1_n74, s5_mul1_1_1_n73, s5_mul1_1_1_n72,
         s5_mul1_1_1_n71, s5_mul1_1_1_n70, s5_mul1_1_1_n69, s5_mul1_1_1_n68,
         s5_mul1_1_1_n67, s5_mul1_1_1_n66, s5_mul1_1_1_n65, s5_mul1_1_1_n64,
         s5_mul1_1_1_n63, s5_mul1_1_1_n62, s5_mul1_1_1_n61, s5_mul1_1_1_n60,
         s5_mul1_1_1_n59, s5_mul1_1_1_n58, s5_mul1_1_1_n57, s5_mul1_1_1_n56,
         s5_mul1_1_1_n55, s5_mul1_1_1_n54, s5_mul1_1_1_n53, s5_mul1_1_0_n76,
         s5_mul1_1_0_n75, s5_mul1_1_0_n74, s5_mul1_1_0_n73, s5_mul1_1_0_n72,
         s5_mul1_1_0_n71, s5_mul1_1_0_n70, s5_mul1_1_0_n69, s5_mul1_1_0_n68,
         s5_mul1_1_0_n67, s5_mul1_1_0_n66, s5_mul1_1_0_n65, s5_mul1_1_0_n64,
         s5_mul1_1_0_n63, s5_mul1_1_0_n62, s5_mul1_1_0_n61, s5_mul1_1_0_n60,
         s5_mul1_1_0_n59, s5_mul1_1_0_n58, s5_mul1_1_0_n57, s5_mul1_1_0_n56,
         s5_mul1_1_0_n55, s5_mul1_1_0_n54, s5_mul1_1_0_n53, s5_mul1_0_2_n76,
         s5_mul1_0_2_n75, s5_mul1_0_2_n74, s5_mul1_0_2_n73, s5_mul1_0_2_n72,
         s5_mul1_0_2_n71, s5_mul1_0_2_n70, s5_mul1_0_2_n69, s5_mul1_0_2_n68,
         s5_mul1_0_2_n67, s5_mul1_0_2_n66, s5_mul1_0_2_n65, s5_mul1_0_2_n64,
         s5_mul1_0_2_n63, s5_mul1_0_2_n62, s5_mul1_0_2_n61, s5_mul1_0_2_n60,
         s5_mul1_0_2_n59, s5_mul1_0_2_n58, s5_mul1_0_2_n57, s5_mul1_0_2_n56,
         s5_mul1_0_2_n55, s5_mul1_0_2_n54, s5_mul1_0_2_n53, s5_mul1_0_1_n76,
         s5_mul1_0_1_n75, s5_mul1_0_1_n74, s5_mul1_0_1_n73, s5_mul1_0_1_n72,
         s5_mul1_0_1_n71, s5_mul1_0_1_n70, s5_mul1_0_1_n69, s5_mul1_0_1_n68,
         s5_mul1_0_1_n67, s5_mul1_0_1_n66, s5_mul1_0_1_n65, s5_mul1_0_1_n64,
         s5_mul1_0_1_n63, s5_mul1_0_1_n62, s5_mul1_0_1_n61, s5_mul1_0_1_n60,
         s5_mul1_0_1_n59, s5_mul1_0_1_n58, s5_mul1_0_1_n57, s5_mul1_0_1_n56,
         s5_mul1_0_1_n55, s5_mul1_0_1_n54, s5_mul1_0_1_n53, s5_mul1_0_0_n76,
         s5_mul1_0_0_n75, s5_mul1_0_0_n74, s5_mul1_0_0_n73, s5_mul1_0_0_n72,
         s5_mul1_0_0_n71, s5_mul1_0_0_n70, s5_mul1_0_0_n69, s5_mul1_0_0_n68,
         s5_mul1_0_0_n67, s5_mul1_0_0_n66, s5_mul1_0_0_n65, s5_mul1_0_0_n64,
         s5_mul1_0_0_n63, s5_mul1_0_0_n62, s5_mul1_0_0_n61, s5_mul1_0_0_n60,
         s5_mul1_0_0_n59, s5_mul1_0_0_n58, s5_mul1_0_0_n57, s5_mul1_0_0_n56,
         s5_mul1_0_0_n55, s5_mul1_0_0_n54, s5_mul1_0_0_n53, s5_mul2_2_2_n76,
         s5_mul2_2_2_n75, s5_mul2_2_2_n74, s5_mul2_2_2_n73, s5_mul2_2_2_n72,
         s5_mul2_2_2_n71, s5_mul2_2_2_n70, s5_mul2_2_2_n69, s5_mul2_2_2_n68,
         s5_mul2_2_2_n67, s5_mul2_2_2_n66, s5_mul2_2_2_n65, s5_mul2_2_2_n64,
         s5_mul2_2_2_n63, s5_mul2_2_2_n62, s5_mul2_2_2_n61, s5_mul2_2_2_n60,
         s5_mul2_2_2_n59, s5_mul2_2_2_n58, s5_mul2_2_2_n57, s5_mul2_2_2_n56,
         s5_mul2_2_2_n55, s5_mul2_2_2_n54, s5_mul2_2_2_n53, s5_mul2_2_1_n76,
         s5_mul2_2_1_n75, s5_mul2_2_1_n74, s5_mul2_2_1_n73, s5_mul2_2_1_n72,
         s5_mul2_2_1_n71, s5_mul2_2_1_n70, s5_mul2_2_1_n69, s5_mul2_2_1_n68,
         s5_mul2_2_1_n67, s5_mul2_2_1_n66, s5_mul2_2_1_n65, s5_mul2_2_1_n64,
         s5_mul2_2_1_n63, s5_mul2_2_1_n62, s5_mul2_2_1_n61, s5_mul2_2_1_n60,
         s5_mul2_2_1_n59, s5_mul2_2_1_n58, s5_mul2_2_1_n57, s5_mul2_2_1_n56,
         s5_mul2_2_1_n55, s5_mul2_2_1_n54, s5_mul2_2_1_n53, s5_mul2_2_0_n76,
         s5_mul2_2_0_n75, s5_mul2_2_0_n74, s5_mul2_2_0_n73, s5_mul2_2_0_n72,
         s5_mul2_2_0_n71, s5_mul2_2_0_n70, s5_mul2_2_0_n69, s5_mul2_2_0_n68,
         s5_mul2_2_0_n67, s5_mul2_2_0_n66, s5_mul2_2_0_n65, s5_mul2_2_0_n64,
         s5_mul2_2_0_n63, s5_mul2_2_0_n62, s5_mul2_2_0_n61, s5_mul2_2_0_n60,
         s5_mul2_2_0_n59, s5_mul2_2_0_n58, s5_mul2_2_0_n57, s5_mul2_2_0_n56,
         s5_mul2_2_0_n55, s5_mul2_2_0_n54, s5_mul2_2_0_n53, s5_mul2_1_2_n76,
         s5_mul2_1_2_n75, s5_mul2_1_2_n74, s5_mul2_1_2_n73, s5_mul2_1_2_n72,
         s5_mul2_1_2_n71, s5_mul2_1_2_n70, s5_mul2_1_2_n69, s5_mul2_1_2_n68,
         s5_mul2_1_2_n67, s5_mul2_1_2_n66, s5_mul2_1_2_n65, s5_mul2_1_2_n64,
         s5_mul2_1_2_n63, s5_mul2_1_2_n62, s5_mul2_1_2_n61, s5_mul2_1_2_n60,
         s5_mul2_1_2_n59, s5_mul2_1_2_n58, s5_mul2_1_2_n57, s5_mul2_1_2_n56,
         s5_mul2_1_2_n55, s5_mul2_1_2_n54, s5_mul2_1_2_n53, s5_mul2_1_1_n76,
         s5_mul2_1_1_n75, s5_mul2_1_1_n74, s5_mul2_1_1_n73, s5_mul2_1_1_n72,
         s5_mul2_1_1_n71, s5_mul2_1_1_n70, s5_mul2_1_1_n69, s5_mul2_1_1_n68,
         s5_mul2_1_1_n67, s5_mul2_1_1_n66, s5_mul2_1_1_n65, s5_mul2_1_1_n64,
         s5_mul2_1_1_n63, s5_mul2_1_1_n62, s5_mul2_1_1_n61, s5_mul2_1_1_n60,
         s5_mul2_1_1_n59, s5_mul2_1_1_n58, s5_mul2_1_1_n57, s5_mul2_1_1_n56,
         s5_mul2_1_1_n55, s5_mul2_1_1_n54, s5_mul2_1_1_n53, s5_mul2_1_0_n76,
         s5_mul2_1_0_n75, s5_mul2_1_0_n74, s5_mul2_1_0_n73, s5_mul2_1_0_n72,
         s5_mul2_1_0_n71, s5_mul2_1_0_n70, s5_mul2_1_0_n69, s5_mul2_1_0_n68,
         s5_mul2_1_0_n67, s5_mul2_1_0_n66, s5_mul2_1_0_n65, s5_mul2_1_0_n64,
         s5_mul2_1_0_n63, s5_mul2_1_0_n62, s5_mul2_1_0_n61, s5_mul2_1_0_n60,
         s5_mul2_1_0_n59, s5_mul2_1_0_n58, s5_mul2_1_0_n57, s5_mul2_1_0_n56,
         s5_mul2_1_0_n55, s5_mul2_1_0_n54, s5_mul2_1_0_n53, s5_mul2_0_2_n76,
         s5_mul2_0_2_n75, s5_mul2_0_2_n74, s5_mul2_0_2_n73, s5_mul2_0_2_n72,
         s5_mul2_0_2_n71, s5_mul2_0_2_n70, s5_mul2_0_2_n69, s5_mul2_0_2_n68,
         s5_mul2_0_2_n67, s5_mul2_0_2_n66, s5_mul2_0_2_n65, s5_mul2_0_2_n64,
         s5_mul2_0_2_n63, s5_mul2_0_2_n62, s5_mul2_0_2_n61, s5_mul2_0_2_n60,
         s5_mul2_0_2_n59, s5_mul2_0_2_n58, s5_mul2_0_2_n57, s5_mul2_0_2_n56,
         s5_mul2_0_2_n55, s5_mul2_0_2_n54, s5_mul2_0_2_n53, s5_mul2_0_1_n76,
         s5_mul2_0_1_n75, s5_mul2_0_1_n74, s5_mul2_0_1_n73, s5_mul2_0_1_n72,
         s5_mul2_0_1_n71, s5_mul2_0_1_n70, s5_mul2_0_1_n69, s5_mul2_0_1_n68,
         s5_mul2_0_1_n67, s5_mul2_0_1_n66, s5_mul2_0_1_n65, s5_mul2_0_1_n64,
         s5_mul2_0_1_n63, s5_mul2_0_1_n62, s5_mul2_0_1_n61, s5_mul2_0_1_n60,
         s5_mul2_0_1_n59, s5_mul2_0_1_n58, s5_mul2_0_1_n57, s5_mul2_0_1_n56,
         s5_mul2_0_1_n55, s5_mul2_0_1_n54, s5_mul2_0_1_n53, s5_mul2_0_0_n76,
         s5_mul2_0_0_n75, s5_mul2_0_0_n74, s5_mul2_0_0_n73, s5_mul2_0_0_n72,
         s5_mul2_0_0_n71, s5_mul2_0_0_n70, s5_mul2_0_0_n69, s5_mul2_0_0_n68,
         s5_mul2_0_0_n67, s5_mul2_0_0_n66, s5_mul2_0_0_n65, s5_mul2_0_0_n64,
         s5_mul2_0_0_n63, s5_mul2_0_0_n62, s5_mul2_0_0_n61, s5_mul2_0_0_n60,
         s5_mul2_0_0_n59, s5_mul2_0_0_n58, s5_mul2_0_0_n57, s5_mul2_0_0_n56,
         s5_mul2_0_0_n55, s5_mul2_0_0_n54, s5_mul2_0_0_n53, s6_2_n9, s6_2_n8,
         s6_2_n7, s6_1_n9, s6_1_n8, s6_1_n7, s6_0_n9, s6_0_n8, s6_0_n7;
  wire   [23:0] stage1Out;
  wire   [35:0] stage2Out;
  wire   [35:0] stage3Out;
  wire   [35:0] stage4Out;
  wire   [23:0] stage5Out;
  wire   [23:0] stage6Out;
  wire   [23:0] regOut1;
  wire   [35:0] s2_refreshed;
  wire   [23:0] s2_xorResult;
  wire   [11:0] s2_sqsc_out;
  wire   [8:0] s2_sqsc_in;
  wire   [17:0] s3_refreshed;
  wire   [11:0] s3_xorResult;
  wire   [5:0] s3_scale_out;
  wire   [2:0] s3_scale_in;
  wire   [35:0] s4_refreshed;
  wire   [35:0] s4_concat;
  wire   [71:0] s5_regOut;
  wire   [71:0] s5_refreshed;
  wire   [71:0] s5_concat;

  DFF_X1 regOut1_reg_2__7_ ( .D(stage6Out[23]), .CK(clk), .Q(regOut1[23]), 
        .QN() );
  DFF_X1 regOut2_reg_2__7_ ( .D(regOut1[23]), .CK(clk), .Q(sboxOut[23]), .QN()
         );
  DFF_X1 regOut1_reg_2__6_ ( .D(stage6Out[22]), .CK(clk), .Q(regOut1[22]), 
        .QN() );
  DFF_X1 regOut2_reg_2__6_ ( .D(regOut1[22]), .CK(clk), .Q(sboxOut[22]), .QN()
         );
  DFF_X1 regOut1_reg_2__5_ ( .D(stage6Out[21]), .CK(clk), .Q(regOut1[21]), 
        .QN() );
  DFF_X1 regOut2_reg_2__5_ ( .D(regOut1[21]), .CK(clk), .Q(sboxOut[21]), .QN()
         );
  DFF_X1 regOut1_reg_2__4_ ( .D(stage6Out[20]), .CK(clk), .Q(regOut1[20]), 
        .QN() );
  DFF_X1 regOut2_reg_2__4_ ( .D(regOut1[20]), .CK(clk), .Q(sboxOut[20]), .QN()
         );
  DFF_X1 regOut1_reg_2__3_ ( .D(stage6Out[19]), .CK(clk), .Q(regOut1[19]), 
        .QN() );
  DFF_X1 regOut2_reg_2__3_ ( .D(regOut1[19]), .CK(clk), .Q(sboxOut[19]), .QN()
         );
  DFF_X1 regOut1_reg_2__2_ ( .D(stage6Out[18]), .CK(clk), .Q(regOut1[18]), 
        .QN() );
  DFF_X1 regOut2_reg_2__2_ ( .D(regOut1[18]), .CK(clk), .Q(sboxOut[18]), .QN()
         );
  DFF_X1 regOut1_reg_2__1_ ( .D(stage6Out[17]), .CK(clk), .Q(regOut1[17]), 
        .QN() );
  DFF_X1 regOut2_reg_2__1_ ( .D(regOut1[17]), .CK(clk), .Q(sboxOut[17]), .QN()
         );
  DFF_X1 regOut1_reg_2__0_ ( .D(stage6Out[16]), .CK(clk), .Q(regOut1[16]), 
        .QN() );
  DFF_X1 regOut2_reg_2__0_ ( .D(regOut1[16]), .CK(clk), .Q(sboxOut[16]), .QN()
         );
  DFF_X1 regOut1_reg_1__7_ ( .D(stage6Out[15]), .CK(clk), .Q(regOut1[15]), 
        .QN() );
  DFF_X1 regOut2_reg_1__7_ ( .D(regOut1[15]), .CK(clk), .Q(sboxOut[15]), .QN()
         );
  DFF_X1 regOut1_reg_1__6_ ( .D(stage6Out[14]), .CK(clk), .Q(regOut1[14]), 
        .QN() );
  DFF_X1 regOut2_reg_1__6_ ( .D(regOut1[14]), .CK(clk), .Q(sboxOut[14]), .QN()
         );
  DFF_X1 regOut1_reg_1__5_ ( .D(stage6Out[13]), .CK(clk), .Q(regOut1[13]), 
        .QN() );
  DFF_X1 regOut2_reg_1__5_ ( .D(regOut1[13]), .CK(clk), .Q(sboxOut[13]), .QN()
         );
  DFF_X1 regOut1_reg_1__4_ ( .D(stage6Out[12]), .CK(clk), .Q(regOut1[12]), 
        .QN() );
  DFF_X1 regOut2_reg_1__4_ ( .D(regOut1[12]), .CK(clk), .Q(sboxOut[12]), .QN()
         );
  DFF_X1 regOut1_reg_1__3_ ( .D(stage6Out[11]), .CK(clk), .Q(regOut1[11]), 
        .QN() );
  DFF_X1 regOut2_reg_1__3_ ( .D(regOut1[11]), .CK(clk), .Q(sboxOut[11]), .QN()
         );
  DFF_X1 regOut1_reg_1__2_ ( .D(stage6Out[10]), .CK(clk), .Q(regOut1[10]), 
        .QN() );
  DFF_X1 regOut2_reg_1__2_ ( .D(regOut1[10]), .CK(clk), .Q(sboxOut[10]), .QN()
         );
  DFF_X1 regOut1_reg_1__1_ ( .D(stage6Out[9]), .CK(clk), .Q(regOut1[9]), .QN()
         );
  DFF_X1 regOut2_reg_1__1_ ( .D(regOut1[9]), .CK(clk), .Q(sboxOut[9]), .QN()
         );
  DFF_X1 regOut1_reg_1__0_ ( .D(stage6Out[8]), .CK(clk), .Q(regOut1[8]), .QN()
         );
  DFF_X1 regOut2_reg_1__0_ ( .D(regOut1[8]), .CK(clk), .Q(sboxOut[8]), .QN()
         );
  DFF_X1 regOut1_reg_0__7_ ( .D(stage6Out[7]), .CK(clk), .Q(regOut1[7]), .QN()
         );
  DFF_X1 regOut2_reg_0__7_ ( .D(regOut1[7]), .CK(clk), .Q(sboxOut[7]), .QN()
         );
  DFF_X1 regOut1_reg_0__6_ ( .D(stage6Out[6]), .CK(clk), .Q(regOut1[6]), .QN()
         );
  DFF_X1 regOut2_reg_0__6_ ( .D(regOut1[6]), .CK(clk), .Q(), .QN(sboxOut[6])
         );
  DFF_X1 regOut1_reg_0__5_ ( .D(stage6Out[5]), .CK(clk), .Q(regOut1[5]), .QN()
         );
  DFF_X1 regOut2_reg_0__5_ ( .D(regOut1[5]), .CK(clk), .Q(), .QN(sboxOut[5])
         );
  DFF_X1 regOut1_reg_0__4_ ( .D(stage6Out[4]), .CK(clk), .Q(regOut1[4]), .QN()
         );
  DFF_X1 regOut2_reg_0__4_ ( .D(regOut1[4]), .CK(clk), .Q(sboxOut[4]), .QN()
         );
  DFF_X1 regOut1_reg_0__3_ ( .D(stage6Out[3]), .CK(clk), .Q(regOut1[3]), .QN()
         );
  DFF_X1 regOut2_reg_0__3_ ( .D(regOut1[3]), .CK(clk), .Q(sboxOut[3]), .QN()
         );
  DFF_X1 regOut1_reg_0__2_ ( .D(stage6Out[2]), .CK(clk), .Q(regOut1[2]), .QN()
         );
  DFF_X1 regOut2_reg_0__2_ ( .D(regOut1[2]), .CK(clk), .Q(sboxOut[2]), .QN()
         );
  DFF_X1 regOut1_reg_0__1_ ( .D(stage6Out[1]), .CK(clk), .Q(regOut1[1]), .QN()
         );
  DFF_X1 regOut2_reg_0__1_ ( .D(regOut1[1]), .CK(clk), .Q(), .QN(sboxOut[1])
         );
  DFF_X1 regOut1_reg_0__0_ ( .D(stage6Out[0]), .CK(clk), .Q(regOut1[0]), .QN()
         );
  DFF_X1 regOut2_reg_0__0_ ( .D(regOut1[0]), .CK(clk), .Q(), .QN(sboxOut[0])
         );
  DFF_X1 s1_stage1Out_reg_0__0_ ( .D(s1_linMapOut_0__0_), .CK(clk), .Q(
        stage1Out[0]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__1_ ( .D(s1_linMapOut_0__1_), .CK(clk), .Q(
        stage1Out[1]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__2_ ( .D(sboxIn[0]), .CK(clk), .Q(stage1Out[2]), 
        .QN() );
  DFF_X1 s1_stage1Out_reg_0__3_ ( .D(s1_linMapOut_0__3_), .CK(clk), .Q(
        stage1Out[3]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__4_ ( .D(s1_linMapOut_0__4_), .CK(clk), .Q(
        stage1Out[4]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__5_ ( .D(s1_linMapOut_0__5_), .CK(clk), .Q(
        stage1Out[5]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__6_ ( .D(s1_linMapOut_0__6_), .CK(clk), .Q(
        stage1Out[6]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__7_ ( .D(s1_linMapOut_0__7_), .CK(clk), .Q(
        stage1Out[7]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__0_ ( .D(s1_linMapOut_1__0_), .CK(clk), .Q(
        stage1Out[8]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__1_ ( .D(s1_linMapOut_1__1_), .CK(clk), .Q(
        stage1Out[9]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__2_ ( .D(sboxIn[8]), .CK(clk), .Q(stage1Out[10]), 
        .QN() );
  DFF_X1 s1_stage1Out_reg_1__3_ ( .D(s1_linMapOut_1__3_), .CK(clk), .Q(
        stage1Out[11]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__4_ ( .D(s1_linMapOut_1__4_), .CK(clk), .Q(
        stage1Out[12]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__5_ ( .D(s1_linMapOut_1__5_), .CK(clk), .Q(
        stage1Out[13]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__6_ ( .D(s1_linMapOut_1__6_), .CK(clk), .Q(
        stage1Out[14]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__7_ ( .D(s1_linMapOut_1__7_), .CK(clk), .Q(
        stage1Out[15]), .QN() );
  DFF_X1 s1_stage1Out_reg_2__0_ ( .D(s1_linMapOut_2__0_), .CK(clk), .Q(
        stage1Out[16]), .QN() );
  DFF_X1 s1_stage1Out_reg_2__1_ ( .D(s1_linMapOut_2__1_), .CK(clk), .Q(
        stage1Out[17]), .QN() );
  DFF_X1 s1_stage1Out_reg_2__2_ ( .D(sboxIn[16]), .CK(clk), .Q(stage1Out[18]), 
        .QN() );
  DFF_X1 s1_stage1Out_reg_2__3_ ( .D(s1_linMapOut_2__3_), .CK(clk), .Q(
        stage1Out[19]), .QN() );
  DFF_X1 s1_stage1Out_reg_2__4_ ( .D(s1_linMapOut_2__4_), .CK(clk), .Q(
        stage1Out[20]), .QN() );
  DFF_X1 s1_stage1Out_reg_2__5_ ( .D(s1_linMapOut_2__5_), .CK(clk), .Q(
        stage1Out[21]), .QN() );
  DFF_X1 s1_stage1Out_reg_2__6_ ( .D(s1_linMapOut_2__6_), .CK(clk), .Q(
        stage1Out[22]), .QN() );
  DFF_X1 s1_stage1Out_reg_2__7_ ( .D(s1_linMapOut_2__7_), .CK(clk), .Q(
        stage1Out[23]), .QN() );
  XNOR2_X1 s1_input_mapping_2_U14 ( .A(s1_input_mapping_2_n23), .B(
        s1_input_mapping_2_n22), .ZN(s1_linMapOut_2__7_) );
  XOR2_X1 s1_input_mapping_2_U13 ( .A(sboxIn[20]), .B(s1_linMapOut_2__1_), .Z(
        s1_linMapOut_2__6_) );
  XNOR2_X1 s1_input_mapping_2_U12 ( .A(s1_input_mapping_2_n21), .B(
        s1_input_mapping_2_n20), .ZN(s1_linMapOut_2__5_) );
  XNOR2_X1 s1_input_mapping_2_U11 ( .A(sboxIn[16]), .B(s1_input_mapping_2_n22), 
        .ZN(s1_linMapOut_2__4_) );
  XNOR2_X1 s1_input_mapping_2_U10 ( .A(sboxIn[23]), .B(s1_input_mapping_2_n21), 
        .ZN(s1_input_mapping_2_n22) );
  XNOR2_X1 s1_input_mapping_2_U9 ( .A(s1_input_mapping_2_n19), .B(
        s1_input_mapping_2_n18), .ZN(s1_linMapOut_2__3_) );
  XNOR2_X1 s1_input_mapping_2_U8 ( .A(s1_input_mapping_2_n20), .B(sboxIn[19]), 
        .ZN(s1_input_mapping_2_n18) );
  XNOR2_X1 s1_input_mapping_2_U7 ( .A(sboxIn[23]), .B(sboxIn[20]), .ZN(
        s1_input_mapping_2_n19) );
  XOR2_X1 s1_input_mapping_2_U6 ( .A(sboxIn[16]), .B(s1_input_mapping_2_n21), 
        .Z(s1_linMapOut_2__1_) );
  XOR2_X1 s1_input_mapping_2_U5 ( .A(sboxIn[22]), .B(sboxIn[21]), .Z(
        s1_input_mapping_2_n21) );
  XNOR2_X1 s1_input_mapping_2_U4 ( .A(s1_input_mapping_2_n23), .B(
        s1_input_mapping_2_n17), .ZN(s1_linMapOut_2__0_) );
  XNOR2_X1 s1_input_mapping_2_U3 ( .A(sboxIn[22]), .B(sboxIn[19]), .ZN(
        s1_input_mapping_2_n17) );
  XNOR2_X1 s1_input_mapping_2_U2 ( .A(sboxIn[18]), .B(s1_input_mapping_2_n20), 
        .ZN(s1_input_mapping_2_n23) );
  XNOR2_X1 s1_input_mapping_2_U1 ( .A(sboxIn[16]), .B(sboxIn[17]), .ZN(
        s1_input_mapping_2_n20) );
  XNOR2_X1 s1_input_mapping_1_U14 ( .A(s1_input_mapping_1_n23), .B(
        s1_input_mapping_1_n22), .ZN(s1_linMapOut_1__7_) );
  XOR2_X1 s1_input_mapping_1_U13 ( .A(sboxIn[12]), .B(s1_linMapOut_1__1_), .Z(
        s1_linMapOut_1__6_) );
  XNOR2_X1 s1_input_mapping_1_U12 ( .A(s1_input_mapping_1_n21), .B(
        s1_input_mapping_1_n20), .ZN(s1_linMapOut_1__5_) );
  XNOR2_X1 s1_input_mapping_1_U11 ( .A(sboxIn[8]), .B(s1_input_mapping_1_n22), 
        .ZN(s1_linMapOut_1__4_) );
  XNOR2_X1 s1_input_mapping_1_U10 ( .A(sboxIn[15]), .B(s1_input_mapping_1_n21), 
        .ZN(s1_input_mapping_1_n22) );
  XNOR2_X1 s1_input_mapping_1_U9 ( .A(s1_input_mapping_1_n19), .B(
        s1_input_mapping_1_n18), .ZN(s1_linMapOut_1__3_) );
  XNOR2_X1 s1_input_mapping_1_U8 ( .A(s1_input_mapping_1_n20), .B(sboxIn[11]), 
        .ZN(s1_input_mapping_1_n18) );
  XNOR2_X1 s1_input_mapping_1_U7 ( .A(sboxIn[15]), .B(sboxIn[12]), .ZN(
        s1_input_mapping_1_n19) );
  XOR2_X1 s1_input_mapping_1_U6 ( .A(sboxIn[8]), .B(s1_input_mapping_1_n21), 
        .Z(s1_linMapOut_1__1_) );
  XOR2_X1 s1_input_mapping_1_U5 ( .A(sboxIn[14]), .B(sboxIn[13]), .Z(
        s1_input_mapping_1_n21) );
  XNOR2_X1 s1_input_mapping_1_U4 ( .A(s1_input_mapping_1_n23), .B(
        s1_input_mapping_1_n17), .ZN(s1_linMapOut_1__0_) );
  XNOR2_X1 s1_input_mapping_1_U3 ( .A(sboxIn[14]), .B(sboxIn[11]), .ZN(
        s1_input_mapping_1_n17) );
  XNOR2_X1 s1_input_mapping_1_U2 ( .A(sboxIn[10]), .B(s1_input_mapping_1_n20), 
        .ZN(s1_input_mapping_1_n23) );
  XNOR2_X1 s1_input_mapping_1_U1 ( .A(sboxIn[8]), .B(sboxIn[9]), .ZN(
        s1_input_mapping_1_n20) );
  XNOR2_X1 s1_input_mapping_0_U14 ( .A(s1_input_mapping_0_n23), .B(
        s1_input_mapping_0_n22), .ZN(s1_linMapOut_0__7_) );
  XOR2_X1 s1_input_mapping_0_U13 ( .A(sboxIn[4]), .B(s1_linMapOut_0__1_), .Z(
        s1_linMapOut_0__6_) );
  XNOR2_X1 s1_input_mapping_0_U12 ( .A(s1_input_mapping_0_n21), .B(
        s1_input_mapping_0_n20), .ZN(s1_linMapOut_0__5_) );
  XNOR2_X1 s1_input_mapping_0_U11 ( .A(sboxIn[0]), .B(s1_input_mapping_0_n22), 
        .ZN(s1_linMapOut_0__4_) );
  XNOR2_X1 s1_input_mapping_0_U10 ( .A(sboxIn[7]), .B(s1_input_mapping_0_n21), 
        .ZN(s1_input_mapping_0_n22) );
  XNOR2_X1 s1_input_mapping_0_U9 ( .A(s1_input_mapping_0_n19), .B(
        s1_input_mapping_0_n18), .ZN(s1_linMapOut_0__3_) );
  XNOR2_X1 s1_input_mapping_0_U8 ( .A(s1_input_mapping_0_n20), .B(sboxIn[3]), 
        .ZN(s1_input_mapping_0_n18) );
  XNOR2_X1 s1_input_mapping_0_U7 ( .A(sboxIn[7]), .B(sboxIn[4]), .ZN(
        s1_input_mapping_0_n19) );
  XOR2_X1 s1_input_mapping_0_U6 ( .A(sboxIn[0]), .B(s1_input_mapping_0_n21), 
        .Z(s1_linMapOut_0__1_) );
  XOR2_X1 s1_input_mapping_0_U5 ( .A(sboxIn[6]), .B(sboxIn[5]), .Z(
        s1_input_mapping_0_n21) );
  XNOR2_X1 s1_input_mapping_0_U4 ( .A(s1_input_mapping_0_n23), .B(
        s1_input_mapping_0_n17), .ZN(s1_linMapOut_0__0_) );
  XNOR2_X1 s1_input_mapping_0_U3 ( .A(sboxIn[6]), .B(sboxIn[3]), .ZN(
        s1_input_mapping_0_n17) );
  XNOR2_X1 s1_input_mapping_0_U2 ( .A(sboxIn[2]), .B(s1_input_mapping_0_n20), 
        .ZN(s1_input_mapping_0_n23) );
  XNOR2_X1 s1_input_mapping_0_U1 ( .A(sboxIn[0]), .B(sboxIn[1]), .ZN(
        s1_input_mapping_0_n20) );
  XNOR2_X1 s2_U98 ( .A(s2_n48), .B(s2_n47), .ZN(s2_refreshed[33]) );
  XNOR2_X1 s2_U97 ( .A(randomS2[1]), .B(randomS2[5]), .ZN(s2_n47) );
  XOR2_X1 s2_U96 ( .A(s2_gf2_mul_out_2__2__1_), .B(s2_sqsc_out[9]), .Z(s2_n48)
         );
  XNOR2_X1 s2_U95 ( .A(s2_n46), .B(s2_n45), .ZN(s2_refreshed[32]) );
  XNOR2_X1 s2_U94 ( .A(randomS2[0]), .B(randomS2[4]), .ZN(s2_n45) );
  XOR2_X1 s2_U93 ( .A(s2_gf2_mul_out_2__2__0_), .B(s2_sqsc_out[8]), .Z(s2_n46)
         );
  XNOR2_X1 s2_U92 ( .A(s2_n44), .B(s2_xorResult[23]), .ZN(s2_refreshed[31]) );
  XNOR2_X1 s2_U91 ( .A(randomS2[11]), .B(randomS2[7]), .ZN(s2_n44) );
  XNOR2_X1 s2_U90 ( .A(s2_n43), .B(s2_xorResult[22]), .ZN(s2_refreshed[30]) );
  XNOR2_X1 s2_U89 ( .A(randomS2[10]), .B(randomS2[6]), .ZN(s2_n43) );
  XNOR2_X1 s2_U88 ( .A(s2_n42), .B(s2_xorResult[21]), .ZN(s2_refreshed[29]) );
  XNOR2_X1 s2_U87 ( .A(randomS2[9]), .B(randomS2[5]), .ZN(s2_n42) );
  XNOR2_X1 s2_U86 ( .A(s2_n41), .B(s2_xorResult[20]), .ZN(s2_refreshed[28]) );
  XNOR2_X1 s2_U85 ( .A(randomS2[8]), .B(randomS2[4]), .ZN(s2_n41) );
  XNOR2_X1 s2_U84 ( .A(s2_n40), .B(s2_xorResult[19]), .ZN(s2_refreshed[27]) );
  XNOR2_X1 s2_U83 ( .A(randomS2[15]), .B(randomS2[11]), .ZN(s2_n40) );
  XNOR2_X1 s2_U82 ( .A(s2_n39), .B(s2_xorResult[18]), .ZN(s2_refreshed[26]) );
  XNOR2_X1 s2_U81 ( .A(randomS2[14]), .B(randomS2[10]), .ZN(s2_n39) );
  XNOR2_X1 s2_U80 ( .A(s2_n38), .B(s2_xorResult[17]), .ZN(s2_refreshed[25]) );
  XNOR2_X1 s2_U79 ( .A(randomS2[13]), .B(randomS2[9]), .ZN(s2_n38) );
  XNOR2_X1 s2_U78 ( .A(s2_n37), .B(s2_xorResult[16]), .ZN(s2_refreshed[24]) );
  XNOR2_X1 s2_U77 ( .A(randomS2[12]), .B(randomS2[8]), .ZN(s2_n37) );
  XNOR2_X1 s2_U76 ( .A(s2_n36), .B(s2_xorResult[15]), .ZN(s2_refreshed[23]) );
  XNOR2_X1 s2_U75 ( .A(randomS2[19]), .B(randomS2[15]), .ZN(s2_n36) );
  XNOR2_X1 s2_U74 ( .A(s2_n35), .B(s2_xorResult[14]), .ZN(s2_refreshed[22]) );
  XNOR2_X1 s2_U73 ( .A(randomS2[18]), .B(randomS2[14]), .ZN(s2_n35) );
  XNOR2_X1 s2_U72 ( .A(s2_n34), .B(s2_xorResult[13]), .ZN(s2_refreshed[21]) );
  XNOR2_X1 s2_U71 ( .A(randomS2[17]), .B(randomS2[13]), .ZN(s2_n34) );
  XNOR2_X1 s2_U70 ( .A(s2_n33), .B(s2_xorResult[12]), .ZN(s2_refreshed[20]) );
  XNOR2_X1 s2_U69 ( .A(randomS2[16]), .B(randomS2[12]), .ZN(s2_n33) );
  XNOR2_X1 s2_U68 ( .A(s2_n32), .B(s2_n31), .ZN(s2_refreshed[17]) );
  XNOR2_X1 s2_U67 ( .A(randomS2[21]), .B(randomS2[17]), .ZN(s2_n31) );
  XOR2_X1 s2_U66 ( .A(s2_gf2_mul_out_1__1__1_), .B(s2_sqsc_out[5]), .Z(s2_n32)
         );
  XNOR2_X1 s2_U65 ( .A(s2_n30), .B(s2_n29), .ZN(s2_refreshed[16]) );
  XNOR2_X1 s2_U64 ( .A(randomS2[20]), .B(randomS2[16]), .ZN(s2_n29) );
  XOR2_X1 s2_U63 ( .A(s2_gf2_mul_out_1__1__0_), .B(s2_sqsc_out[4]), .Z(s2_n30)
         );
  XNOR2_X1 s2_U62 ( .A(s2_n28), .B(s2_xorResult[11]), .ZN(s2_refreshed[15]) );
  XNOR2_X1 s2_U61 ( .A(randomS2[27]), .B(randomS2[23]), .ZN(s2_n28) );
  XNOR2_X1 s2_U60 ( .A(s2_n27), .B(s2_xorResult[10]), .ZN(s2_refreshed[14]) );
  XNOR2_X1 s2_U59 ( .A(randomS2[26]), .B(randomS2[22]), .ZN(s2_n27) );
  XNOR2_X1 s2_U58 ( .A(s2_n26), .B(s2_xorResult[9]), .ZN(s2_refreshed[13]) );
  XNOR2_X1 s2_U57 ( .A(randomS2[25]), .B(randomS2[21]), .ZN(s2_n26) );
  XNOR2_X1 s2_U56 ( .A(s2_n25), .B(s2_xorResult[8]), .ZN(s2_refreshed[12]) );
  XNOR2_X1 s2_U55 ( .A(randomS2[24]), .B(randomS2[20]), .ZN(s2_n25) );
  XNOR2_X1 s2_U54 ( .A(s2_n24), .B(s2_xorResult[7]), .ZN(s2_refreshed[11]) );
  XNOR2_X1 s2_U53 ( .A(randomS2[31]), .B(randomS2[27]), .ZN(s2_n24) );
  XNOR2_X1 s2_U52 ( .A(s2_n23), .B(s2_xorResult[6]), .ZN(s2_refreshed[10]) );
  XNOR2_X1 s2_U51 ( .A(randomS2[30]), .B(randomS2[26]), .ZN(s2_n23) );
  XNOR2_X1 s2_U50 ( .A(s2_n22), .B(s2_xorResult[5]), .ZN(s2_refreshed[9]) );
  XNOR2_X1 s2_U49 ( .A(randomS2[29]), .B(randomS2[25]), .ZN(s2_n22) );
  XNOR2_X1 s2_U48 ( .A(s2_n21), .B(s2_xorResult[4]), .ZN(s2_refreshed[8]) );
  XNOR2_X1 s2_U47 ( .A(randomS2[28]), .B(randomS2[24]), .ZN(s2_n21) );
  XNOR2_X1 s2_U46 ( .A(s2_n20), .B(s2_xorResult[3]), .ZN(s2_refreshed[7]) );
  XNOR2_X1 s2_U45 ( .A(randomS2[35]), .B(randomS2[31]), .ZN(s2_n20) );
  XNOR2_X1 s2_U44 ( .A(s2_n19), .B(s2_xorResult[2]), .ZN(s2_refreshed[6]) );
  XNOR2_X1 s2_U43 ( .A(randomS2[34]), .B(randomS2[30]), .ZN(s2_n19) );
  XNOR2_X1 s2_U42 ( .A(s2_n18), .B(s2_xorResult[1]), .ZN(s2_refreshed[5]) );
  XNOR2_X1 s2_U41 ( .A(randomS2[33]), .B(randomS2[29]), .ZN(s2_n18) );
  XNOR2_X1 s2_U40 ( .A(s2_n17), .B(s2_xorResult[0]), .ZN(s2_refreshed[4]) );
  XNOR2_X1 s2_U39 ( .A(randomS2[32]), .B(randomS2[28]), .ZN(s2_n17) );
  XNOR2_X1 s2_U38 ( .A(s2_n16), .B(s2_n15), .ZN(s2_refreshed[1]) );
  XNOR2_X1 s2_U37 ( .A(randomS2[1]), .B(randomS2[33]), .ZN(s2_n15) );
  XOR2_X1 s2_U36 ( .A(s2_gf2_mul_out_0__0__1_), .B(s2_sqsc_out[1]), .Z(s2_n16)
         );
  XNOR2_X1 s2_U35 ( .A(s2_n14), .B(s2_n13), .ZN(s2_refreshed[0]) );
  XNOR2_X1 s2_U34 ( .A(randomS2[0]), .B(randomS2[32]), .ZN(s2_n13) );
  XOR2_X1 s2_U33 ( .A(s2_gf2_mul_out_0__0__0_), .B(s2_sqsc_out[0]), .Z(s2_n14)
         );
  XOR2_X1 s2_U32 ( .A(stage1Out[18]), .B(stage1Out[22]), .Z(s2_sqsc_in[7]) );
  XNOR2_X1 s2_U31 ( .A(s2_n11), .B(s2_n12), .ZN(s2_refreshed[35]) );
  XNOR2_X1 s2_U30 ( .A(s2_gf2_mul_out_2__2__3_), .B(s2_sqsc_out[11]), .ZN(
        s2_n12) );
  XOR2_X1 s2_U29 ( .A(randomS2[7]), .B(randomS2[3]), .Z(s2_n11) );
  XOR2_X1 s2_U28 ( .A(stage1Out[10]), .B(stage1Out[14]), .Z(s2_sqsc_in[4]) );
  XNOR2_X1 s2_U27 ( .A(s2_n9), .B(s2_n10), .ZN(s2_refreshed[19]) );
  XNOR2_X1 s2_U26 ( .A(s2_gf2_mul_out_1__1__3_), .B(s2_sqsc_out[7]), .ZN(
        s2_n10) );
  XOR2_X1 s2_U25 ( .A(randomS2[19]), .B(randomS2[23]), .Z(s2_n9) );
  XOR2_X1 s2_U24 ( .A(stage1Out[2]), .B(stage1Out[6]), .Z(s2_sqsc_in[1]) );
  XNOR2_X1 s2_U23 ( .A(s2_n7), .B(s2_n8), .ZN(s2_refreshed[3]) );
  XNOR2_X1 s2_U22 ( .A(s2_gf2_mul_out_0__0__3_), .B(s2_sqsc_out[3]), .ZN(s2_n8) );
  XOR2_X1 s2_U21 ( .A(randomS2[35]), .B(randomS2[3]), .Z(s2_n7) );
  XOR2_X1 s2_U20 ( .A(stage1Out[21]), .B(stage1Out[17]), .Z(s2_sqsc_in[6]) );
  XOR2_X1 s2_U19 ( .A(stage1Out[13]), .B(stage1Out[9]), .Z(s2_sqsc_in[3]) );
  XOR2_X1 s2_U18 ( .A(stage1Out[5]), .B(stage1Out[1]), .Z(s2_sqsc_in[0]) );
  XOR2_X1 s2_U17 ( .A(stage1Out[19]), .B(stage1Out[23]), .Z(s2_sqsc_in[8]) );
  XNOR2_X1 s2_U16 ( .A(s2_n5), .B(s2_n6), .ZN(s2_refreshed[34]) );
  XNOR2_X1 s2_U15 ( .A(s2_gf2_mul_out_2__2__2_), .B(s2_sqsc_out[10]), .ZN(
        s2_n6) );
  XOR2_X1 s2_U14 ( .A(randomS2[6]), .B(randomS2[2]), .Z(s2_n5) );
  XOR2_X1 s2_U13 ( .A(stage1Out[11]), .B(stage1Out[15]), .Z(s2_sqsc_in[5]) );
  XNOR2_X1 s2_U12 ( .A(s2_n3), .B(s2_n4), .ZN(s2_refreshed[18]) );
  XNOR2_X1 s2_U11 ( .A(s2_gf2_mul_out_1__1__2_), .B(s2_sqsc_out[6]), .ZN(s2_n4) );
  XOR2_X1 s2_U10 ( .A(randomS2[18]), .B(randomS2[22]), .Z(s2_n3) );
  XOR2_X1 s2_U9 ( .A(stage1Out[3]), .B(stage1Out[7]), .Z(s2_sqsc_in[2]) );
  XNOR2_X1 s2_U8 ( .A(s2_n1), .B(s2_n2), .ZN(s2_refreshed[2]) );
  XNOR2_X1 s2_U7 ( .A(s2_gf2_mul_out_0__0__2_), .B(s2_sqsc_out[2]), .ZN(s2_n2)
         );
  XOR2_X1 s2_U6 ( .A(randomS2[34]), .B(randomS2[2]), .Z(s2_n1) );
  XOR2_X1 s2_U5 ( .A(stage1Out[20]), .B(stage1Out[16]), .Z(s2_sqsc_out[8]) );
  XOR2_X1 s2_U4 ( .A(stage1Out[12]), .B(stage1Out[8]), .Z(s2_sqsc_out[4]) );
  XOR2_X1 s2_U3 ( .A(stage1Out[4]), .B(stage1Out[0]), .Z(s2_sqsc_out[0]) );
  DFF_X1 s2_regOut_reg_0__0__0_ ( .D(stage1Out[0]), .CK(clk), .Q(stage2Out[0]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__0__1_ ( .D(stage1Out[1]), .CK(clk), .Q(stage2Out[1]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__0__2_ ( .D(stage1Out[2]), .CK(clk), .Q(stage2Out[2]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__0__3_ ( .D(stage1Out[3]), .CK(clk), .Q(stage2Out[3]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__1__0_ ( .D(s2_refreshed[0]), .CK(clk), .Q(
        s2_regOut_0__1__0_), .QN() );
  DFF_X1 s2_regOut_reg_0__1__1_ ( .D(s2_refreshed[1]), .CK(clk), .Q(
        s2_regOut_0__1__1_), .QN() );
  DFF_X1 s2_regOut_reg_0__1__2_ ( .D(s2_refreshed[2]), .CK(clk), .Q(
        s2_regOut_0__1__2_), .QN() );
  DFF_X1 s2_regOut_reg_0__1__3_ ( .D(s2_refreshed[3]), .CK(clk), .Q(
        s2_regOut_0__1__3_), .QN() );
  DFF_X1 s2_regOut_reg_0__2__0_ ( .D(s2_refreshed[4]), .CK(clk), .Q(
        s2_regOut_0__2__0_), .QN() );
  DFF_X1 s2_regOut_reg_0__2__1_ ( .D(s2_refreshed[5]), .CK(clk), .Q(
        s2_regOut_0__2__1_), .QN() );
  DFF_X1 s2_regOut_reg_0__2__2_ ( .D(s2_refreshed[6]), .CK(clk), .Q(
        s2_regOut_0__2__2_), .QN() );
  DFF_X1 s2_regOut_reg_0__2__3_ ( .D(s2_refreshed[7]), .CK(clk), .Q(
        s2_regOut_0__2__3_), .QN() );
  DFF_X1 s2_regOut_reg_0__3__0_ ( .D(s2_refreshed[8]), .CK(clk), .Q(
        s2_regOut_0__3__0_), .QN() );
  DFF_X1 s2_regOut_reg_0__3__1_ ( .D(s2_refreshed[9]), .CK(clk), .Q(
        s2_regOut_0__3__1_), .QN() );
  DFF_X1 s2_regOut_reg_0__3__2_ ( .D(s2_refreshed[10]), .CK(clk), .Q(
        s2_regOut_0__3__2_), .QN() );
  DFF_X1 s2_regOut_reg_0__3__3_ ( .D(s2_refreshed[11]), .CK(clk), .Q(
        s2_regOut_0__3__3_), .QN() );
  DFF_X1 s2_regOut_reg_0__4__0_ ( .D(stage1Out[4]), .CK(clk), .Q(stage2Out[8]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__4__1_ ( .D(stage1Out[5]), .CK(clk), .Q(stage2Out[9]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__4__2_ ( .D(stage1Out[6]), .CK(clk), .Q(stage2Out[10]), .QN() );
  DFF_X1 s2_regOut_reg_0__4__3_ ( .D(stage1Out[7]), .CK(clk), .Q(stage2Out[11]), .QN() );
  DFF_X1 s2_regOut_reg_1__0__0_ ( .D(stage1Out[8]), .CK(clk), .Q(stage2Out[12]), .QN() );
  DFF_X1 s2_regOut_reg_1__0__1_ ( .D(stage1Out[9]), .CK(clk), .Q(stage2Out[13]), .QN() );
  DFF_X1 s2_regOut_reg_1__0__2_ ( .D(stage1Out[10]), .CK(clk), .Q(
        stage2Out[14]), .QN() );
  DFF_X1 s2_regOut_reg_1__0__3_ ( .D(stage1Out[11]), .CK(clk), .Q(
        stage2Out[15]), .QN() );
  DFF_X1 s2_regOut_reg_1__1__0_ ( .D(s2_refreshed[12]), .CK(clk), .Q(
        s2_regOut_1__1__0_), .QN() );
  DFF_X1 s2_regOut_reg_1__1__1_ ( .D(s2_refreshed[13]), .CK(clk), .Q(
        s2_regOut_1__1__1_), .QN() );
  DFF_X1 s2_regOut_reg_1__1__2_ ( .D(s2_refreshed[14]), .CK(clk), .Q(
        s2_regOut_1__1__2_), .QN() );
  DFF_X1 s2_regOut_reg_1__1__3_ ( .D(s2_refreshed[15]), .CK(clk), .Q(
        s2_regOut_1__1__3_), .QN() );
  DFF_X1 s2_regOut_reg_1__2__0_ ( .D(s2_refreshed[16]), .CK(clk), .Q(
        s2_regOut_1__2__0_), .QN() );
  DFF_X1 s2_regOut_reg_1__2__1_ ( .D(s2_refreshed[17]), .CK(clk), .Q(
        s2_regOut_1__2__1_), .QN() );
  DFF_X1 s2_regOut_reg_1__2__2_ ( .D(s2_refreshed[18]), .CK(clk), .Q(
        s2_regOut_1__2__2_), .QN() );
  DFF_X1 s2_regOut_reg_1__2__3_ ( .D(s2_refreshed[19]), .CK(clk), .Q(
        s2_regOut_1__2__3_), .QN() );
  DFF_X1 s2_regOut_reg_1__3__0_ ( .D(s2_refreshed[20]), .CK(clk), .Q(
        s2_regOut_1__3__0_), .QN() );
  DFF_X1 s2_regOut_reg_1__3__1_ ( .D(s2_refreshed[21]), .CK(clk), .Q(
        s2_regOut_1__3__1_), .QN() );
  DFF_X1 s2_regOut_reg_1__3__2_ ( .D(s2_refreshed[22]), .CK(clk), .Q(
        s2_regOut_1__3__2_), .QN() );
  DFF_X1 s2_regOut_reg_1__3__3_ ( .D(s2_refreshed[23]), .CK(clk), .Q(
        s2_regOut_1__3__3_), .QN() );
  DFF_X1 s2_regOut_reg_1__4__0_ ( .D(stage1Out[12]), .CK(clk), .Q(
        stage2Out[20]), .QN() );
  DFF_X1 s2_regOut_reg_1__4__1_ ( .D(stage1Out[13]), .CK(clk), .Q(
        stage2Out[21]), .QN() );
  DFF_X1 s2_regOut_reg_1__4__2_ ( .D(stage1Out[14]), .CK(clk), .Q(
        stage2Out[22]), .QN() );
  DFF_X1 s2_regOut_reg_1__4__3_ ( .D(stage1Out[15]), .CK(clk), .Q(
        stage2Out[23]), .QN() );
  DFF_X1 s2_regOut_reg_2__0__0_ ( .D(stage1Out[16]), .CK(clk), .Q(
        stage2Out[24]), .QN() );
  DFF_X1 s2_regOut_reg_2__0__1_ ( .D(stage1Out[17]), .CK(clk), .Q(
        stage2Out[25]), .QN() );
  DFF_X1 s2_regOut_reg_2__0__2_ ( .D(stage1Out[18]), .CK(clk), .Q(
        stage2Out[26]), .QN() );
  DFF_X1 s2_regOut_reg_2__0__3_ ( .D(stage1Out[19]), .CK(clk), .Q(
        stage2Out[27]), .QN() );
  DFF_X1 s2_regOut_reg_2__1__0_ ( .D(s2_refreshed[24]), .CK(clk), .Q(
        s2_regOut_2__1__0_), .QN() );
  DFF_X1 s2_regOut_reg_2__1__1_ ( .D(s2_refreshed[25]), .CK(clk), .Q(
        s2_regOut_2__1__1_), .QN() );
  DFF_X1 s2_regOut_reg_2__1__2_ ( .D(s2_refreshed[26]), .CK(clk), .Q(
        s2_regOut_2__1__2_), .QN() );
  DFF_X1 s2_regOut_reg_2__1__3_ ( .D(s2_refreshed[27]), .CK(clk), .Q(
        s2_regOut_2__1__3_), .QN() );
  DFF_X1 s2_regOut_reg_2__2__0_ ( .D(s2_refreshed[28]), .CK(clk), .Q(
        s2_regOut_2__2__0_), .QN() );
  DFF_X1 s2_regOut_reg_2__2__1_ ( .D(s2_refreshed[29]), .CK(clk), .Q(
        s2_regOut_2__2__1_), .QN() );
  DFF_X1 s2_regOut_reg_2__2__2_ ( .D(s2_refreshed[30]), .CK(clk), .Q(
        s2_regOut_2__2__2_), .QN() );
  DFF_X1 s2_regOut_reg_2__2__3_ ( .D(s2_refreshed[31]), .CK(clk), .Q(
        s2_regOut_2__2__3_), .QN() );
  DFF_X1 s2_regOut_reg_2__3__0_ ( .D(s2_refreshed[32]), .CK(clk), .Q(
        s2_regOut_2__3__0_), .QN() );
  DFF_X1 s2_regOut_reg_2__3__1_ ( .D(s2_refreshed[33]), .CK(clk), .Q(
        s2_regOut_2__3__1_), .QN() );
  DFF_X1 s2_regOut_reg_2__3__2_ ( .D(s2_refreshed[34]), .CK(clk), .Q(
        s2_regOut_2__3__2_), .QN() );
  DFF_X1 s2_regOut_reg_2__3__3_ ( .D(s2_refreshed[35]), .CK(clk), .Q(
        s2_regOut_2__3__3_), .QN() );
  DFF_X1 s2_regOut_reg_2__4__0_ ( .D(stage1Out[20]), .CK(clk), .Q(
        stage2Out[32]), .QN() );
  DFF_X1 s2_regOut_reg_2__4__1_ ( .D(stage1Out[21]), .CK(clk), .Q(
        stage2Out[33]), .QN() );
  DFF_X1 s2_regOut_reg_2__4__2_ ( .D(stage1Out[22]), .CK(clk), .Q(
        stage2Out[34]), .QN() );
  DFF_X1 s2_regOut_reg_2__4__3_ ( .D(stage1Out[23]), .CK(clk), .Q(
        stage2Out[35]), .QN() );
  XOR2_X1 s2_sqsc_2_U3 ( .A(s2_sqsc_out[8]), .B(s2_sqsc_in[6]), .Z(
        s2_sqsc_out[9]) );
  XOR2_X1 s2_sqsc_2_U2 ( .A(s2_sqsc_out[8]), .B(s2_sqsc_in[7]), .Z(
        s2_sqsc_out[11]) );
  XOR2_X1 s2_sqsc_2_U1 ( .A(s2_sqsc_in[6]), .B(s2_sqsc_in[8]), .Z(
        s2_sqsc_out[10]) );
  XOR2_X1 s2_sqsc_1_U3 ( .A(s2_sqsc_out[4]), .B(s2_sqsc_in[3]), .Z(
        s2_sqsc_out[5]) );
  XOR2_X1 s2_sqsc_1_U2 ( .A(s2_sqsc_out[4]), .B(s2_sqsc_in[4]), .Z(
        s2_sqsc_out[7]) );
  XOR2_X1 s2_sqsc_1_U1 ( .A(s2_sqsc_in[3]), .B(s2_sqsc_in[5]), .Z(
        s2_sqsc_out[6]) );
  XOR2_X1 s2_sqsc_0_U3 ( .A(s2_sqsc_out[0]), .B(s2_sqsc_in[0]), .Z(
        s2_sqsc_out[1]) );
  XOR2_X1 s2_sqsc_0_U2 ( .A(s2_sqsc_out[0]), .B(s2_sqsc_in[1]), .Z(
        s2_sqsc_out[3]) );
  XOR2_X1 s2_sqsc_0_U1 ( .A(s2_sqsc_in[0]), .B(s2_sqsc_in[2]), .Z(
        s2_sqsc_out[2]) );
  AOI221_X1 s2_mul1_2_2_U28 ( .B1(stage1Out[18]), .B2(stage1Out[19]), .C1(
        stage1Out[22]), .C2(stage1Out[23]), .A(s2_mul1_2_2_n73), .ZN(
        s2_mul1_2_2_n75) );
  OAI22_X1 s2_mul1_2_2_U27 ( .A1(stage1Out[18]), .A2(stage1Out[19]), .B1(
        stage1Out[23]), .B2(stage1Out[22]), .ZN(s2_mul1_2_2_n73) );
  XNOR2_X1 s2_mul1_2_2_U26 ( .A(s2_mul1_2_2_n72), .B(s2_mul1_2_2_n71), .ZN(
        s2_gf2_mul_out_2__2__1_) );
  NAND2_X1 s2_mul1_2_2_U25 ( .A1(stage1Out[17]), .A2(stage1Out[21]), .ZN(
        s2_mul1_2_2_n71) );
  XOR2_X1 s2_mul1_2_2_U24 ( .A(s2_mul1_2_2_n76), .B(s2_mul1_2_2_n70), .Z(
        s2_mul1_2_2_n72) );
  OAI22_X1 s2_mul1_2_2_U23 ( .A1(s2_mul1_2_2_n69), .A2(s2_mul1_2_2_n68), .B1(
        s2_mul1_2_2_n67), .B2(s2_mul1_2_2_n66), .ZN(s2_mul1_2_2_n76) );
  NAND2_X1 s2_mul1_2_2_U22 ( .A1(s2_mul1_2_2_n65), .A2(s2_mul1_2_2_n69), .ZN(
        s2_mul1_2_2_n66) );
  XNOR2_X1 s2_mul1_2_2_U21 ( .A(s2_mul1_2_2_n64), .B(s2_mul1_2_2_n63), .ZN(
        s2_mul1_2_2_n68) );
  NAND2_X1 s2_mul1_2_2_U20 ( .A1(s2_mul1_2_2_n65), .A2(s2_mul1_2_2_n67), .ZN(
        s2_mul1_2_2_n63) );
  INV_X1 s2_mul1_2_2_U19 ( .A(s2_mul1_2_2_n62), .ZN(s2_mul1_2_2_n69) );
  XNOR2_X1 s2_mul1_2_2_U18 ( .A(s2_mul1_2_2_n61), .B(s2_mul1_2_2_n60), .ZN(
        s2_gf2_mul_out_2__2__0_) );
  NAND2_X1 s2_mul1_2_2_U17 ( .A1(stage1Out[20]), .A2(stage1Out[16]), .ZN(
        s2_mul1_2_2_n60) );
  XOR2_X1 s2_mul1_2_2_U16 ( .A(s2_mul1_2_2_n70), .B(s2_mul1_2_2_n74), .Z(
        s2_mul1_2_2_n61) );
  XNOR2_X1 s2_mul1_2_2_U15 ( .A(s2_mul1_2_2_n59), .B(s2_mul1_2_2_n58), .ZN(
        s2_mul1_2_2_n74) );
  NAND2_X1 s2_mul1_2_2_U14 ( .A1(s2_mul1_2_2_n65), .A2(s2_mul1_2_2_n62), .ZN(
        s2_mul1_2_2_n58) );
  XOR2_X1 s2_mul1_2_2_U13 ( .A(stage1Out[17]), .B(stage1Out[19]), .Z(
        s2_mul1_2_2_n62) );
  XOR2_X1 s2_mul1_2_2_U12 ( .A(stage1Out[21]), .B(stage1Out[23]), .Z(
        s2_mul1_2_2_n65) );
  NOR2_X1 s2_mul1_2_2_U11 ( .A1(s2_mul1_2_2_n67), .A2(s2_mul1_2_2_n64), .ZN(
        s2_mul1_2_2_n59) );
  XNOR2_X1 s2_mul1_2_2_U10 ( .A(stage1Out[20]), .B(stage1Out[22]), .ZN(
        s2_mul1_2_2_n64) );
  XNOR2_X1 s2_mul1_2_2_U9 ( .A(stage1Out[16]), .B(stage1Out[18]), .ZN(
        s2_mul1_2_2_n67) );
  AOI221_X1 s2_mul1_2_2_U8 ( .B1(stage1Out[16]), .B2(stage1Out[17]), .C1(
        stage1Out[20]), .C2(stage1Out[21]), .A(s2_mul1_2_2_n57), .ZN(
        s2_mul1_2_2_n70) );
  OAI22_X1 s2_mul1_2_2_U7 ( .A1(stage1Out[16]), .A2(stage1Out[17]), .B1(
        stage1Out[21]), .B2(stage1Out[20]), .ZN(s2_mul1_2_2_n57) );
  XNOR2_X1 s2_mul1_2_2_U6 ( .A(s2_mul1_2_2_n55), .B(s2_mul1_2_2_n56), .ZN(
        s2_gf2_mul_out_2__2__3_) );
  XOR2_X1 s2_mul1_2_2_U5 ( .A(s2_mul1_2_2_n76), .B(s2_mul1_2_2_n75), .Z(
        s2_mul1_2_2_n56) );
  NAND2_X1 s2_mul1_2_2_U4 ( .A1(stage1Out[19]), .A2(stage1Out[23]), .ZN(
        s2_mul1_2_2_n55) );
  XNOR2_X1 s2_mul1_2_2_U3 ( .A(s2_mul1_2_2_n53), .B(s2_mul1_2_2_n54), .ZN(
        s2_gf2_mul_out_2__2__2_) );
  XOR2_X1 s2_mul1_2_2_U2 ( .A(s2_mul1_2_2_n74), .B(s2_mul1_2_2_n75), .Z(
        s2_mul1_2_2_n54) );
  NAND2_X1 s2_mul1_2_2_U1 ( .A1(stage1Out[18]), .A2(stage1Out[22]), .ZN(
        s2_mul1_2_2_n53) );
  XNOR2_X1 s2_mul1_2_1_U28 ( .A(s2_mul1_2_1_n76), .B(s2_mul1_2_1_n75), .ZN(
        s2_xorResult[23]) );
  NAND2_X1 s2_mul1_2_1_U27 ( .A1(stage1Out[11]), .A2(stage1Out[23]), .ZN(
        s2_mul1_2_1_n75) );
  XOR2_X1 s2_mul1_2_1_U26 ( .A(s2_mul1_2_1_n74), .B(s2_mul1_2_1_n73), .Z(
        s2_mul1_2_1_n76) );
  XNOR2_X1 s2_mul1_2_1_U25 ( .A(s2_mul1_2_1_n72), .B(s2_mul1_2_1_n71), .ZN(
        s2_xorResult[22]) );
  NAND2_X1 s2_mul1_2_1_U24 ( .A1(stage1Out[22]), .A2(stage1Out[10]), .ZN(
        s2_mul1_2_1_n71) );
  XOR2_X1 s2_mul1_2_1_U23 ( .A(s2_mul1_2_1_n73), .B(s2_mul1_2_1_n70), .Z(
        s2_mul1_2_1_n72) );
  AOI221_X1 s2_mul1_2_1_U22 ( .B1(stage1Out[10]), .B2(stage1Out[11]), .C1(
        stage1Out[22]), .C2(stage1Out[23]), .A(s2_mul1_2_1_n69), .ZN(
        s2_mul1_2_1_n73) );
  OAI22_X1 s2_mul1_2_1_U21 ( .A1(stage1Out[10]), .A2(stage1Out[11]), .B1(
        stage1Out[23]), .B2(stage1Out[22]), .ZN(s2_mul1_2_1_n69) );
  XNOR2_X1 s2_mul1_2_1_U20 ( .A(s2_mul1_2_1_n68), .B(s2_mul1_2_1_n67), .ZN(
        s2_xorResult[21]) );
  NAND2_X1 s2_mul1_2_1_U19 ( .A1(stage1Out[9]), .A2(stage1Out[21]), .ZN(
        s2_mul1_2_1_n67) );
  XOR2_X1 s2_mul1_2_1_U18 ( .A(s2_mul1_2_1_n74), .B(s2_mul1_2_1_n66), .Z(
        s2_mul1_2_1_n68) );
  OAI22_X1 s2_mul1_2_1_U17 ( .A1(s2_mul1_2_1_n65), .A2(s2_mul1_2_1_n64), .B1(
        s2_mul1_2_1_n63), .B2(s2_mul1_2_1_n62), .ZN(s2_mul1_2_1_n74) );
  NAND2_X1 s2_mul1_2_1_U16 ( .A1(s2_mul1_2_1_n61), .A2(s2_mul1_2_1_n65), .ZN(
        s2_mul1_2_1_n62) );
  XNOR2_X1 s2_mul1_2_1_U15 ( .A(s2_mul1_2_1_n60), .B(s2_mul1_2_1_n59), .ZN(
        s2_mul1_2_1_n64) );
  NAND2_X1 s2_mul1_2_1_U14 ( .A1(s2_mul1_2_1_n61), .A2(s2_mul1_2_1_n63), .ZN(
        s2_mul1_2_1_n59) );
  INV_X1 s2_mul1_2_1_U13 ( .A(s2_mul1_2_1_n58), .ZN(s2_mul1_2_1_n65) );
  XNOR2_X1 s2_mul1_2_1_U12 ( .A(s2_mul1_2_1_n57), .B(s2_mul1_2_1_n56), .ZN(
        s2_xorResult[20]) );
  NAND2_X1 s2_mul1_2_1_U11 ( .A1(stage1Out[20]), .A2(stage1Out[8]), .ZN(
        s2_mul1_2_1_n56) );
  XOR2_X1 s2_mul1_2_1_U10 ( .A(s2_mul1_2_1_n66), .B(s2_mul1_2_1_n70), .Z(
        s2_mul1_2_1_n57) );
  XNOR2_X1 s2_mul1_2_1_U9 ( .A(s2_mul1_2_1_n55), .B(s2_mul1_2_1_n54), .ZN(
        s2_mul1_2_1_n70) );
  NAND2_X1 s2_mul1_2_1_U8 ( .A1(s2_mul1_2_1_n61), .A2(s2_mul1_2_1_n58), .ZN(
        s2_mul1_2_1_n54) );
  XOR2_X1 s2_mul1_2_1_U7 ( .A(stage1Out[9]), .B(stage1Out[11]), .Z(
        s2_mul1_2_1_n58) );
  XOR2_X1 s2_mul1_2_1_U6 ( .A(stage1Out[21]), .B(stage1Out[23]), .Z(
        s2_mul1_2_1_n61) );
  NOR2_X1 s2_mul1_2_1_U5 ( .A1(s2_mul1_2_1_n63), .A2(s2_mul1_2_1_n60), .ZN(
        s2_mul1_2_1_n55) );
  XNOR2_X1 s2_mul1_2_1_U4 ( .A(stage1Out[20]), .B(stage1Out[22]), .ZN(
        s2_mul1_2_1_n60) );
  XNOR2_X1 s2_mul1_2_1_U3 ( .A(stage1Out[8]), .B(stage1Out[10]), .ZN(
        s2_mul1_2_1_n63) );
  AOI221_X1 s2_mul1_2_1_U2 ( .B1(stage1Out[8]), .B2(stage1Out[9]), .C1(
        stage1Out[20]), .C2(stage1Out[21]), .A(s2_mul1_2_1_n53), .ZN(
        s2_mul1_2_1_n66) );
  OAI22_X1 s2_mul1_2_1_U1 ( .A1(stage1Out[8]), .A2(stage1Out[9]), .B1(
        stage1Out[21]), .B2(stage1Out[20]), .ZN(s2_mul1_2_1_n53) );
  XNOR2_X1 s2_mul1_2_0_U28 ( .A(s2_mul1_2_0_n76), .B(s2_mul1_2_0_n75), .ZN(
        s2_xorResult[19]) );
  NAND2_X1 s2_mul1_2_0_U27 ( .A1(stage1Out[3]), .A2(stage1Out[23]), .ZN(
        s2_mul1_2_0_n75) );
  XOR2_X1 s2_mul1_2_0_U26 ( .A(s2_mul1_2_0_n74), .B(s2_mul1_2_0_n73), .Z(
        s2_mul1_2_0_n76) );
  XNOR2_X1 s2_mul1_2_0_U25 ( .A(s2_mul1_2_0_n72), .B(s2_mul1_2_0_n71), .ZN(
        s2_xorResult[18]) );
  NAND2_X1 s2_mul1_2_0_U24 ( .A1(stage1Out[22]), .A2(stage1Out[2]), .ZN(
        s2_mul1_2_0_n71) );
  XOR2_X1 s2_mul1_2_0_U23 ( .A(s2_mul1_2_0_n73), .B(s2_mul1_2_0_n70), .Z(
        s2_mul1_2_0_n72) );
  AOI221_X1 s2_mul1_2_0_U22 ( .B1(stage1Out[2]), .B2(stage1Out[3]), .C1(
        stage1Out[22]), .C2(stage1Out[23]), .A(s2_mul1_2_0_n69), .ZN(
        s2_mul1_2_0_n73) );
  OAI22_X1 s2_mul1_2_0_U21 ( .A1(stage1Out[2]), .A2(stage1Out[3]), .B1(
        stage1Out[23]), .B2(stage1Out[22]), .ZN(s2_mul1_2_0_n69) );
  XNOR2_X1 s2_mul1_2_0_U20 ( .A(s2_mul1_2_0_n68), .B(s2_mul1_2_0_n67), .ZN(
        s2_xorResult[17]) );
  NAND2_X1 s2_mul1_2_0_U19 ( .A1(stage1Out[1]), .A2(stage1Out[21]), .ZN(
        s2_mul1_2_0_n67) );
  XOR2_X1 s2_mul1_2_0_U18 ( .A(s2_mul1_2_0_n74), .B(s2_mul1_2_0_n66), .Z(
        s2_mul1_2_0_n68) );
  OAI22_X1 s2_mul1_2_0_U17 ( .A1(s2_mul1_2_0_n65), .A2(s2_mul1_2_0_n64), .B1(
        s2_mul1_2_0_n63), .B2(s2_mul1_2_0_n62), .ZN(s2_mul1_2_0_n74) );
  NAND2_X1 s2_mul1_2_0_U16 ( .A1(s2_mul1_2_0_n61), .A2(s2_mul1_2_0_n65), .ZN(
        s2_mul1_2_0_n62) );
  XNOR2_X1 s2_mul1_2_0_U15 ( .A(s2_mul1_2_0_n60), .B(s2_mul1_2_0_n59), .ZN(
        s2_mul1_2_0_n64) );
  NAND2_X1 s2_mul1_2_0_U14 ( .A1(s2_mul1_2_0_n61), .A2(s2_mul1_2_0_n63), .ZN(
        s2_mul1_2_0_n59) );
  INV_X1 s2_mul1_2_0_U13 ( .A(s2_mul1_2_0_n58), .ZN(s2_mul1_2_0_n65) );
  XNOR2_X1 s2_mul1_2_0_U12 ( .A(s2_mul1_2_0_n57), .B(s2_mul1_2_0_n56), .ZN(
        s2_xorResult[16]) );
  NAND2_X1 s2_mul1_2_0_U11 ( .A1(stage1Out[20]), .A2(stage1Out[0]), .ZN(
        s2_mul1_2_0_n56) );
  XOR2_X1 s2_mul1_2_0_U10 ( .A(s2_mul1_2_0_n66), .B(s2_mul1_2_0_n70), .Z(
        s2_mul1_2_0_n57) );
  XNOR2_X1 s2_mul1_2_0_U9 ( .A(s2_mul1_2_0_n55), .B(s2_mul1_2_0_n54), .ZN(
        s2_mul1_2_0_n70) );
  NAND2_X1 s2_mul1_2_0_U8 ( .A1(s2_mul1_2_0_n61), .A2(s2_mul1_2_0_n58), .ZN(
        s2_mul1_2_0_n54) );
  XOR2_X1 s2_mul1_2_0_U7 ( .A(stage1Out[1]), .B(stage1Out[3]), .Z(
        s2_mul1_2_0_n58) );
  XOR2_X1 s2_mul1_2_0_U6 ( .A(stage1Out[21]), .B(stage1Out[23]), .Z(
        s2_mul1_2_0_n61) );
  NOR2_X1 s2_mul1_2_0_U5 ( .A1(s2_mul1_2_0_n63), .A2(s2_mul1_2_0_n60), .ZN(
        s2_mul1_2_0_n55) );
  XNOR2_X1 s2_mul1_2_0_U4 ( .A(stage1Out[20]), .B(stage1Out[22]), .ZN(
        s2_mul1_2_0_n60) );
  XNOR2_X1 s2_mul1_2_0_U3 ( .A(stage1Out[0]), .B(stage1Out[2]), .ZN(
        s2_mul1_2_0_n63) );
  AOI221_X1 s2_mul1_2_0_U2 ( .B1(stage1Out[0]), .B2(stage1Out[1]), .C1(
        stage1Out[20]), .C2(stage1Out[21]), .A(s2_mul1_2_0_n53), .ZN(
        s2_mul1_2_0_n66) );
  OAI22_X1 s2_mul1_2_0_U1 ( .A1(stage1Out[0]), .A2(stage1Out[1]), .B1(
        stage1Out[21]), .B2(stage1Out[20]), .ZN(s2_mul1_2_0_n53) );
  XNOR2_X1 s2_mul1_1_2_U28 ( .A(s2_mul1_1_2_n76), .B(s2_mul1_1_2_n75), .ZN(
        s2_xorResult[15]) );
  NAND2_X1 s2_mul1_1_2_U27 ( .A1(stage1Out[19]), .A2(stage1Out[15]), .ZN(
        s2_mul1_1_2_n75) );
  XOR2_X1 s2_mul1_1_2_U26 ( .A(s2_mul1_1_2_n74), .B(s2_mul1_1_2_n73), .Z(
        s2_mul1_1_2_n76) );
  XNOR2_X1 s2_mul1_1_2_U25 ( .A(s2_mul1_1_2_n72), .B(s2_mul1_1_2_n71), .ZN(
        s2_xorResult[14]) );
  NAND2_X1 s2_mul1_1_2_U24 ( .A1(stage1Out[14]), .A2(stage1Out[18]), .ZN(
        s2_mul1_1_2_n71) );
  XOR2_X1 s2_mul1_1_2_U23 ( .A(s2_mul1_1_2_n73), .B(s2_mul1_1_2_n70), .Z(
        s2_mul1_1_2_n72) );
  AOI221_X1 s2_mul1_1_2_U22 ( .B1(stage1Out[18]), .B2(stage1Out[19]), .C1(
        stage1Out[14]), .C2(stage1Out[15]), .A(s2_mul1_1_2_n69), .ZN(
        s2_mul1_1_2_n73) );
  OAI22_X1 s2_mul1_1_2_U21 ( .A1(stage1Out[18]), .A2(stage1Out[19]), .B1(
        stage1Out[15]), .B2(stage1Out[14]), .ZN(s2_mul1_1_2_n69) );
  XNOR2_X1 s2_mul1_1_2_U20 ( .A(s2_mul1_1_2_n68), .B(s2_mul1_1_2_n67), .ZN(
        s2_xorResult[13]) );
  NAND2_X1 s2_mul1_1_2_U19 ( .A1(stage1Out[17]), .A2(stage1Out[13]), .ZN(
        s2_mul1_1_2_n67) );
  XOR2_X1 s2_mul1_1_2_U18 ( .A(s2_mul1_1_2_n74), .B(s2_mul1_1_2_n66), .Z(
        s2_mul1_1_2_n68) );
  OAI22_X1 s2_mul1_1_2_U17 ( .A1(s2_mul1_1_2_n65), .A2(s2_mul1_1_2_n64), .B1(
        s2_mul1_1_2_n63), .B2(s2_mul1_1_2_n62), .ZN(s2_mul1_1_2_n74) );
  NAND2_X1 s2_mul1_1_2_U16 ( .A1(s2_mul1_1_2_n61), .A2(s2_mul1_1_2_n65), .ZN(
        s2_mul1_1_2_n62) );
  XNOR2_X1 s2_mul1_1_2_U15 ( .A(s2_mul1_1_2_n60), .B(s2_mul1_1_2_n59), .ZN(
        s2_mul1_1_2_n64) );
  NAND2_X1 s2_mul1_1_2_U14 ( .A1(s2_mul1_1_2_n61), .A2(s2_mul1_1_2_n63), .ZN(
        s2_mul1_1_2_n59) );
  INV_X1 s2_mul1_1_2_U13 ( .A(s2_mul1_1_2_n58), .ZN(s2_mul1_1_2_n65) );
  XNOR2_X1 s2_mul1_1_2_U12 ( .A(s2_mul1_1_2_n57), .B(s2_mul1_1_2_n56), .ZN(
        s2_xorResult[12]) );
  NAND2_X1 s2_mul1_1_2_U11 ( .A1(stage1Out[12]), .A2(stage1Out[16]), .ZN(
        s2_mul1_1_2_n56) );
  XOR2_X1 s2_mul1_1_2_U10 ( .A(s2_mul1_1_2_n66), .B(s2_mul1_1_2_n70), .Z(
        s2_mul1_1_2_n57) );
  XNOR2_X1 s2_mul1_1_2_U9 ( .A(s2_mul1_1_2_n55), .B(s2_mul1_1_2_n54), .ZN(
        s2_mul1_1_2_n70) );
  NAND2_X1 s2_mul1_1_2_U8 ( .A1(s2_mul1_1_2_n61), .A2(s2_mul1_1_2_n58), .ZN(
        s2_mul1_1_2_n54) );
  XOR2_X1 s2_mul1_1_2_U7 ( .A(stage1Out[17]), .B(stage1Out[19]), .Z(
        s2_mul1_1_2_n58) );
  XOR2_X1 s2_mul1_1_2_U6 ( .A(stage1Out[13]), .B(stage1Out[15]), .Z(
        s2_mul1_1_2_n61) );
  NOR2_X1 s2_mul1_1_2_U5 ( .A1(s2_mul1_1_2_n63), .A2(s2_mul1_1_2_n60), .ZN(
        s2_mul1_1_2_n55) );
  XNOR2_X1 s2_mul1_1_2_U4 ( .A(stage1Out[12]), .B(stage1Out[14]), .ZN(
        s2_mul1_1_2_n60) );
  XNOR2_X1 s2_mul1_1_2_U3 ( .A(stage1Out[16]), .B(stage1Out[18]), .ZN(
        s2_mul1_1_2_n63) );
  AOI221_X1 s2_mul1_1_2_U2 ( .B1(stage1Out[16]), .B2(stage1Out[17]), .C1(
        stage1Out[12]), .C2(stage1Out[13]), .A(s2_mul1_1_2_n53), .ZN(
        s2_mul1_1_2_n66) );
  OAI22_X1 s2_mul1_1_2_U1 ( .A1(stage1Out[16]), .A2(stage1Out[17]), .B1(
        stage1Out[13]), .B2(stage1Out[12]), .ZN(s2_mul1_1_2_n53) );
  AOI221_X1 s2_mul1_1_1_U28 ( .B1(stage1Out[10]), .B2(stage1Out[11]), .C1(
        stage1Out[14]), .C2(stage1Out[15]), .A(s2_mul1_1_1_n73), .ZN(
        s2_mul1_1_1_n75) );
  OAI22_X1 s2_mul1_1_1_U27 ( .A1(stage1Out[10]), .A2(stage1Out[11]), .B1(
        stage1Out[15]), .B2(stage1Out[14]), .ZN(s2_mul1_1_1_n73) );
  XNOR2_X1 s2_mul1_1_1_U26 ( .A(s2_mul1_1_1_n72), .B(s2_mul1_1_1_n71), .ZN(
        s2_gf2_mul_out_1__1__1_) );
  NAND2_X1 s2_mul1_1_1_U25 ( .A1(stage1Out[9]), .A2(stage1Out[13]), .ZN(
        s2_mul1_1_1_n71) );
  XOR2_X1 s2_mul1_1_1_U24 ( .A(s2_mul1_1_1_n76), .B(s2_mul1_1_1_n70), .Z(
        s2_mul1_1_1_n72) );
  OAI22_X1 s2_mul1_1_1_U23 ( .A1(s2_mul1_1_1_n69), .A2(s2_mul1_1_1_n68), .B1(
        s2_mul1_1_1_n67), .B2(s2_mul1_1_1_n66), .ZN(s2_mul1_1_1_n76) );
  NAND2_X1 s2_mul1_1_1_U22 ( .A1(s2_mul1_1_1_n65), .A2(s2_mul1_1_1_n69), .ZN(
        s2_mul1_1_1_n66) );
  XNOR2_X1 s2_mul1_1_1_U21 ( .A(s2_mul1_1_1_n64), .B(s2_mul1_1_1_n63), .ZN(
        s2_mul1_1_1_n68) );
  NAND2_X1 s2_mul1_1_1_U20 ( .A1(s2_mul1_1_1_n65), .A2(s2_mul1_1_1_n67), .ZN(
        s2_mul1_1_1_n63) );
  INV_X1 s2_mul1_1_1_U19 ( .A(s2_mul1_1_1_n62), .ZN(s2_mul1_1_1_n69) );
  XNOR2_X1 s2_mul1_1_1_U18 ( .A(s2_mul1_1_1_n61), .B(s2_mul1_1_1_n60), .ZN(
        s2_gf2_mul_out_1__1__0_) );
  NAND2_X1 s2_mul1_1_1_U17 ( .A1(stage1Out[12]), .A2(stage1Out[8]), .ZN(
        s2_mul1_1_1_n60) );
  XOR2_X1 s2_mul1_1_1_U16 ( .A(s2_mul1_1_1_n70), .B(s2_mul1_1_1_n74), .Z(
        s2_mul1_1_1_n61) );
  XNOR2_X1 s2_mul1_1_1_U15 ( .A(s2_mul1_1_1_n59), .B(s2_mul1_1_1_n58), .ZN(
        s2_mul1_1_1_n74) );
  NAND2_X1 s2_mul1_1_1_U14 ( .A1(s2_mul1_1_1_n65), .A2(s2_mul1_1_1_n62), .ZN(
        s2_mul1_1_1_n58) );
  XOR2_X1 s2_mul1_1_1_U13 ( .A(stage1Out[9]), .B(stage1Out[11]), .Z(
        s2_mul1_1_1_n62) );
  XOR2_X1 s2_mul1_1_1_U12 ( .A(stage1Out[13]), .B(stage1Out[15]), .Z(
        s2_mul1_1_1_n65) );
  NOR2_X1 s2_mul1_1_1_U11 ( .A1(s2_mul1_1_1_n67), .A2(s2_mul1_1_1_n64), .ZN(
        s2_mul1_1_1_n59) );
  XNOR2_X1 s2_mul1_1_1_U10 ( .A(stage1Out[12]), .B(stage1Out[14]), .ZN(
        s2_mul1_1_1_n64) );
  XNOR2_X1 s2_mul1_1_1_U9 ( .A(stage1Out[8]), .B(stage1Out[10]), .ZN(
        s2_mul1_1_1_n67) );
  AOI221_X1 s2_mul1_1_1_U8 ( .B1(stage1Out[8]), .B2(stage1Out[9]), .C1(
        stage1Out[12]), .C2(stage1Out[13]), .A(s2_mul1_1_1_n57), .ZN(
        s2_mul1_1_1_n70) );
  OAI22_X1 s2_mul1_1_1_U7 ( .A1(stage1Out[8]), .A2(stage1Out[9]), .B1(
        stage1Out[13]), .B2(stage1Out[12]), .ZN(s2_mul1_1_1_n57) );
  XNOR2_X1 s2_mul1_1_1_U6 ( .A(s2_mul1_1_1_n55), .B(s2_mul1_1_1_n56), .ZN(
        s2_gf2_mul_out_1__1__3_) );
  XOR2_X1 s2_mul1_1_1_U5 ( .A(s2_mul1_1_1_n76), .B(s2_mul1_1_1_n75), .Z(
        s2_mul1_1_1_n56) );
  NAND2_X1 s2_mul1_1_1_U4 ( .A1(stage1Out[11]), .A2(stage1Out[15]), .ZN(
        s2_mul1_1_1_n55) );
  XNOR2_X1 s2_mul1_1_1_U3 ( .A(s2_mul1_1_1_n53), .B(s2_mul1_1_1_n54), .ZN(
        s2_gf2_mul_out_1__1__2_) );
  XOR2_X1 s2_mul1_1_1_U2 ( .A(s2_mul1_1_1_n74), .B(s2_mul1_1_1_n75), .Z(
        s2_mul1_1_1_n54) );
  NAND2_X1 s2_mul1_1_1_U1 ( .A1(stage1Out[10]), .A2(stage1Out[14]), .ZN(
        s2_mul1_1_1_n53) );
  XNOR2_X1 s2_mul1_1_0_U28 ( .A(s2_mul1_1_0_n76), .B(s2_mul1_1_0_n75), .ZN(
        s2_xorResult[11]) );
  NAND2_X1 s2_mul1_1_0_U27 ( .A1(stage1Out[3]), .A2(stage1Out[15]), .ZN(
        s2_mul1_1_0_n75) );
  XOR2_X1 s2_mul1_1_0_U26 ( .A(s2_mul1_1_0_n74), .B(s2_mul1_1_0_n73), .Z(
        s2_mul1_1_0_n76) );
  XNOR2_X1 s2_mul1_1_0_U25 ( .A(s2_mul1_1_0_n72), .B(s2_mul1_1_0_n71), .ZN(
        s2_xorResult[10]) );
  NAND2_X1 s2_mul1_1_0_U24 ( .A1(stage1Out[14]), .A2(stage1Out[2]), .ZN(
        s2_mul1_1_0_n71) );
  XOR2_X1 s2_mul1_1_0_U23 ( .A(s2_mul1_1_0_n73), .B(s2_mul1_1_0_n70), .Z(
        s2_mul1_1_0_n72) );
  AOI221_X1 s2_mul1_1_0_U22 ( .B1(stage1Out[2]), .B2(stage1Out[3]), .C1(
        stage1Out[14]), .C2(stage1Out[15]), .A(s2_mul1_1_0_n69), .ZN(
        s2_mul1_1_0_n73) );
  OAI22_X1 s2_mul1_1_0_U21 ( .A1(stage1Out[2]), .A2(stage1Out[3]), .B1(
        stage1Out[15]), .B2(stage1Out[14]), .ZN(s2_mul1_1_0_n69) );
  XNOR2_X1 s2_mul1_1_0_U20 ( .A(s2_mul1_1_0_n68), .B(s2_mul1_1_0_n67), .ZN(
        s2_xorResult[9]) );
  NAND2_X1 s2_mul1_1_0_U19 ( .A1(stage1Out[1]), .A2(stage1Out[13]), .ZN(
        s2_mul1_1_0_n67) );
  XOR2_X1 s2_mul1_1_0_U18 ( .A(s2_mul1_1_0_n74), .B(s2_mul1_1_0_n66), .Z(
        s2_mul1_1_0_n68) );
  OAI22_X1 s2_mul1_1_0_U17 ( .A1(s2_mul1_1_0_n65), .A2(s2_mul1_1_0_n64), .B1(
        s2_mul1_1_0_n63), .B2(s2_mul1_1_0_n62), .ZN(s2_mul1_1_0_n74) );
  NAND2_X1 s2_mul1_1_0_U16 ( .A1(s2_mul1_1_0_n61), .A2(s2_mul1_1_0_n65), .ZN(
        s2_mul1_1_0_n62) );
  XNOR2_X1 s2_mul1_1_0_U15 ( .A(s2_mul1_1_0_n60), .B(s2_mul1_1_0_n59), .ZN(
        s2_mul1_1_0_n64) );
  NAND2_X1 s2_mul1_1_0_U14 ( .A1(s2_mul1_1_0_n61), .A2(s2_mul1_1_0_n63), .ZN(
        s2_mul1_1_0_n59) );
  INV_X1 s2_mul1_1_0_U13 ( .A(s2_mul1_1_0_n58), .ZN(s2_mul1_1_0_n65) );
  XNOR2_X1 s2_mul1_1_0_U12 ( .A(s2_mul1_1_0_n57), .B(s2_mul1_1_0_n56), .ZN(
        s2_xorResult[8]) );
  NAND2_X1 s2_mul1_1_0_U11 ( .A1(stage1Out[12]), .A2(stage1Out[0]), .ZN(
        s2_mul1_1_0_n56) );
  XOR2_X1 s2_mul1_1_0_U10 ( .A(s2_mul1_1_0_n66), .B(s2_mul1_1_0_n70), .Z(
        s2_mul1_1_0_n57) );
  XNOR2_X1 s2_mul1_1_0_U9 ( .A(s2_mul1_1_0_n55), .B(s2_mul1_1_0_n54), .ZN(
        s2_mul1_1_0_n70) );
  NAND2_X1 s2_mul1_1_0_U8 ( .A1(s2_mul1_1_0_n61), .A2(s2_mul1_1_0_n58), .ZN(
        s2_mul1_1_0_n54) );
  XOR2_X1 s2_mul1_1_0_U7 ( .A(stage1Out[1]), .B(stage1Out[3]), .Z(
        s2_mul1_1_0_n58) );
  XOR2_X1 s2_mul1_1_0_U6 ( .A(stage1Out[13]), .B(stage1Out[15]), .Z(
        s2_mul1_1_0_n61) );
  NOR2_X1 s2_mul1_1_0_U5 ( .A1(s2_mul1_1_0_n63), .A2(s2_mul1_1_0_n60), .ZN(
        s2_mul1_1_0_n55) );
  XNOR2_X1 s2_mul1_1_0_U4 ( .A(stage1Out[12]), .B(stage1Out[14]), .ZN(
        s2_mul1_1_0_n60) );
  XNOR2_X1 s2_mul1_1_0_U3 ( .A(stage1Out[0]), .B(stage1Out[2]), .ZN(
        s2_mul1_1_0_n63) );
  AOI221_X1 s2_mul1_1_0_U2 ( .B1(stage1Out[0]), .B2(stage1Out[1]), .C1(
        stage1Out[12]), .C2(stage1Out[13]), .A(s2_mul1_1_0_n53), .ZN(
        s2_mul1_1_0_n66) );
  OAI22_X1 s2_mul1_1_0_U1 ( .A1(stage1Out[0]), .A2(stage1Out[1]), .B1(
        stage1Out[13]), .B2(stage1Out[12]), .ZN(s2_mul1_1_0_n53) );
  XNOR2_X1 s2_mul1_0_2_U28 ( .A(s2_mul1_0_2_n76), .B(s2_mul1_0_2_n75), .ZN(
        s2_xorResult[7]) );
  NAND2_X1 s2_mul1_0_2_U27 ( .A1(stage1Out[19]), .A2(stage1Out[7]), .ZN(
        s2_mul1_0_2_n75) );
  XOR2_X1 s2_mul1_0_2_U26 ( .A(s2_mul1_0_2_n74), .B(s2_mul1_0_2_n73), .Z(
        s2_mul1_0_2_n76) );
  XNOR2_X1 s2_mul1_0_2_U25 ( .A(s2_mul1_0_2_n72), .B(s2_mul1_0_2_n71), .ZN(
        s2_xorResult[6]) );
  NAND2_X1 s2_mul1_0_2_U24 ( .A1(stage1Out[6]), .A2(stage1Out[18]), .ZN(
        s2_mul1_0_2_n71) );
  XOR2_X1 s2_mul1_0_2_U23 ( .A(s2_mul1_0_2_n73), .B(s2_mul1_0_2_n70), .Z(
        s2_mul1_0_2_n72) );
  AOI221_X1 s2_mul1_0_2_U22 ( .B1(stage1Out[18]), .B2(stage1Out[19]), .C1(
        stage1Out[6]), .C2(stage1Out[7]), .A(s2_mul1_0_2_n69), .ZN(
        s2_mul1_0_2_n73) );
  OAI22_X1 s2_mul1_0_2_U21 ( .A1(stage1Out[18]), .A2(stage1Out[19]), .B1(
        stage1Out[7]), .B2(stage1Out[6]), .ZN(s2_mul1_0_2_n69) );
  XNOR2_X1 s2_mul1_0_2_U20 ( .A(s2_mul1_0_2_n68), .B(s2_mul1_0_2_n67), .ZN(
        s2_xorResult[5]) );
  NAND2_X1 s2_mul1_0_2_U19 ( .A1(stage1Out[17]), .A2(stage1Out[5]), .ZN(
        s2_mul1_0_2_n67) );
  XOR2_X1 s2_mul1_0_2_U18 ( .A(s2_mul1_0_2_n74), .B(s2_mul1_0_2_n66), .Z(
        s2_mul1_0_2_n68) );
  OAI22_X1 s2_mul1_0_2_U17 ( .A1(s2_mul1_0_2_n65), .A2(s2_mul1_0_2_n64), .B1(
        s2_mul1_0_2_n63), .B2(s2_mul1_0_2_n62), .ZN(s2_mul1_0_2_n74) );
  NAND2_X1 s2_mul1_0_2_U16 ( .A1(s2_mul1_0_2_n61), .A2(s2_mul1_0_2_n65), .ZN(
        s2_mul1_0_2_n62) );
  XNOR2_X1 s2_mul1_0_2_U15 ( .A(s2_mul1_0_2_n60), .B(s2_mul1_0_2_n59), .ZN(
        s2_mul1_0_2_n64) );
  NAND2_X1 s2_mul1_0_2_U14 ( .A1(s2_mul1_0_2_n61), .A2(s2_mul1_0_2_n63), .ZN(
        s2_mul1_0_2_n59) );
  INV_X1 s2_mul1_0_2_U13 ( .A(s2_mul1_0_2_n58), .ZN(s2_mul1_0_2_n65) );
  XNOR2_X1 s2_mul1_0_2_U12 ( .A(s2_mul1_0_2_n57), .B(s2_mul1_0_2_n56), .ZN(
        s2_xorResult[4]) );
  NAND2_X1 s2_mul1_0_2_U11 ( .A1(stage1Out[4]), .A2(stage1Out[16]), .ZN(
        s2_mul1_0_2_n56) );
  XOR2_X1 s2_mul1_0_2_U10 ( .A(s2_mul1_0_2_n66), .B(s2_mul1_0_2_n70), .Z(
        s2_mul1_0_2_n57) );
  XNOR2_X1 s2_mul1_0_2_U9 ( .A(s2_mul1_0_2_n55), .B(s2_mul1_0_2_n54), .ZN(
        s2_mul1_0_2_n70) );
  NAND2_X1 s2_mul1_0_2_U8 ( .A1(s2_mul1_0_2_n61), .A2(s2_mul1_0_2_n58), .ZN(
        s2_mul1_0_2_n54) );
  XOR2_X1 s2_mul1_0_2_U7 ( .A(stage1Out[17]), .B(stage1Out[19]), .Z(
        s2_mul1_0_2_n58) );
  XOR2_X1 s2_mul1_0_2_U6 ( .A(stage1Out[5]), .B(stage1Out[7]), .Z(
        s2_mul1_0_2_n61) );
  NOR2_X1 s2_mul1_0_2_U5 ( .A1(s2_mul1_0_2_n63), .A2(s2_mul1_0_2_n60), .ZN(
        s2_mul1_0_2_n55) );
  XNOR2_X1 s2_mul1_0_2_U4 ( .A(stage1Out[4]), .B(stage1Out[6]), .ZN(
        s2_mul1_0_2_n60) );
  XNOR2_X1 s2_mul1_0_2_U3 ( .A(stage1Out[16]), .B(stage1Out[18]), .ZN(
        s2_mul1_0_2_n63) );
  AOI221_X1 s2_mul1_0_2_U2 ( .B1(stage1Out[16]), .B2(stage1Out[17]), .C1(
        stage1Out[4]), .C2(stage1Out[5]), .A(s2_mul1_0_2_n53), .ZN(
        s2_mul1_0_2_n66) );
  OAI22_X1 s2_mul1_0_2_U1 ( .A1(stage1Out[16]), .A2(stage1Out[17]), .B1(
        stage1Out[5]), .B2(stage1Out[4]), .ZN(s2_mul1_0_2_n53) );
  XNOR2_X1 s2_mul1_0_1_U28 ( .A(s2_mul1_0_1_n76), .B(s2_mul1_0_1_n75), .ZN(
        s2_xorResult[3]) );
  NAND2_X1 s2_mul1_0_1_U27 ( .A1(stage1Out[11]), .A2(stage1Out[7]), .ZN(
        s2_mul1_0_1_n75) );
  XOR2_X1 s2_mul1_0_1_U26 ( .A(s2_mul1_0_1_n74), .B(s2_mul1_0_1_n73), .Z(
        s2_mul1_0_1_n76) );
  XNOR2_X1 s2_mul1_0_1_U25 ( .A(s2_mul1_0_1_n72), .B(s2_mul1_0_1_n71), .ZN(
        s2_xorResult[2]) );
  NAND2_X1 s2_mul1_0_1_U24 ( .A1(stage1Out[6]), .A2(stage1Out[10]), .ZN(
        s2_mul1_0_1_n71) );
  XOR2_X1 s2_mul1_0_1_U23 ( .A(s2_mul1_0_1_n73), .B(s2_mul1_0_1_n70), .Z(
        s2_mul1_0_1_n72) );
  AOI221_X1 s2_mul1_0_1_U22 ( .B1(stage1Out[10]), .B2(stage1Out[11]), .C1(
        stage1Out[6]), .C2(stage1Out[7]), .A(s2_mul1_0_1_n69), .ZN(
        s2_mul1_0_1_n73) );
  OAI22_X1 s2_mul1_0_1_U21 ( .A1(stage1Out[10]), .A2(stage1Out[11]), .B1(
        stage1Out[7]), .B2(stage1Out[6]), .ZN(s2_mul1_0_1_n69) );
  XNOR2_X1 s2_mul1_0_1_U20 ( .A(s2_mul1_0_1_n68), .B(s2_mul1_0_1_n67), .ZN(
        s2_xorResult[1]) );
  NAND2_X1 s2_mul1_0_1_U19 ( .A1(stage1Out[9]), .A2(stage1Out[5]), .ZN(
        s2_mul1_0_1_n67) );
  XOR2_X1 s2_mul1_0_1_U18 ( .A(s2_mul1_0_1_n74), .B(s2_mul1_0_1_n66), .Z(
        s2_mul1_0_1_n68) );
  OAI22_X1 s2_mul1_0_1_U17 ( .A1(s2_mul1_0_1_n65), .A2(s2_mul1_0_1_n64), .B1(
        s2_mul1_0_1_n63), .B2(s2_mul1_0_1_n62), .ZN(s2_mul1_0_1_n74) );
  NAND2_X1 s2_mul1_0_1_U16 ( .A1(s2_mul1_0_1_n61), .A2(s2_mul1_0_1_n65), .ZN(
        s2_mul1_0_1_n62) );
  XNOR2_X1 s2_mul1_0_1_U15 ( .A(s2_mul1_0_1_n60), .B(s2_mul1_0_1_n59), .ZN(
        s2_mul1_0_1_n64) );
  NAND2_X1 s2_mul1_0_1_U14 ( .A1(s2_mul1_0_1_n61), .A2(s2_mul1_0_1_n63), .ZN(
        s2_mul1_0_1_n59) );
  INV_X1 s2_mul1_0_1_U13 ( .A(s2_mul1_0_1_n58), .ZN(s2_mul1_0_1_n65) );
  XNOR2_X1 s2_mul1_0_1_U12 ( .A(s2_mul1_0_1_n57), .B(s2_mul1_0_1_n56), .ZN(
        s2_xorResult[0]) );
  NAND2_X1 s2_mul1_0_1_U11 ( .A1(stage1Out[4]), .A2(stage1Out[8]), .ZN(
        s2_mul1_0_1_n56) );
  XOR2_X1 s2_mul1_0_1_U10 ( .A(s2_mul1_0_1_n66), .B(s2_mul1_0_1_n70), .Z(
        s2_mul1_0_1_n57) );
  XNOR2_X1 s2_mul1_0_1_U9 ( .A(s2_mul1_0_1_n55), .B(s2_mul1_0_1_n54), .ZN(
        s2_mul1_0_1_n70) );
  NAND2_X1 s2_mul1_0_1_U8 ( .A1(s2_mul1_0_1_n61), .A2(s2_mul1_0_1_n58), .ZN(
        s2_mul1_0_1_n54) );
  XOR2_X1 s2_mul1_0_1_U7 ( .A(stage1Out[9]), .B(stage1Out[11]), .Z(
        s2_mul1_0_1_n58) );
  XOR2_X1 s2_mul1_0_1_U6 ( .A(stage1Out[5]), .B(stage1Out[7]), .Z(
        s2_mul1_0_1_n61) );
  NOR2_X1 s2_mul1_0_1_U5 ( .A1(s2_mul1_0_1_n63), .A2(s2_mul1_0_1_n60), .ZN(
        s2_mul1_0_1_n55) );
  XNOR2_X1 s2_mul1_0_1_U4 ( .A(stage1Out[4]), .B(stage1Out[6]), .ZN(
        s2_mul1_0_1_n60) );
  XNOR2_X1 s2_mul1_0_1_U3 ( .A(stage1Out[8]), .B(stage1Out[10]), .ZN(
        s2_mul1_0_1_n63) );
  AOI221_X1 s2_mul1_0_1_U2 ( .B1(stage1Out[8]), .B2(stage1Out[9]), .C1(
        stage1Out[4]), .C2(stage1Out[5]), .A(s2_mul1_0_1_n53), .ZN(
        s2_mul1_0_1_n66) );
  OAI22_X1 s2_mul1_0_1_U1 ( .A1(stage1Out[8]), .A2(stage1Out[9]), .B1(
        stage1Out[5]), .B2(stage1Out[4]), .ZN(s2_mul1_0_1_n53) );
  AOI221_X1 s2_mul1_0_0_U28 ( .B1(stage1Out[2]), .B2(stage1Out[3]), .C1(
        stage1Out[6]), .C2(stage1Out[7]), .A(s2_mul1_0_0_n73), .ZN(
        s2_mul1_0_0_n75) );
  OAI22_X1 s2_mul1_0_0_U27 ( .A1(stage1Out[2]), .A2(stage1Out[3]), .B1(
        stage1Out[7]), .B2(stage1Out[6]), .ZN(s2_mul1_0_0_n73) );
  XNOR2_X1 s2_mul1_0_0_U26 ( .A(s2_mul1_0_0_n72), .B(s2_mul1_0_0_n71), .ZN(
        s2_gf2_mul_out_0__0__1_) );
  NAND2_X1 s2_mul1_0_0_U25 ( .A1(stage1Out[1]), .A2(stage1Out[5]), .ZN(
        s2_mul1_0_0_n71) );
  XOR2_X1 s2_mul1_0_0_U24 ( .A(s2_mul1_0_0_n76), .B(s2_mul1_0_0_n70), .Z(
        s2_mul1_0_0_n72) );
  OAI22_X1 s2_mul1_0_0_U23 ( .A1(s2_mul1_0_0_n69), .A2(s2_mul1_0_0_n68), .B1(
        s2_mul1_0_0_n67), .B2(s2_mul1_0_0_n66), .ZN(s2_mul1_0_0_n76) );
  NAND2_X1 s2_mul1_0_0_U22 ( .A1(s2_mul1_0_0_n65), .A2(s2_mul1_0_0_n69), .ZN(
        s2_mul1_0_0_n66) );
  XNOR2_X1 s2_mul1_0_0_U21 ( .A(s2_mul1_0_0_n64), .B(s2_mul1_0_0_n63), .ZN(
        s2_mul1_0_0_n68) );
  NAND2_X1 s2_mul1_0_0_U20 ( .A1(s2_mul1_0_0_n65), .A2(s2_mul1_0_0_n67), .ZN(
        s2_mul1_0_0_n63) );
  INV_X1 s2_mul1_0_0_U19 ( .A(s2_mul1_0_0_n62), .ZN(s2_mul1_0_0_n69) );
  XNOR2_X1 s2_mul1_0_0_U18 ( .A(s2_mul1_0_0_n61), .B(s2_mul1_0_0_n60), .ZN(
        s2_gf2_mul_out_0__0__0_) );
  NAND2_X1 s2_mul1_0_0_U17 ( .A1(stage1Out[4]), .A2(stage1Out[0]), .ZN(
        s2_mul1_0_0_n60) );
  XOR2_X1 s2_mul1_0_0_U16 ( .A(s2_mul1_0_0_n70), .B(s2_mul1_0_0_n74), .Z(
        s2_mul1_0_0_n61) );
  XNOR2_X1 s2_mul1_0_0_U15 ( .A(s2_mul1_0_0_n59), .B(s2_mul1_0_0_n58), .ZN(
        s2_mul1_0_0_n74) );
  NAND2_X1 s2_mul1_0_0_U14 ( .A1(s2_mul1_0_0_n65), .A2(s2_mul1_0_0_n62), .ZN(
        s2_mul1_0_0_n58) );
  XOR2_X1 s2_mul1_0_0_U13 ( .A(stage1Out[1]), .B(stage1Out[3]), .Z(
        s2_mul1_0_0_n62) );
  XOR2_X1 s2_mul1_0_0_U12 ( .A(stage1Out[5]), .B(stage1Out[7]), .Z(
        s2_mul1_0_0_n65) );
  NOR2_X1 s2_mul1_0_0_U11 ( .A1(s2_mul1_0_0_n67), .A2(s2_mul1_0_0_n64), .ZN(
        s2_mul1_0_0_n59) );
  XNOR2_X1 s2_mul1_0_0_U10 ( .A(stage1Out[4]), .B(stage1Out[6]), .ZN(
        s2_mul1_0_0_n64) );
  XNOR2_X1 s2_mul1_0_0_U9 ( .A(stage1Out[0]), .B(stage1Out[2]), .ZN(
        s2_mul1_0_0_n67) );
  AOI221_X1 s2_mul1_0_0_U8 ( .B1(stage1Out[0]), .B2(stage1Out[1]), .C1(
        stage1Out[4]), .C2(stage1Out[5]), .A(s2_mul1_0_0_n57), .ZN(
        s2_mul1_0_0_n70) );
  OAI22_X1 s2_mul1_0_0_U7 ( .A1(stage1Out[0]), .A2(stage1Out[1]), .B1(
        stage1Out[5]), .B2(stage1Out[4]), .ZN(s2_mul1_0_0_n57) );
  XNOR2_X1 s2_mul1_0_0_U6 ( .A(s2_mul1_0_0_n55), .B(s2_mul1_0_0_n56), .ZN(
        s2_gf2_mul_out_0__0__3_) );
  XOR2_X1 s2_mul1_0_0_U5 ( .A(s2_mul1_0_0_n76), .B(s2_mul1_0_0_n75), .Z(
        s2_mul1_0_0_n56) );
  NAND2_X1 s2_mul1_0_0_U4 ( .A1(stage1Out[3]), .A2(stage1Out[7]), .ZN(
        s2_mul1_0_0_n55) );
  XNOR2_X1 s2_mul1_0_0_U3 ( .A(s2_mul1_0_0_n53), .B(s2_mul1_0_0_n54), .ZN(
        s2_gf2_mul_out_0__0__2_) );
  XOR2_X1 s2_mul1_0_0_U2 ( .A(s2_mul1_0_0_n74), .B(s2_mul1_0_0_n75), .Z(
        s2_mul1_0_0_n54) );
  NAND2_X1 s2_mul1_0_0_U1 ( .A1(stage1Out[2]), .A2(stage1Out[6]), .ZN(
        s2_mul1_0_0_n53) );
  XOR2_X1 s2_compr_0_0_U4 ( .A(s2_regOut_0__1__3_), .B(s2_regOut_0__2__3_), 
        .Z(s2_chain_0__1__3_) );
  XOR2_X1 s2_compr_0_0_U3 ( .A(s2_regOut_0__1__2_), .B(s2_regOut_0__2__2_), 
        .Z(s2_chain_0__1__2_) );
  XOR2_X1 s2_compr_0_0_U2 ( .A(s2_regOut_0__1__1_), .B(s2_regOut_0__2__1_), 
        .Z(s2_chain_0__1__1_) );
  XOR2_X1 s2_compr_0_0_U1 ( .A(s2_regOut_0__1__0_), .B(s2_regOut_0__2__0_), 
        .Z(s2_chain_0__1__0_) );
  XOR2_X2 s2_compr_0_1_U4 ( .A(s2_chain_0__1__1_), .B(s2_regOut_0__3__1_), .Z(
        stage2Out[5]) );
  XOR2_X2 s2_compr_0_1_U3 ( .A(s2_chain_0__1__0_), .B(s2_regOut_0__3__0_), .Z(
        stage2Out[4]) );
  XOR2_X2 s2_compr_0_1_U2 ( .A(s2_chain_0__1__2_), .B(s2_regOut_0__3__2_), .Z(
        stage2Out[6]) );
  XOR2_X2 s2_compr_0_1_U1 ( .A(s2_chain_0__1__3_), .B(s2_regOut_0__3__3_), .Z(
        stage2Out[7]) );
  XOR2_X1 s2_compr_1_0_U4 ( .A(s2_regOut_1__1__3_), .B(s2_regOut_1__2__3_), 
        .Z(s2_chain_1__1__3_) );
  XOR2_X1 s2_compr_1_0_U3 ( .A(s2_regOut_1__1__2_), .B(s2_regOut_1__2__2_), 
        .Z(s2_chain_1__1__2_) );
  XOR2_X1 s2_compr_1_0_U2 ( .A(s2_regOut_1__1__1_), .B(s2_regOut_1__2__1_), 
        .Z(s2_chain_1__1__1_) );
  XOR2_X1 s2_compr_1_0_U1 ( .A(s2_regOut_1__1__0_), .B(s2_regOut_1__2__0_), 
        .Z(s2_chain_1__1__0_) );
  XOR2_X2 s2_compr_1_1_U4 ( .A(s2_chain_1__1__1_), .B(s2_regOut_1__3__1_), .Z(
        stage2Out[17]) );
  XOR2_X2 s2_compr_1_1_U3 ( .A(s2_chain_1__1__0_), .B(s2_regOut_1__3__0_), .Z(
        stage2Out[16]) );
  XOR2_X2 s2_compr_1_1_U2 ( .A(s2_chain_1__1__2_), .B(s2_regOut_1__3__2_), .Z(
        stage2Out[18]) );
  XOR2_X2 s2_compr_1_1_U1 ( .A(s2_chain_1__1__3_), .B(s2_regOut_1__3__3_), .Z(
        stage2Out[19]) );
  XOR2_X1 s2_compr_2_0_U4 ( .A(s2_regOut_2__1__3_), .B(s2_regOut_2__2__3_), 
        .Z(s2_chain_2__1__3_) );
  XOR2_X1 s2_compr_2_0_U3 ( .A(s2_regOut_2__1__2_), .B(s2_regOut_2__2__2_), 
        .Z(s2_chain_2__1__2_) );
  XOR2_X1 s2_compr_2_0_U2 ( .A(s2_regOut_2__1__1_), .B(s2_regOut_2__2__1_), 
        .Z(s2_chain_2__1__1_) );
  XOR2_X1 s2_compr_2_0_U1 ( .A(s2_regOut_2__1__0_), .B(s2_regOut_2__2__0_), 
        .Z(s2_chain_2__1__0_) );
  XOR2_X2 s2_compr_2_1_U4 ( .A(s2_chain_2__1__1_), .B(s2_regOut_2__3__1_), .Z(
        stage2Out[29]) );
  XOR2_X2 s2_compr_2_1_U3 ( .A(s2_chain_2__1__0_), .B(s2_regOut_2__3__0_), .Z(
        stage2Out[28]) );
  XOR2_X2 s2_compr_2_1_U2 ( .A(s2_chain_2__1__2_), .B(s2_regOut_2__3__2_), .Z(
        stage2Out[30]) );
  XOR2_X2 s2_compr_2_1_U1 ( .A(s2_chain_2__1__3_), .B(s2_regOut_2__3__3_), .Z(
        stage2Out[31]) );
  XNOR2_X1 s3_U50 ( .A(s3_n24), .B(s3_n23), .ZN(s3_refreshed[17]) );
  XNOR2_X1 s3_U49 ( .A(randomS3[1]), .B(randomS3[3]), .ZN(s3_n23) );
  XOR2_X1 s3_U48 ( .A(s3_gf2_mul_out_2__2__1_), .B(s3_scale_out[5]), .Z(s3_n24) );
  XNOR2_X1 s3_U47 ( .A(s3_n22), .B(s3_xorResult[11]), .ZN(s3_refreshed[15]) );
  XNOR2_X1 s3_U46 ( .A(randomS3[5]), .B(randomS3[3]), .ZN(s3_n22) );
  XNOR2_X1 s3_U45 ( .A(s3_n21), .B(s3_xorResult[10]), .ZN(s3_refreshed[14]) );
  XNOR2_X1 s3_U44 ( .A(randomS3[4]), .B(randomS3[2]), .ZN(s3_n21) );
  XNOR2_X1 s3_U43 ( .A(s3_n20), .B(s3_xorResult[9]), .ZN(s3_refreshed[13]) );
  XNOR2_X1 s3_U42 ( .A(randomS3[7]), .B(randomS3[5]), .ZN(s3_n20) );
  XNOR2_X1 s3_U41 ( .A(s3_n19), .B(s3_xorResult[8]), .ZN(s3_refreshed[12]) );
  XNOR2_X1 s3_U40 ( .A(randomS3[6]), .B(randomS3[4]), .ZN(s3_n19) );
  XNOR2_X1 s3_U39 ( .A(s3_n18), .B(s3_xorResult[7]), .ZN(s3_refreshed[11]) );
  XNOR2_X1 s3_U38 ( .A(randomS3[9]), .B(randomS3[7]), .ZN(s3_n18) );
  XNOR2_X1 s3_U37 ( .A(s3_n17), .B(s3_xorResult[6]), .ZN(s3_refreshed[10]) );
  XNOR2_X1 s3_U36 ( .A(randomS3[8]), .B(randomS3[6]), .ZN(s3_n17) );
  XNOR2_X1 s3_U35 ( .A(s3_n16), .B(s3_n15), .ZN(s3_refreshed[9]) );
  XNOR2_X1 s3_U34 ( .A(randomS3[11]), .B(randomS3[9]), .ZN(s3_n15) );
  XOR2_X1 s3_U33 ( .A(s3_gf2_mul_out_1__1__1_), .B(s3_scale_out[3]), .Z(s3_n16) );
  XNOR2_X1 s3_U32 ( .A(s3_n14), .B(s3_xorResult[5]), .ZN(s3_refreshed[7]) );
  XNOR2_X1 s3_U31 ( .A(randomS3[13]), .B(randomS3[11]), .ZN(s3_n14) );
  XNOR2_X1 s3_U30 ( .A(s3_n13), .B(s3_xorResult[4]), .ZN(s3_refreshed[6]) );
  XNOR2_X1 s3_U29 ( .A(randomS3[12]), .B(randomS3[10]), .ZN(s3_n13) );
  XNOR2_X1 s3_U28 ( .A(s3_n12), .B(s3_xorResult[3]), .ZN(s3_refreshed[5]) );
  XNOR2_X1 s3_U27 ( .A(randomS3[15]), .B(randomS3[13]), .ZN(s3_n12) );
  XNOR2_X1 s3_U26 ( .A(s3_n11), .B(s3_xorResult[2]), .ZN(s3_refreshed[4]) );
  XNOR2_X1 s3_U25 ( .A(randomS3[14]), .B(randomS3[12]), .ZN(s3_n11) );
  XNOR2_X1 s3_U24 ( .A(s3_n10), .B(s3_xorResult[1]), .ZN(s3_refreshed[3]) );
  XNOR2_X1 s3_U23 ( .A(randomS3[17]), .B(randomS3[15]), .ZN(s3_n10) );
  XNOR2_X1 s3_U22 ( .A(s3_n9), .B(s3_xorResult[0]), .ZN(s3_refreshed[2]) );
  XNOR2_X1 s3_U21 ( .A(randomS3[16]), .B(randomS3[14]), .ZN(s3_n9) );
  XNOR2_X1 s3_U20 ( .A(s3_n8), .B(s3_n7), .ZN(s3_refreshed[1]) );
  XNOR2_X1 s3_U19 ( .A(randomS3[1]), .B(randomS3[17]), .ZN(s3_n7) );
  XOR2_X1 s3_U18 ( .A(s3_gf2_mul_out_0__0__1_), .B(s3_scale_out[1]), .Z(s3_n8)
         );
  XOR2_X1 s3_U17 ( .A(stage2Out[28]), .B(stage2Out[30]), .Z(s3_scale_in[2]) );
  XNOR2_X1 s3_U16 ( .A(s3_n5), .B(s3_n6), .ZN(s3_refreshed[16]) );
  XNOR2_X1 s3_U15 ( .A(s3_gf2_mul_out_2__2__0_), .B(s3_scale_out[4]), .ZN(
        s3_n6) );
  XOR2_X1 s3_U14 ( .A(randomS3[2]), .B(randomS3[0]), .Z(s3_n5) );
  XOR2_X1 s3_U13 ( .A(stage2Out[16]), .B(stage2Out[18]), .Z(s3_scale_in[1]) );
  XNOR2_X1 s3_U12 ( .A(s3_n3), .B(s3_n4), .ZN(s3_refreshed[8]) );
  XNOR2_X1 s3_U11 ( .A(s3_gf2_mul_out_1__1__0_), .B(s3_scale_out[2]), .ZN(
        s3_n4) );
  XOR2_X1 s3_U10 ( .A(randomS3[8]), .B(randomS3[10]), .Z(s3_n3) );
  XOR2_X1 s3_U9 ( .A(stage2Out[4]), .B(stage2Out[6]), .Z(s3_scale_in[0]) );
  XNOR2_X1 s3_U8 ( .A(s3_n1), .B(s3_n2), .ZN(s3_refreshed[0]) );
  XNOR2_X1 s3_U7 ( .A(s3_gf2_mul_out_0__0__0_), .B(s3_scale_out[0]), .ZN(s3_n2) );
  XOR2_X1 s3_U6 ( .A(randomS3[16]), .B(randomS3[0]), .Z(s3_n1) );
  XOR2_X1 s3_U5 ( .A(stage2Out[31]), .B(stage2Out[29]), .Z(s3_scale_out[5]) );
  XOR2_X1 s3_U4 ( .A(stage2Out[19]), .B(stage2Out[17]), .Z(s3_scale_out[3]) );
  XOR2_X1 s3_U3 ( .A(stage2Out[7]), .B(stage2Out[5]), .Z(s3_scale_out[1]) );
  DFF_X1 s3_regOut_reg_0__0__0_ ( .D(stage2Out[0]), .CK(clk), .Q(stage3Out[0]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__0__1_ ( .D(stage2Out[1]), .CK(clk), .Q(stage3Out[1]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__1__0_ ( .D(stage2Out[2]), .CK(clk), .Q(stage3Out[2]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__1__1_ ( .D(stage2Out[3]), .CK(clk), .Q(stage3Out[3]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__2__0_ ( .D(stage2Out[4]), .CK(clk), .Q(stage3Out[4]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__2__1_ ( .D(stage2Out[5]), .CK(clk), .Q(stage3Out[5]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__3__0_ ( .D(s3_refreshed[0]), .CK(clk), .Q(
        s3_regOut_0__3__0_), .QN() );
  DFF_X1 s3_regOut_reg_0__3__1_ ( .D(s3_refreshed[1]), .CK(clk), .Q(
        s3_regOut_0__3__1_), .QN() );
  DFF_X1 s3_regOut_reg_0__4__0_ ( .D(s3_refreshed[2]), .CK(clk), .Q(
        s3_regOut_0__4__0_), .QN() );
  DFF_X1 s3_regOut_reg_0__4__1_ ( .D(s3_refreshed[3]), .CK(clk), .Q(
        s3_regOut_0__4__1_), .QN() );
  DFF_X1 s3_regOut_reg_0__5__0_ ( .D(s3_refreshed[4]), .CK(clk), .Q(
        s3_regOut_0__5__0_), .QN() );
  DFF_X1 s3_regOut_reg_0__5__1_ ( .D(s3_refreshed[5]), .CK(clk), .Q(
        s3_regOut_0__5__1_), .QN() );
  DFF_X1 s3_regOut_reg_0__6__0_ ( .D(stage2Out[6]), .CK(clk), .Q(stage3Out[6]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__6__1_ ( .D(stage2Out[7]), .CK(clk), .Q(stage3Out[7]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__7__0_ ( .D(stage2Out[8]), .CK(clk), .Q(stage3Out[8]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__7__1_ ( .D(stage2Out[9]), .CK(clk), .Q(stage3Out[9]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__8__0_ ( .D(stage2Out[10]), .CK(clk), .Q(
        stage3Out[10]), .QN() );
  DFF_X1 s3_regOut_reg_0__8__1_ ( .D(stage2Out[11]), .CK(clk), .Q(
        stage3Out[11]), .QN() );
  DFF_X1 s3_regOut_reg_1__0__0_ ( .D(stage2Out[12]), .CK(clk), .Q(
        stage3Out[12]), .QN() );
  DFF_X1 s3_regOut_reg_1__0__1_ ( .D(stage2Out[13]), .CK(clk), .Q(
        stage3Out[13]), .QN() );
  DFF_X1 s3_regOut_reg_1__1__0_ ( .D(stage2Out[14]), .CK(clk), .Q(
        stage3Out[14]), .QN() );
  DFF_X1 s3_regOut_reg_1__1__1_ ( .D(stage2Out[15]), .CK(clk), .Q(
        stage3Out[15]), .QN() );
  DFF_X1 s3_regOut_reg_1__2__0_ ( .D(stage2Out[16]), .CK(clk), .Q(
        stage3Out[16]), .QN() );
  DFF_X1 s3_regOut_reg_1__2__1_ ( .D(stage2Out[17]), .CK(clk), .Q(
        stage3Out[17]), .QN() );
  DFF_X1 s3_regOut_reg_1__3__0_ ( .D(s3_refreshed[6]), .CK(clk), .Q(
        s3_regOut_1__3__0_), .QN() );
  DFF_X1 s3_regOut_reg_1__3__1_ ( .D(s3_refreshed[7]), .CK(clk), .Q(
        s3_regOut_1__3__1_), .QN() );
  DFF_X1 s3_regOut_reg_1__4__0_ ( .D(s3_refreshed[8]), .CK(clk), .Q(
        s3_regOut_1__4__0_), .QN() );
  DFF_X1 s3_regOut_reg_1__4__1_ ( .D(s3_refreshed[9]), .CK(clk), .Q(
        s3_regOut_1__4__1_), .QN() );
  DFF_X1 s3_regOut_reg_1__5__0_ ( .D(s3_refreshed[10]), .CK(clk), .Q(
        s3_regOut_1__5__0_), .QN() );
  DFF_X1 s3_regOut_reg_1__5__1_ ( .D(s3_refreshed[11]), .CK(clk), .Q(
        s3_regOut_1__5__1_), .QN() );
  DFF_X1 s3_regOut_reg_1__6__0_ ( .D(stage2Out[18]), .CK(clk), .Q(
        stage3Out[18]), .QN() );
  DFF_X1 s3_regOut_reg_1__6__1_ ( .D(stage2Out[19]), .CK(clk), .Q(
        stage3Out[19]), .QN() );
  DFF_X1 s3_regOut_reg_1__7__0_ ( .D(stage2Out[20]), .CK(clk), .Q(
        stage3Out[20]), .QN() );
  DFF_X1 s3_regOut_reg_1__7__1_ ( .D(stage2Out[21]), .CK(clk), .Q(
        stage3Out[21]), .QN() );
  DFF_X1 s3_regOut_reg_1__8__0_ ( .D(stage2Out[22]), .CK(clk), .Q(
        stage3Out[22]), .QN() );
  DFF_X1 s3_regOut_reg_1__8__1_ ( .D(stage2Out[23]), .CK(clk), .Q(
        stage3Out[23]), .QN() );
  DFF_X1 s3_regOut_reg_2__0__0_ ( .D(stage2Out[24]), .CK(clk), .Q(
        stage3Out[24]), .QN() );
  DFF_X1 s3_regOut_reg_2__0__1_ ( .D(stage2Out[25]), .CK(clk), .Q(
        stage3Out[25]), .QN() );
  DFF_X1 s3_regOut_reg_2__1__0_ ( .D(stage2Out[26]), .CK(clk), .Q(
        stage3Out[26]), .QN() );
  DFF_X1 s3_regOut_reg_2__1__1_ ( .D(stage2Out[27]), .CK(clk), .Q(
        stage3Out[27]), .QN() );
  DFF_X1 s3_regOut_reg_2__2__0_ ( .D(stage2Out[28]), .CK(clk), .Q(
        stage3Out[28]), .QN() );
  DFF_X1 s3_regOut_reg_2__2__1_ ( .D(stage2Out[29]), .CK(clk), .Q(
        stage3Out[29]), .QN() );
  DFF_X1 s3_regOut_reg_2__3__0_ ( .D(s3_refreshed[12]), .CK(clk), .Q(
        s3_regOut_2__3__0_), .QN() );
  DFF_X1 s3_regOut_reg_2__3__1_ ( .D(s3_refreshed[13]), .CK(clk), .Q(
        s3_regOut_2__3__1_), .QN() );
  DFF_X1 s3_regOut_reg_2__4__0_ ( .D(s3_refreshed[14]), .CK(clk), .Q(
        s3_regOut_2__4__0_), .QN() );
  DFF_X1 s3_regOut_reg_2__4__1_ ( .D(s3_refreshed[15]), .CK(clk), .Q(
        s3_regOut_2__4__1_), .QN() );
  DFF_X1 s3_regOut_reg_2__5__0_ ( .D(s3_refreshed[16]), .CK(clk), .Q(
        s3_regOut_2__5__0_), .QN() );
  DFF_X1 s3_regOut_reg_2__5__1_ ( .D(s3_refreshed[17]), .CK(clk), .Q(
        s3_regOut_2__5__1_), .QN() );
  DFF_X1 s3_regOut_reg_2__6__0_ ( .D(stage2Out[30]), .CK(clk), .Q(
        stage3Out[30]), .QN() );
  DFF_X1 s3_regOut_reg_2__6__1_ ( .D(stage2Out[31]), .CK(clk), .Q(
        stage3Out[31]), .QN() );
  DFF_X1 s3_regOut_reg_2__7__0_ ( .D(stage2Out[32]), .CK(clk), .Q(
        stage3Out[32]), .QN() );
  DFF_X1 s3_regOut_reg_2__7__1_ ( .D(stage2Out[33]), .CK(clk), .Q(
        stage3Out[33]), .QN() );
  DFF_X1 s3_regOut_reg_2__8__0_ ( .D(stage2Out[34]), .CK(clk), .Q(
        stage3Out[34]), .QN() );
  DFF_X1 s3_regOut_reg_2__8__1_ ( .D(stage2Out[35]), .CK(clk), .Q(
        stage3Out[35]), .QN() );
  XOR2_X1 s3_sqsc_2_U1 ( .A(s3_scale_in[2]), .B(s3_scale_out[5]), .Z(
        s3_scale_out[4]) );
  XOR2_X1 s3_sqsc_1_U1 ( .A(s3_scale_in[1]), .B(s3_scale_out[3]), .Z(
        s3_scale_out[2]) );
  XOR2_X1 s3_sqsc_0_U1 ( .A(s3_scale_in[0]), .B(s3_scale_out[1]), .Z(
        s3_scale_out[0]) );
  XNOR2_X1 s3_mul1_2_2_U6 ( .A(s3_mul1_2_2_n14), .B(s3_mul1_2_2_n13), .ZN(
        s3_gf2_mul_out_2__2__1_) );
  NAND2_X1 s3_mul1_2_2_U5 ( .A1(stage2Out[31]), .A2(stage2Out[29]), .ZN(
        s3_mul1_2_2_n14) );
  OAI22_X1 s3_mul1_2_2_U4 ( .A1(stage2Out[28]), .A2(stage2Out[29]), .B1(
        stage2Out[30]), .B2(stage2Out[31]), .ZN(s3_mul1_2_2_n12) );
  AOI221_X1 s3_mul1_2_2_U3 ( .B1(stage2Out[28]), .B2(stage2Out[29]), .C1(
        stage2Out[31]), .C2(stage2Out[30]), .A(s3_mul1_2_2_n12), .ZN(
        s3_mul1_2_2_n13) );
  XNOR2_X1 s3_mul1_2_2_U2 ( .A(s3_mul1_2_2_n11), .B(s3_mul1_2_2_n13), .ZN(
        s3_gf2_mul_out_2__2__0_) );
  NAND2_X1 s3_mul1_2_2_U1 ( .A1(stage2Out[30]), .A2(stage2Out[28]), .ZN(
        s3_mul1_2_2_n11) );
  XNOR2_X1 s3_mul1_2_1_U6 ( .A(s3_mul1_2_1_n14), .B(s3_mul1_2_1_n13), .ZN(
        s3_xorResult[11]) );
  NAND2_X1 s3_mul1_2_1_U5 ( .A1(stage2Out[31]), .A2(stage2Out[17]), .ZN(
        s3_mul1_2_1_n14) );
  XNOR2_X1 s3_mul1_2_1_U4 ( .A(s3_mul1_2_1_n13), .B(s3_mul1_2_1_n12), .ZN(
        s3_xorResult[10]) );
  NAND2_X1 s3_mul1_2_1_U3 ( .A1(stage2Out[16]), .A2(stage2Out[30]), .ZN(
        s3_mul1_2_1_n12) );
  AOI221_X1 s3_mul1_2_1_U2 ( .B1(stage2Out[16]), .B2(stage2Out[17]), .C1(
        stage2Out[31]), .C2(stage2Out[30]), .A(s3_mul1_2_1_n11), .ZN(
        s3_mul1_2_1_n13) );
  OAI22_X1 s3_mul1_2_1_U1 ( .A1(stage2Out[16]), .A2(stage2Out[17]), .B1(
        stage2Out[30]), .B2(stage2Out[31]), .ZN(s3_mul1_2_1_n11) );
  XNOR2_X1 s3_mul1_2_0_U6 ( .A(s3_mul1_2_0_n14), .B(s3_mul1_2_0_n13), .ZN(
        s3_xorResult[9]) );
  NAND2_X1 s3_mul1_2_0_U5 ( .A1(stage2Out[31]), .A2(stage2Out[5]), .ZN(
        s3_mul1_2_0_n14) );
  XNOR2_X1 s3_mul1_2_0_U4 ( .A(s3_mul1_2_0_n13), .B(s3_mul1_2_0_n12), .ZN(
        s3_xorResult[8]) );
  NAND2_X1 s3_mul1_2_0_U3 ( .A1(stage2Out[4]), .A2(stage2Out[30]), .ZN(
        s3_mul1_2_0_n12) );
  AOI221_X1 s3_mul1_2_0_U2 ( .B1(stage2Out[4]), .B2(stage2Out[5]), .C1(
        stage2Out[31]), .C2(stage2Out[30]), .A(s3_mul1_2_0_n11), .ZN(
        s3_mul1_2_0_n13) );
  OAI22_X1 s3_mul1_2_0_U1 ( .A1(stage2Out[4]), .A2(stage2Out[5]), .B1(
        stage2Out[30]), .B2(stage2Out[31]), .ZN(s3_mul1_2_0_n11) );
  XNOR2_X1 s3_mul1_1_2_U6 ( .A(s3_mul1_1_2_n14), .B(s3_mul1_1_2_n13), .ZN(
        s3_xorResult[7]) );
  NAND2_X1 s3_mul1_1_2_U5 ( .A1(stage2Out[19]), .A2(stage2Out[29]), .ZN(
        s3_mul1_1_2_n14) );
  XNOR2_X1 s3_mul1_1_2_U4 ( .A(s3_mul1_1_2_n13), .B(s3_mul1_1_2_n12), .ZN(
        s3_xorResult[6]) );
  NAND2_X1 s3_mul1_1_2_U3 ( .A1(stage2Out[28]), .A2(stage2Out[18]), .ZN(
        s3_mul1_1_2_n12) );
  AOI221_X1 s3_mul1_1_2_U2 ( .B1(stage2Out[28]), .B2(stage2Out[29]), .C1(
        stage2Out[19]), .C2(stage2Out[18]), .A(s3_mul1_1_2_n11), .ZN(
        s3_mul1_1_2_n13) );
  OAI22_X1 s3_mul1_1_2_U1 ( .A1(stage2Out[28]), .A2(stage2Out[29]), .B1(
        stage2Out[18]), .B2(stage2Out[19]), .ZN(s3_mul1_1_2_n11) );
  XNOR2_X1 s3_mul1_1_1_U6 ( .A(s3_mul1_1_1_n14), .B(s3_mul1_1_1_n13), .ZN(
        s3_gf2_mul_out_1__1__1_) );
  NAND2_X1 s3_mul1_1_1_U5 ( .A1(stage2Out[19]), .A2(stage2Out[17]), .ZN(
        s3_mul1_1_1_n14) );
  OAI22_X1 s3_mul1_1_1_U4 ( .A1(stage2Out[16]), .A2(stage2Out[17]), .B1(
        stage2Out[18]), .B2(stage2Out[19]), .ZN(s3_mul1_1_1_n12) );
  AOI221_X1 s3_mul1_1_1_U3 ( .B1(stage2Out[16]), .B2(stage2Out[17]), .C1(
        stage2Out[19]), .C2(stage2Out[18]), .A(s3_mul1_1_1_n12), .ZN(
        s3_mul1_1_1_n13) );
  XNOR2_X1 s3_mul1_1_1_U2 ( .A(s3_mul1_1_1_n11), .B(s3_mul1_1_1_n13), .ZN(
        s3_gf2_mul_out_1__1__0_) );
  NAND2_X1 s3_mul1_1_1_U1 ( .A1(stage2Out[18]), .A2(stage2Out[16]), .ZN(
        s3_mul1_1_1_n11) );
  XNOR2_X1 s3_mul1_1_0_U6 ( .A(s3_mul1_1_0_n14), .B(s3_mul1_1_0_n13), .ZN(
        s3_xorResult[5]) );
  NAND2_X1 s3_mul1_1_0_U5 ( .A1(stage2Out[19]), .A2(stage2Out[5]), .ZN(
        s3_mul1_1_0_n14) );
  XNOR2_X1 s3_mul1_1_0_U4 ( .A(s3_mul1_1_0_n13), .B(s3_mul1_1_0_n12), .ZN(
        s3_xorResult[4]) );
  NAND2_X1 s3_mul1_1_0_U3 ( .A1(stage2Out[4]), .A2(stage2Out[18]), .ZN(
        s3_mul1_1_0_n12) );
  AOI221_X1 s3_mul1_1_0_U2 ( .B1(stage2Out[4]), .B2(stage2Out[5]), .C1(
        stage2Out[19]), .C2(stage2Out[18]), .A(s3_mul1_1_0_n11), .ZN(
        s3_mul1_1_0_n13) );
  OAI22_X1 s3_mul1_1_0_U1 ( .A1(stage2Out[4]), .A2(stage2Out[5]), .B1(
        stage2Out[18]), .B2(stage2Out[19]), .ZN(s3_mul1_1_0_n11) );
  XNOR2_X1 s3_mul1_0_2_U6 ( .A(s3_mul1_0_2_n14), .B(s3_mul1_0_2_n13), .ZN(
        s3_xorResult[3]) );
  NAND2_X1 s3_mul1_0_2_U5 ( .A1(stage2Out[7]), .A2(stage2Out[29]), .ZN(
        s3_mul1_0_2_n14) );
  XNOR2_X1 s3_mul1_0_2_U4 ( .A(s3_mul1_0_2_n13), .B(s3_mul1_0_2_n12), .ZN(
        s3_xorResult[2]) );
  NAND2_X1 s3_mul1_0_2_U3 ( .A1(stage2Out[28]), .A2(stage2Out[6]), .ZN(
        s3_mul1_0_2_n12) );
  AOI221_X1 s3_mul1_0_2_U2 ( .B1(stage2Out[28]), .B2(stage2Out[29]), .C1(
        stage2Out[7]), .C2(stage2Out[6]), .A(s3_mul1_0_2_n11), .ZN(
        s3_mul1_0_2_n13) );
  OAI22_X1 s3_mul1_0_2_U1 ( .A1(stage2Out[28]), .A2(stage2Out[29]), .B1(
        stage2Out[6]), .B2(stage2Out[7]), .ZN(s3_mul1_0_2_n11) );
  XNOR2_X1 s3_mul1_0_1_U6 ( .A(s3_mul1_0_1_n14), .B(s3_mul1_0_1_n13), .ZN(
        s3_xorResult[1]) );
  NAND2_X1 s3_mul1_0_1_U5 ( .A1(stage2Out[7]), .A2(stage2Out[17]), .ZN(
        s3_mul1_0_1_n14) );
  XNOR2_X1 s3_mul1_0_1_U4 ( .A(s3_mul1_0_1_n13), .B(s3_mul1_0_1_n12), .ZN(
        s3_xorResult[0]) );
  NAND2_X1 s3_mul1_0_1_U3 ( .A1(stage2Out[16]), .A2(stage2Out[6]), .ZN(
        s3_mul1_0_1_n12) );
  AOI221_X1 s3_mul1_0_1_U2 ( .B1(stage2Out[16]), .B2(stage2Out[17]), .C1(
        stage2Out[7]), .C2(stage2Out[6]), .A(s3_mul1_0_1_n11), .ZN(
        s3_mul1_0_1_n13) );
  OAI22_X1 s3_mul1_0_1_U1 ( .A1(stage2Out[16]), .A2(stage2Out[17]), .B1(
        stage2Out[6]), .B2(stage2Out[7]), .ZN(s3_mul1_0_1_n11) );
  XNOR2_X1 s3_mul1_0_0_U6 ( .A(s3_mul1_0_0_n14), .B(s3_mul1_0_0_n13), .ZN(
        s3_gf2_mul_out_0__0__1_) );
  NAND2_X1 s3_mul1_0_0_U5 ( .A1(stage2Out[7]), .A2(stage2Out[5]), .ZN(
        s3_mul1_0_0_n14) );
  OAI22_X1 s3_mul1_0_0_U4 ( .A1(stage2Out[4]), .A2(stage2Out[5]), .B1(
        stage2Out[6]), .B2(stage2Out[7]), .ZN(s3_mul1_0_0_n12) );
  AOI221_X1 s3_mul1_0_0_U3 ( .B1(stage2Out[4]), .B2(stage2Out[5]), .C1(
        stage2Out[7]), .C2(stage2Out[6]), .A(s3_mul1_0_0_n12), .ZN(
        s3_mul1_0_0_n13) );
  XNOR2_X1 s3_mul1_0_0_U2 ( .A(s3_mul1_0_0_n11), .B(s3_mul1_0_0_n13), .ZN(
        s3_gf2_mul_out_0__0__0_) );
  NAND2_X1 s3_mul1_0_0_U1 ( .A1(stage2Out[6]), .A2(stage2Out[4]), .ZN(
        s3_mul1_0_0_n11) );
  XOR2_X1 s3_compr_0_0_U2 ( .A(s3_regOut_0__3__1_), .B(s3_regOut_0__4__1_), 
        .Z(s3_chain_0__1__1_) );
  XOR2_X1 s3_compr_0_0_U1 ( .A(s3_regOut_0__3__0_), .B(s3_regOut_0__4__0_), 
        .Z(s3_chain_0__1__0_) );
  XOR2_X2 s3_compr_0_1_U2 ( .A(s3_chain_0__1__0_), .B(s3_regOut_0__5__0_), .Z(
        s4_inv_out_0__1_) );
  XOR2_X2 s3_compr_0_1_U1 ( .A(s3_chain_0__1__1_), .B(s3_regOut_0__5__1_), .Z(
        s4_inv_out_0__0_) );
  XOR2_X1 s3_compr_1_0_U2 ( .A(s3_regOut_1__3__1_), .B(s3_regOut_1__4__1_), 
        .Z(s3_chain_1__1__1_) );
  XOR2_X1 s3_compr_1_0_U1 ( .A(s3_regOut_1__3__0_), .B(s3_regOut_1__4__0_), 
        .Z(s3_chain_1__1__0_) );
  XOR2_X2 s3_compr_1_1_U2 ( .A(s3_chain_1__1__0_), .B(s3_regOut_1__5__0_), .Z(
        s4_inv_out_1__1_) );
  XOR2_X2 s3_compr_1_1_U1 ( .A(s3_chain_1__1__1_), .B(s3_regOut_1__5__1_), .Z(
        s4_inv_out_1__0_) );
  XOR2_X1 s3_compr_2_0_U2 ( .A(s3_regOut_2__3__1_), .B(s3_regOut_2__4__1_), 
        .Z(s3_chain_2__1__1_) );
  XOR2_X1 s3_compr_2_0_U1 ( .A(s3_regOut_2__3__0_), .B(s3_regOut_2__4__0_), 
        .Z(s3_chain_2__1__0_) );
  XOR2_X2 s3_compr_2_1_U2 ( .A(s3_chain_2__1__0_), .B(s3_regOut_2__5__0_), .Z(
        s4_inv_out_2__1_) );
  XOR2_X2 s3_compr_2_1_U1 ( .A(s3_chain_2__1__1_), .B(s3_regOut_2__5__1_), .Z(
        s4_inv_out_2__0_) );
  XNOR2_X1 s4_U74 ( .A(s4_n36), .B(s4_concat[35]), .ZN(s4_refreshed[35]) );
  XNOR2_X1 s4_U73 ( .A(randomS4[3]), .B(randomS4[7]), .ZN(s4_n36) );
  XNOR2_X1 s4_U72 ( .A(s4_n35), .B(s4_concat[34]), .ZN(s4_refreshed[34]) );
  XNOR2_X1 s4_U71 ( .A(randomS4[2]), .B(randomS4[6]), .ZN(s4_n35) );
  XNOR2_X1 s4_U70 ( .A(s4_n34), .B(s4_concat[33]), .ZN(s4_refreshed[33]) );
  XNOR2_X1 s4_U69 ( .A(randomS4[1]), .B(randomS4[5]), .ZN(s4_n34) );
  XNOR2_X1 s4_U68 ( .A(s4_n33), .B(s4_concat[32]), .ZN(s4_refreshed[32]) );
  XNOR2_X1 s4_U67 ( .A(randomS4[0]), .B(randomS4[4]), .ZN(s4_n33) );
  XNOR2_X1 s4_U66 ( .A(s4_n32), .B(s4_concat[31]), .ZN(s4_refreshed[31]) );
  XNOR2_X1 s4_U65 ( .A(randomS4[11]), .B(randomS4[7]), .ZN(s4_n32) );
  XNOR2_X1 s4_U64 ( .A(s4_n31), .B(s4_concat[30]), .ZN(s4_refreshed[30]) );
  XNOR2_X1 s4_U63 ( .A(randomS4[10]), .B(randomS4[6]), .ZN(s4_n31) );
  XNOR2_X1 s4_U62 ( .A(s4_n30), .B(s4_concat[29]), .ZN(s4_refreshed[29]) );
  XNOR2_X1 s4_U61 ( .A(randomS4[9]), .B(randomS4[5]), .ZN(s4_n30) );
  XNOR2_X1 s4_U60 ( .A(s4_n29), .B(s4_concat[28]), .ZN(s4_refreshed[28]) );
  XNOR2_X1 s4_U59 ( .A(randomS4[8]), .B(randomS4[4]), .ZN(s4_n29) );
  XNOR2_X1 s4_U58 ( .A(s4_n28), .B(s4_concat[27]), .ZN(s4_refreshed[27]) );
  XNOR2_X1 s4_U57 ( .A(randomS4[15]), .B(randomS4[11]), .ZN(s4_n28) );
  XNOR2_X1 s4_U56 ( .A(s4_n27), .B(s4_concat[26]), .ZN(s4_refreshed[26]) );
  XNOR2_X1 s4_U55 ( .A(randomS4[14]), .B(randomS4[10]), .ZN(s4_n27) );
  XNOR2_X1 s4_U54 ( .A(s4_n26), .B(s4_concat[25]), .ZN(s4_refreshed[25]) );
  XNOR2_X1 s4_U53 ( .A(randomS4[13]), .B(randomS4[9]), .ZN(s4_n26) );
  XNOR2_X1 s4_U52 ( .A(s4_n25), .B(s4_concat[24]), .ZN(s4_refreshed[24]) );
  XNOR2_X1 s4_U51 ( .A(randomS4[12]), .B(randomS4[8]), .ZN(s4_n25) );
  XNOR2_X1 s4_U50 ( .A(s4_n24), .B(s4_concat[23]), .ZN(s4_refreshed[23]) );
  XNOR2_X1 s4_U49 ( .A(randomS4[19]), .B(randomS4[15]), .ZN(s4_n24) );
  XNOR2_X1 s4_U48 ( .A(s4_n23), .B(s4_concat[22]), .ZN(s4_refreshed[22]) );
  XNOR2_X1 s4_U47 ( .A(randomS4[18]), .B(randomS4[14]), .ZN(s4_n23) );
  XNOR2_X1 s4_U46 ( .A(s4_n22), .B(s4_concat[21]), .ZN(s4_refreshed[21]) );
  XNOR2_X1 s4_U45 ( .A(randomS4[17]), .B(randomS4[13]), .ZN(s4_n22) );
  XNOR2_X1 s4_U44 ( .A(s4_n21), .B(s4_concat[20]), .ZN(s4_refreshed[20]) );
  XNOR2_X1 s4_U43 ( .A(randomS4[16]), .B(randomS4[12]), .ZN(s4_n21) );
  XNOR2_X1 s4_U42 ( .A(s4_n20), .B(s4_concat[19]), .ZN(s4_refreshed[19]) );
  XNOR2_X1 s4_U41 ( .A(randomS4[23]), .B(randomS4[19]), .ZN(s4_n20) );
  XNOR2_X1 s4_U40 ( .A(s4_n19), .B(s4_concat[18]), .ZN(s4_refreshed[18]) );
  XNOR2_X1 s4_U39 ( .A(randomS4[22]), .B(randomS4[18]), .ZN(s4_n19) );
  XNOR2_X1 s4_U38 ( .A(s4_n18), .B(s4_concat[17]), .ZN(s4_refreshed[17]) );
  XNOR2_X1 s4_U37 ( .A(randomS4[21]), .B(randomS4[17]), .ZN(s4_n18) );
  XNOR2_X1 s4_U36 ( .A(s4_n17), .B(s4_concat[16]), .ZN(s4_refreshed[16]) );
  XNOR2_X1 s4_U35 ( .A(randomS4[20]), .B(randomS4[16]), .ZN(s4_n17) );
  XNOR2_X1 s4_U34 ( .A(s4_n16), .B(s4_concat[15]), .ZN(s4_refreshed[15]) );
  XNOR2_X1 s4_U33 ( .A(randomS4[27]), .B(randomS4[23]), .ZN(s4_n16) );
  XNOR2_X1 s4_U32 ( .A(s4_n15), .B(s4_concat[14]), .ZN(s4_refreshed[14]) );
  XNOR2_X1 s4_U31 ( .A(randomS4[26]), .B(randomS4[22]), .ZN(s4_n15) );
  XNOR2_X1 s4_U30 ( .A(s4_n14), .B(s4_concat[13]), .ZN(s4_refreshed[13]) );
  XNOR2_X1 s4_U29 ( .A(randomS4[25]), .B(randomS4[21]), .ZN(s4_n14) );
  XNOR2_X1 s4_U28 ( .A(s4_n13), .B(s4_concat[12]), .ZN(s4_refreshed[12]) );
  XNOR2_X1 s4_U27 ( .A(randomS4[24]), .B(randomS4[20]), .ZN(s4_n13) );
  XNOR2_X1 s4_U26 ( .A(s4_n12), .B(s4_concat[11]), .ZN(s4_refreshed[11]) );
  XNOR2_X1 s4_U25 ( .A(randomS4[31]), .B(randomS4[27]), .ZN(s4_n12) );
  XNOR2_X1 s4_U24 ( .A(s4_n11), .B(s4_concat[10]), .ZN(s4_refreshed[10]) );
  XNOR2_X1 s4_U23 ( .A(randomS4[30]), .B(randomS4[26]), .ZN(s4_n11) );
  XNOR2_X1 s4_U22 ( .A(s4_n10), .B(s4_concat[9]), .ZN(s4_refreshed[9]) );
  XNOR2_X1 s4_U21 ( .A(randomS4[29]), .B(randomS4[25]), .ZN(s4_n10) );
  XNOR2_X1 s4_U20 ( .A(s4_n9), .B(s4_concat[8]), .ZN(s4_refreshed[8]) );
  XNOR2_X1 s4_U19 ( .A(randomS4[28]), .B(randomS4[24]), .ZN(s4_n9) );
  XNOR2_X1 s4_U18 ( .A(s4_n8), .B(s4_concat[7]), .ZN(s4_refreshed[7]) );
  XNOR2_X1 s4_U17 ( .A(randomS4[35]), .B(randomS4[31]), .ZN(s4_n8) );
  XNOR2_X1 s4_U16 ( .A(s4_n7), .B(s4_concat[6]), .ZN(s4_refreshed[6]) );
  XNOR2_X1 s4_U15 ( .A(randomS4[34]), .B(randomS4[30]), .ZN(s4_n7) );
  XNOR2_X1 s4_U14 ( .A(s4_n6), .B(s4_concat[5]), .ZN(s4_refreshed[5]) );
  XNOR2_X1 s4_U13 ( .A(randomS4[33]), .B(randomS4[29]), .ZN(s4_n6) );
  XNOR2_X1 s4_U12 ( .A(s4_n5), .B(s4_concat[4]), .ZN(s4_refreshed[4]) );
  XNOR2_X1 s4_U11 ( .A(randomS4[32]), .B(randomS4[28]), .ZN(s4_n5) );
  XNOR2_X1 s4_U10 ( .A(s4_n4), .B(s4_concat[3]), .ZN(s4_refreshed[3]) );
  XNOR2_X1 s4_U9 ( .A(randomS4[3]), .B(randomS4[35]), .ZN(s4_n4) );
  XNOR2_X1 s4_U8 ( .A(s4_n3), .B(s4_concat[2]), .ZN(s4_refreshed[2]) );
  XNOR2_X1 s4_U7 ( .A(randomS4[2]), .B(randomS4[34]), .ZN(s4_n3) );
  XNOR2_X1 s4_U6 ( .A(s4_n2), .B(s4_concat[1]), .ZN(s4_refreshed[1]) );
  XNOR2_X1 s4_U5 ( .A(randomS4[1]), .B(randomS4[33]), .ZN(s4_n2) );
  XNOR2_X1 s4_U4 ( .A(s4_n1), .B(s4_concat[0]), .ZN(s4_refreshed[0]) );
  XNOR2_X1 s4_U3 ( .A(randomS4[0]), .B(randomS4[32]), .ZN(s4_n1) );
  DFF_X1 s4_regOut_reg_0__0__0_ ( .D(stage3Out[0]), .CK(clk), .Q(stage4Out[0]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__0__1_ ( .D(stage3Out[1]), .CK(clk), .Q(stage4Out[1]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__0__2_ ( .D(stage3Out[2]), .CK(clk), .Q(stage4Out[2]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__0__3_ ( .D(stage3Out[3]), .CK(clk), .Q(stage4Out[3]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__1__0_ ( .D(s4_refreshed[0]), .CK(clk), .Q(
        s4_regOut_0__1__0_), .QN() );
  DFF_X1 s4_regOut_reg_0__1__1_ ( .D(s4_refreshed[1]), .CK(clk), .Q(
        s4_regOut_0__1__1_), .QN() );
  DFF_X1 s4_regOut_reg_0__1__2_ ( .D(s4_refreshed[2]), .CK(clk), .Q(
        s4_regOut_0__1__2_), .QN() );
  DFF_X1 s4_regOut_reg_0__1__3_ ( .D(s4_refreshed[3]), .CK(clk), .Q(
        s4_regOut_0__1__3_), .QN() );
  DFF_X1 s4_regOut_reg_0__2__0_ ( .D(s4_refreshed[4]), .CK(clk), .Q(
        s4_regOut_0__2__0_), .QN() );
  DFF_X1 s4_regOut_reg_0__2__1_ ( .D(s4_refreshed[5]), .CK(clk), .Q(
        s4_regOut_0__2__1_), .QN() );
  DFF_X1 s4_regOut_reg_0__2__2_ ( .D(s4_refreshed[6]), .CK(clk), .Q(
        s4_regOut_0__2__2_), .QN() );
  DFF_X1 s4_regOut_reg_0__2__3_ ( .D(s4_refreshed[7]), .CK(clk), .Q(
        s4_regOut_0__2__3_), .QN() );
  DFF_X1 s4_regOut_reg_0__3__0_ ( .D(s4_refreshed[8]), .CK(clk), .Q(
        s4_regOut_0__3__0_), .QN() );
  DFF_X1 s4_regOut_reg_0__3__1_ ( .D(s4_refreshed[9]), .CK(clk), .Q(
        s4_regOut_0__3__1_), .QN() );
  DFF_X1 s4_regOut_reg_0__3__2_ ( .D(s4_refreshed[10]), .CK(clk), .Q(
        s4_regOut_0__3__2_), .QN() );
  DFF_X1 s4_regOut_reg_0__3__3_ ( .D(s4_refreshed[11]), .CK(clk), .Q(
        s4_regOut_0__3__3_), .QN() );
  DFF_X1 s4_regOut_reg_0__4__0_ ( .D(stage3Out[8]), .CK(clk), .Q(stage4Out[8]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__4__1_ ( .D(stage3Out[9]), .CK(clk), .Q(stage4Out[9]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__4__2_ ( .D(stage3Out[10]), .CK(clk), .Q(
        stage4Out[10]), .QN() );
  DFF_X1 s4_regOut_reg_0__4__3_ ( .D(stage3Out[11]), .CK(clk), .Q(
        stage4Out[11]), .QN() );
  DFF_X1 s4_regOut_reg_1__0__0_ ( .D(stage3Out[12]), .CK(clk), .Q(
        stage4Out[12]), .QN() );
  DFF_X1 s4_regOut_reg_1__0__1_ ( .D(stage3Out[13]), .CK(clk), .Q(
        stage4Out[13]), .QN() );
  DFF_X1 s4_regOut_reg_1__0__2_ ( .D(stage3Out[14]), .CK(clk), .Q(
        stage4Out[14]), .QN() );
  DFF_X1 s4_regOut_reg_1__0__3_ ( .D(stage3Out[15]), .CK(clk), .Q(
        stage4Out[15]), .QN() );
  DFF_X1 s4_regOut_reg_1__1__0_ ( .D(s4_refreshed[12]), .CK(clk), .Q(
        s4_regOut_1__1__0_), .QN() );
  DFF_X1 s4_regOut_reg_1__1__1_ ( .D(s4_refreshed[13]), .CK(clk), .Q(
        s4_regOut_1__1__1_), .QN() );
  DFF_X1 s4_regOut_reg_1__1__2_ ( .D(s4_refreshed[14]), .CK(clk), .Q(
        s4_regOut_1__1__2_), .QN() );
  DFF_X1 s4_regOut_reg_1__1__3_ ( .D(s4_refreshed[15]), .CK(clk), .Q(
        s4_regOut_1__1__3_), .QN() );
  DFF_X1 s4_regOut_reg_1__2__0_ ( .D(s4_refreshed[16]), .CK(clk), .Q(
        s4_regOut_1__2__0_), .QN() );
  DFF_X1 s4_regOut_reg_1__2__1_ ( .D(s4_refreshed[17]), .CK(clk), .Q(
        s4_regOut_1__2__1_), .QN() );
  DFF_X1 s4_regOut_reg_1__2__2_ ( .D(s4_refreshed[18]), .CK(clk), .Q(
        s4_regOut_1__2__2_), .QN() );
  DFF_X1 s4_regOut_reg_1__2__3_ ( .D(s4_refreshed[19]), .CK(clk), .Q(
        s4_regOut_1__2__3_), .QN() );
  DFF_X1 s4_regOut_reg_1__3__0_ ( .D(s4_refreshed[20]), .CK(clk), .Q(
        s4_regOut_1__3__0_), .QN() );
  DFF_X1 s4_regOut_reg_1__3__1_ ( .D(s4_refreshed[21]), .CK(clk), .Q(
        s4_regOut_1__3__1_), .QN() );
  DFF_X1 s4_regOut_reg_1__3__2_ ( .D(s4_refreshed[22]), .CK(clk), .Q(
        s4_regOut_1__3__2_), .QN() );
  DFF_X1 s4_regOut_reg_1__3__3_ ( .D(s4_refreshed[23]), .CK(clk), .Q(
        s4_regOut_1__3__3_), .QN() );
  DFF_X1 s4_regOut_reg_1__4__0_ ( .D(stage3Out[20]), .CK(clk), .Q(
        stage4Out[20]), .QN() );
  DFF_X1 s4_regOut_reg_1__4__1_ ( .D(stage3Out[21]), .CK(clk), .Q(
        stage4Out[21]), .QN() );
  DFF_X1 s4_regOut_reg_1__4__2_ ( .D(stage3Out[22]), .CK(clk), .Q(
        stage4Out[22]), .QN() );
  DFF_X1 s4_regOut_reg_1__4__3_ ( .D(stage3Out[23]), .CK(clk), .Q(
        stage4Out[23]), .QN() );
  DFF_X1 s4_regOut_reg_2__0__0_ ( .D(stage3Out[24]), .CK(clk), .Q(
        stage4Out[24]), .QN() );
  DFF_X1 s4_regOut_reg_2__0__1_ ( .D(stage3Out[25]), .CK(clk), .Q(
        stage4Out[25]), .QN() );
  DFF_X1 s4_regOut_reg_2__0__2_ ( .D(stage3Out[26]), .CK(clk), .Q(
        stage4Out[26]), .QN() );
  DFF_X1 s4_regOut_reg_2__0__3_ ( .D(stage3Out[27]), .CK(clk), .Q(
        stage4Out[27]), .QN() );
  DFF_X1 s4_regOut_reg_2__1__0_ ( .D(s4_refreshed[24]), .CK(clk), .Q(
        s4_regOut_2__1__0_), .QN() );
  DFF_X1 s4_regOut_reg_2__1__1_ ( .D(s4_refreshed[25]), .CK(clk), .Q(
        s4_regOut_2__1__1_), .QN() );
  DFF_X1 s4_regOut_reg_2__1__2_ ( .D(s4_refreshed[26]), .CK(clk), .Q(
        s4_regOut_2__1__2_), .QN() );
  DFF_X1 s4_regOut_reg_2__1__3_ ( .D(s4_refreshed[27]), .CK(clk), .Q(
        s4_regOut_2__1__3_), .QN() );
  DFF_X1 s4_regOut_reg_2__2__0_ ( .D(s4_refreshed[28]), .CK(clk), .Q(
        s4_regOut_2__2__0_), .QN() );
  DFF_X1 s4_regOut_reg_2__2__1_ ( .D(s4_refreshed[29]), .CK(clk), .Q(
        s4_regOut_2__2__1_), .QN() );
  DFF_X1 s4_regOut_reg_2__2__2_ ( .D(s4_refreshed[30]), .CK(clk), .Q(
        s4_regOut_2__2__2_), .QN() );
  DFF_X1 s4_regOut_reg_2__2__3_ ( .D(s4_refreshed[31]), .CK(clk), .Q(
        s4_regOut_2__2__3_), .QN() );
  DFF_X1 s4_regOut_reg_2__3__0_ ( .D(s4_refreshed[32]), .CK(clk), .Q(
        s4_regOut_2__3__0_), .QN() );
  DFF_X1 s4_regOut_reg_2__3__1_ ( .D(s4_refreshed[33]), .CK(clk), .Q(
        s4_regOut_2__3__1_), .QN() );
  DFF_X1 s4_regOut_reg_2__3__2_ ( .D(s4_refreshed[34]), .CK(clk), .Q(
        s4_regOut_2__3__2_), .QN() );
  DFF_X1 s4_regOut_reg_2__3__3_ ( .D(s4_refreshed[35]), .CK(clk), .Q(
        s4_regOut_2__3__3_), .QN() );
  DFF_X1 s4_regOut_reg_2__4__0_ ( .D(stage3Out[32]), .CK(clk), .Q(
        stage4Out[32]), .QN() );
  DFF_X1 s4_regOut_reg_2__4__1_ ( .D(stage3Out[33]), .CK(clk), .Q(
        stage4Out[33]), .QN() );
  DFF_X1 s4_regOut_reg_2__4__2_ ( .D(stage3Out[34]), .CK(clk), .Q(
        stage4Out[34]), .QN() );
  DFF_X1 s4_regOut_reg_2__4__3_ ( .D(stage3Out[35]), .CK(clk), .Q(
        stage4Out[35]), .QN() );
  XNOR2_X1 s4_mul1_2_2_U6 ( .A(s4_mul1_2_2_n14), .B(s4_mul1_2_2_n13), .ZN(
        s4_concat[33]) );
  NAND2_X1 s4_mul1_2_2_U5 ( .A1(stage3Out[31]), .A2(s4_inv_out_2__1_), .ZN(
        s4_mul1_2_2_n14) );
  XNOR2_X1 s4_mul1_2_2_U4 ( .A(s4_mul1_2_2_n13), .B(s4_mul1_2_2_n12), .ZN(
        s4_concat[32]) );
  NAND2_X1 s4_mul1_2_2_U3 ( .A1(s4_inv_out_2__0_), .A2(stage3Out[30]), .ZN(
        s4_mul1_2_2_n12) );
  AOI221_X1 s4_mul1_2_2_U2 ( .B1(s4_inv_out_2__0_), .B2(s4_inv_out_2__1_), 
        .C1(stage3Out[31]), .C2(stage3Out[30]), .A(s4_mul1_2_2_n11), .ZN(
        s4_mul1_2_2_n13) );
  OAI22_X1 s4_mul1_2_2_U1 ( .A1(s4_inv_out_2__0_), .A2(s4_inv_out_2__1_), .B1(
        stage3Out[30]), .B2(stage3Out[31]), .ZN(s4_mul1_2_2_n11) );
  XNOR2_X1 s4_mul1_2_1_U6 ( .A(s4_mul1_2_1_n14), .B(s4_mul1_2_1_n13), .ZN(
        s4_concat[29]) );
  NAND2_X1 s4_mul1_2_1_U5 ( .A1(stage3Out[31]), .A2(s4_inv_out_1__1_), .ZN(
        s4_mul1_2_1_n14) );
  XNOR2_X1 s4_mul1_2_1_U4 ( .A(s4_mul1_2_1_n13), .B(s4_mul1_2_1_n12), .ZN(
        s4_concat[28]) );
  NAND2_X1 s4_mul1_2_1_U3 ( .A1(s4_inv_out_1__0_), .A2(stage3Out[30]), .ZN(
        s4_mul1_2_1_n12) );
  AOI221_X1 s4_mul1_2_1_U2 ( .B1(s4_inv_out_1__0_), .B2(s4_inv_out_1__1_), 
        .C1(stage3Out[31]), .C2(stage3Out[30]), .A(s4_mul1_2_1_n11), .ZN(
        s4_mul1_2_1_n13) );
  OAI22_X1 s4_mul1_2_1_U1 ( .A1(s4_inv_out_1__0_), .A2(s4_inv_out_1__1_), .B1(
        stage3Out[30]), .B2(stage3Out[31]), .ZN(s4_mul1_2_1_n11) );
  XNOR2_X1 s4_mul1_2_0_U6 ( .A(s4_mul1_2_0_n14), .B(s4_mul1_2_0_n13), .ZN(
        s4_concat[25]) );
  NAND2_X1 s4_mul1_2_0_U5 ( .A1(stage3Out[31]), .A2(s4_inv_out_0__1_), .ZN(
        s4_mul1_2_0_n14) );
  XNOR2_X1 s4_mul1_2_0_U4 ( .A(s4_mul1_2_0_n13), .B(s4_mul1_2_0_n12), .ZN(
        s4_concat[24]) );
  NAND2_X1 s4_mul1_2_0_U3 ( .A1(s4_inv_out_0__0_), .A2(stage3Out[30]), .ZN(
        s4_mul1_2_0_n12) );
  AOI221_X1 s4_mul1_2_0_U2 ( .B1(s4_inv_out_0__0_), .B2(s4_inv_out_0__1_), 
        .C1(stage3Out[31]), .C2(stage3Out[30]), .A(s4_mul1_2_0_n11), .ZN(
        s4_mul1_2_0_n13) );
  OAI22_X1 s4_mul1_2_0_U1 ( .A1(s4_inv_out_0__0_), .A2(s4_inv_out_0__1_), .B1(
        stage3Out[30]), .B2(stage3Out[31]), .ZN(s4_mul1_2_0_n11) );
  XNOR2_X1 s4_mul1_1_2_U6 ( .A(s4_mul1_1_2_n14), .B(s4_mul1_1_2_n13), .ZN(
        s4_concat[21]) );
  NAND2_X1 s4_mul1_1_2_U5 ( .A1(stage3Out[19]), .A2(s4_inv_out_2__1_), .ZN(
        s4_mul1_1_2_n14) );
  XNOR2_X1 s4_mul1_1_2_U4 ( .A(s4_mul1_1_2_n13), .B(s4_mul1_1_2_n12), .ZN(
        s4_concat[20]) );
  NAND2_X1 s4_mul1_1_2_U3 ( .A1(s4_inv_out_2__0_), .A2(stage3Out[18]), .ZN(
        s4_mul1_1_2_n12) );
  AOI221_X1 s4_mul1_1_2_U2 ( .B1(s4_inv_out_2__0_), .B2(s4_inv_out_2__1_), 
        .C1(stage3Out[19]), .C2(stage3Out[18]), .A(s4_mul1_1_2_n11), .ZN(
        s4_mul1_1_2_n13) );
  OAI22_X1 s4_mul1_1_2_U1 ( .A1(s4_inv_out_2__0_), .A2(s4_inv_out_2__1_), .B1(
        stage3Out[18]), .B2(stage3Out[19]), .ZN(s4_mul1_1_2_n11) );
  XNOR2_X1 s4_mul1_1_1_U6 ( .A(s4_mul1_1_1_n14), .B(s4_mul1_1_1_n13), .ZN(
        s4_concat[17]) );
  NAND2_X1 s4_mul1_1_1_U5 ( .A1(stage3Out[19]), .A2(s4_inv_out_1__1_), .ZN(
        s4_mul1_1_1_n14) );
  XNOR2_X1 s4_mul1_1_1_U4 ( .A(s4_mul1_1_1_n13), .B(s4_mul1_1_1_n12), .ZN(
        s4_concat[16]) );
  NAND2_X1 s4_mul1_1_1_U3 ( .A1(s4_inv_out_1__0_), .A2(stage3Out[18]), .ZN(
        s4_mul1_1_1_n12) );
  AOI221_X1 s4_mul1_1_1_U2 ( .B1(s4_inv_out_1__0_), .B2(s4_inv_out_1__1_), 
        .C1(stage3Out[19]), .C2(stage3Out[18]), .A(s4_mul1_1_1_n11), .ZN(
        s4_mul1_1_1_n13) );
  OAI22_X1 s4_mul1_1_1_U1 ( .A1(s4_inv_out_1__0_), .A2(s4_inv_out_1__1_), .B1(
        stage3Out[18]), .B2(stage3Out[19]), .ZN(s4_mul1_1_1_n11) );
  XNOR2_X1 s4_mul1_1_0_U6 ( .A(s4_mul1_1_0_n14), .B(s4_mul1_1_0_n13), .ZN(
        s4_concat[13]) );
  NAND2_X1 s4_mul1_1_0_U5 ( .A1(stage3Out[19]), .A2(s4_inv_out_0__1_), .ZN(
        s4_mul1_1_0_n14) );
  XNOR2_X1 s4_mul1_1_0_U4 ( .A(s4_mul1_1_0_n13), .B(s4_mul1_1_0_n12), .ZN(
        s4_concat[12]) );
  NAND2_X1 s4_mul1_1_0_U3 ( .A1(s4_inv_out_0__0_), .A2(stage3Out[18]), .ZN(
        s4_mul1_1_0_n12) );
  AOI221_X1 s4_mul1_1_0_U2 ( .B1(s4_inv_out_0__0_), .B2(s4_inv_out_0__1_), 
        .C1(stage3Out[19]), .C2(stage3Out[18]), .A(s4_mul1_1_0_n11), .ZN(
        s4_mul1_1_0_n13) );
  OAI22_X1 s4_mul1_1_0_U1 ( .A1(s4_inv_out_0__0_), .A2(s4_inv_out_0__1_), .B1(
        stage3Out[18]), .B2(stage3Out[19]), .ZN(s4_mul1_1_0_n11) );
  XNOR2_X1 s4_mul1_0_2_U6 ( .A(s4_mul1_0_2_n14), .B(s4_mul1_0_2_n13), .ZN(
        s4_concat[9]) );
  NAND2_X1 s4_mul1_0_2_U5 ( .A1(stage3Out[7]), .A2(s4_inv_out_2__1_), .ZN(
        s4_mul1_0_2_n14) );
  XNOR2_X1 s4_mul1_0_2_U4 ( .A(s4_mul1_0_2_n13), .B(s4_mul1_0_2_n12), .ZN(
        s4_concat[8]) );
  NAND2_X1 s4_mul1_0_2_U3 ( .A1(s4_inv_out_2__0_), .A2(stage3Out[6]), .ZN(
        s4_mul1_0_2_n12) );
  AOI221_X1 s4_mul1_0_2_U2 ( .B1(s4_inv_out_2__0_), .B2(s4_inv_out_2__1_), 
        .C1(stage3Out[7]), .C2(stage3Out[6]), .A(s4_mul1_0_2_n11), .ZN(
        s4_mul1_0_2_n13) );
  OAI22_X1 s4_mul1_0_2_U1 ( .A1(s4_inv_out_2__0_), .A2(s4_inv_out_2__1_), .B1(
        stage3Out[6]), .B2(stage3Out[7]), .ZN(s4_mul1_0_2_n11) );
  XNOR2_X1 s4_mul1_0_1_U6 ( .A(s4_mul1_0_1_n14), .B(s4_mul1_0_1_n13), .ZN(
        s4_concat[5]) );
  NAND2_X1 s4_mul1_0_1_U5 ( .A1(stage3Out[7]), .A2(s4_inv_out_1__1_), .ZN(
        s4_mul1_0_1_n14) );
  XNOR2_X1 s4_mul1_0_1_U4 ( .A(s4_mul1_0_1_n13), .B(s4_mul1_0_1_n12), .ZN(
        s4_concat[4]) );
  NAND2_X1 s4_mul1_0_1_U3 ( .A1(s4_inv_out_1__0_), .A2(stage3Out[6]), .ZN(
        s4_mul1_0_1_n12) );
  AOI221_X1 s4_mul1_0_1_U2 ( .B1(s4_inv_out_1__0_), .B2(s4_inv_out_1__1_), 
        .C1(stage3Out[7]), .C2(stage3Out[6]), .A(s4_mul1_0_1_n11), .ZN(
        s4_mul1_0_1_n13) );
  OAI22_X1 s4_mul1_0_1_U1 ( .A1(s4_inv_out_1__0_), .A2(s4_inv_out_1__1_), .B1(
        stage3Out[6]), .B2(stage3Out[7]), .ZN(s4_mul1_0_1_n11) );
  XNOR2_X1 s4_mul1_0_0_U6 ( .A(s4_mul1_0_0_n14), .B(s4_mul1_0_0_n13), .ZN(
        s4_concat[1]) );
  NAND2_X1 s4_mul1_0_0_U5 ( .A1(stage3Out[7]), .A2(s4_inv_out_0__1_), .ZN(
        s4_mul1_0_0_n14) );
  XNOR2_X1 s4_mul1_0_0_U4 ( .A(s4_mul1_0_0_n13), .B(s4_mul1_0_0_n12), .ZN(
        s4_concat[0]) );
  NAND2_X1 s4_mul1_0_0_U3 ( .A1(s4_inv_out_0__0_), .A2(stage3Out[6]), .ZN(
        s4_mul1_0_0_n12) );
  AOI221_X1 s4_mul1_0_0_U2 ( .B1(s4_inv_out_0__0_), .B2(s4_inv_out_0__1_), 
        .C1(stage3Out[7]), .C2(stage3Out[6]), .A(s4_mul1_0_0_n11), .ZN(
        s4_mul1_0_0_n13) );
  OAI22_X1 s4_mul1_0_0_U1 ( .A1(s4_inv_out_0__0_), .A2(s4_inv_out_0__1_), .B1(
        stage3Out[6]), .B2(stage3Out[7]), .ZN(s4_mul1_0_0_n11) );
  XNOR2_X1 s4_mul2_2_2_U6 ( .A(s4_mul2_2_2_n14), .B(s4_mul2_2_2_n13), .ZN(
        s4_concat[35]) );
  NAND2_X1 s4_mul2_2_2_U5 ( .A1(stage3Out[29]), .A2(s4_inv_out_2__1_), .ZN(
        s4_mul2_2_2_n14) );
  XNOR2_X1 s4_mul2_2_2_U4 ( .A(s4_mul2_2_2_n13), .B(s4_mul2_2_2_n12), .ZN(
        s4_concat[34]) );
  NAND2_X1 s4_mul2_2_2_U3 ( .A1(s4_inv_out_2__0_), .A2(stage3Out[28]), .ZN(
        s4_mul2_2_2_n12) );
  AOI221_X1 s4_mul2_2_2_U2 ( .B1(s4_inv_out_2__0_), .B2(s4_inv_out_2__1_), 
        .C1(stage3Out[29]), .C2(stage3Out[28]), .A(s4_mul2_2_2_n11), .ZN(
        s4_mul2_2_2_n13) );
  OAI22_X1 s4_mul2_2_2_U1 ( .A1(s4_inv_out_2__0_), .A2(s4_inv_out_2__1_), .B1(
        stage3Out[28]), .B2(stage3Out[29]), .ZN(s4_mul2_2_2_n11) );
  XNOR2_X1 s4_mul2_2_1_U6 ( .A(s4_mul2_2_1_n14), .B(s4_mul2_2_1_n13), .ZN(
        s4_concat[31]) );
  NAND2_X1 s4_mul2_2_1_U5 ( .A1(stage3Out[29]), .A2(s4_inv_out_1__1_), .ZN(
        s4_mul2_2_1_n14) );
  XNOR2_X1 s4_mul2_2_1_U4 ( .A(s4_mul2_2_1_n13), .B(s4_mul2_2_1_n12), .ZN(
        s4_concat[30]) );
  NAND2_X1 s4_mul2_2_1_U3 ( .A1(s4_inv_out_1__0_), .A2(stage3Out[28]), .ZN(
        s4_mul2_2_1_n12) );
  AOI221_X1 s4_mul2_2_1_U2 ( .B1(s4_inv_out_1__0_), .B2(s4_inv_out_1__1_), 
        .C1(stage3Out[29]), .C2(stage3Out[28]), .A(s4_mul2_2_1_n11), .ZN(
        s4_mul2_2_1_n13) );
  OAI22_X1 s4_mul2_2_1_U1 ( .A1(s4_inv_out_1__0_), .A2(s4_inv_out_1__1_), .B1(
        stage3Out[28]), .B2(stage3Out[29]), .ZN(s4_mul2_2_1_n11) );
  XNOR2_X1 s4_mul2_2_0_U6 ( .A(s4_mul2_2_0_n14), .B(s4_mul2_2_0_n13), .ZN(
        s4_concat[27]) );
  NAND2_X1 s4_mul2_2_0_U5 ( .A1(stage3Out[29]), .A2(s4_inv_out_0__1_), .ZN(
        s4_mul2_2_0_n14) );
  XNOR2_X1 s4_mul2_2_0_U4 ( .A(s4_mul2_2_0_n13), .B(s4_mul2_2_0_n12), .ZN(
        s4_concat[26]) );
  NAND2_X1 s4_mul2_2_0_U3 ( .A1(s4_inv_out_0__0_), .A2(stage3Out[28]), .ZN(
        s4_mul2_2_0_n12) );
  AOI221_X1 s4_mul2_2_0_U2 ( .B1(s4_inv_out_0__0_), .B2(s4_inv_out_0__1_), 
        .C1(stage3Out[29]), .C2(stage3Out[28]), .A(s4_mul2_2_0_n11), .ZN(
        s4_mul2_2_0_n13) );
  OAI22_X1 s4_mul2_2_0_U1 ( .A1(s4_inv_out_0__0_), .A2(s4_inv_out_0__1_), .B1(
        stage3Out[28]), .B2(stage3Out[29]), .ZN(s4_mul2_2_0_n11) );
  XNOR2_X1 s4_mul2_1_2_U6 ( .A(s4_mul2_1_2_n14), .B(s4_mul2_1_2_n13), .ZN(
        s4_concat[23]) );
  NAND2_X1 s4_mul2_1_2_U5 ( .A1(stage3Out[17]), .A2(s4_inv_out_2__1_), .ZN(
        s4_mul2_1_2_n14) );
  XNOR2_X1 s4_mul2_1_2_U4 ( .A(s4_mul2_1_2_n13), .B(s4_mul2_1_2_n12), .ZN(
        s4_concat[22]) );
  NAND2_X1 s4_mul2_1_2_U3 ( .A1(s4_inv_out_2__0_), .A2(stage3Out[16]), .ZN(
        s4_mul2_1_2_n12) );
  AOI221_X1 s4_mul2_1_2_U2 ( .B1(s4_inv_out_2__0_), .B2(s4_inv_out_2__1_), 
        .C1(stage3Out[17]), .C2(stage3Out[16]), .A(s4_mul2_1_2_n11), .ZN(
        s4_mul2_1_2_n13) );
  OAI22_X1 s4_mul2_1_2_U1 ( .A1(s4_inv_out_2__0_), .A2(s4_inv_out_2__1_), .B1(
        stage3Out[16]), .B2(stage3Out[17]), .ZN(s4_mul2_1_2_n11) );
  XNOR2_X1 s4_mul2_1_1_U6 ( .A(s4_mul2_1_1_n14), .B(s4_mul2_1_1_n13), .ZN(
        s4_concat[19]) );
  NAND2_X1 s4_mul2_1_1_U5 ( .A1(stage3Out[17]), .A2(s4_inv_out_1__1_), .ZN(
        s4_mul2_1_1_n14) );
  XNOR2_X1 s4_mul2_1_1_U4 ( .A(s4_mul2_1_1_n13), .B(s4_mul2_1_1_n12), .ZN(
        s4_concat[18]) );
  NAND2_X1 s4_mul2_1_1_U3 ( .A1(s4_inv_out_1__0_), .A2(stage3Out[16]), .ZN(
        s4_mul2_1_1_n12) );
  AOI221_X1 s4_mul2_1_1_U2 ( .B1(s4_inv_out_1__0_), .B2(s4_inv_out_1__1_), 
        .C1(stage3Out[17]), .C2(stage3Out[16]), .A(s4_mul2_1_1_n11), .ZN(
        s4_mul2_1_1_n13) );
  OAI22_X1 s4_mul2_1_1_U1 ( .A1(s4_inv_out_1__0_), .A2(s4_inv_out_1__1_), .B1(
        stage3Out[16]), .B2(stage3Out[17]), .ZN(s4_mul2_1_1_n11) );
  XNOR2_X1 s4_mul2_1_0_U6 ( .A(s4_mul2_1_0_n14), .B(s4_mul2_1_0_n13), .ZN(
        s4_concat[15]) );
  NAND2_X1 s4_mul2_1_0_U5 ( .A1(stage3Out[17]), .A2(s4_inv_out_0__1_), .ZN(
        s4_mul2_1_0_n14) );
  XNOR2_X1 s4_mul2_1_0_U4 ( .A(s4_mul2_1_0_n13), .B(s4_mul2_1_0_n12), .ZN(
        s4_concat[14]) );
  NAND2_X1 s4_mul2_1_0_U3 ( .A1(s4_inv_out_0__0_), .A2(stage3Out[16]), .ZN(
        s4_mul2_1_0_n12) );
  AOI221_X1 s4_mul2_1_0_U2 ( .B1(s4_inv_out_0__0_), .B2(s4_inv_out_0__1_), 
        .C1(stage3Out[17]), .C2(stage3Out[16]), .A(s4_mul2_1_0_n11), .ZN(
        s4_mul2_1_0_n13) );
  OAI22_X1 s4_mul2_1_0_U1 ( .A1(s4_inv_out_0__0_), .A2(s4_inv_out_0__1_), .B1(
        stage3Out[16]), .B2(stage3Out[17]), .ZN(s4_mul2_1_0_n11) );
  XNOR2_X1 s4_mul2_0_2_U6 ( .A(s4_mul2_0_2_n14), .B(s4_mul2_0_2_n13), .ZN(
        s4_concat[11]) );
  NAND2_X1 s4_mul2_0_2_U5 ( .A1(stage3Out[5]), .A2(s4_inv_out_2__1_), .ZN(
        s4_mul2_0_2_n14) );
  XNOR2_X1 s4_mul2_0_2_U4 ( .A(s4_mul2_0_2_n13), .B(s4_mul2_0_2_n12), .ZN(
        s4_concat[10]) );
  NAND2_X1 s4_mul2_0_2_U3 ( .A1(s4_inv_out_2__0_), .A2(stage3Out[4]), .ZN(
        s4_mul2_0_2_n12) );
  AOI221_X1 s4_mul2_0_2_U2 ( .B1(s4_inv_out_2__0_), .B2(s4_inv_out_2__1_), 
        .C1(stage3Out[5]), .C2(stage3Out[4]), .A(s4_mul2_0_2_n11), .ZN(
        s4_mul2_0_2_n13) );
  OAI22_X1 s4_mul2_0_2_U1 ( .A1(s4_inv_out_2__0_), .A2(s4_inv_out_2__1_), .B1(
        stage3Out[4]), .B2(stage3Out[5]), .ZN(s4_mul2_0_2_n11) );
  XNOR2_X1 s4_mul2_0_1_U6 ( .A(s4_mul2_0_1_n14), .B(s4_mul2_0_1_n13), .ZN(
        s4_concat[7]) );
  NAND2_X1 s4_mul2_0_1_U5 ( .A1(stage3Out[5]), .A2(s4_inv_out_1__1_), .ZN(
        s4_mul2_0_1_n14) );
  XNOR2_X1 s4_mul2_0_1_U4 ( .A(s4_mul2_0_1_n13), .B(s4_mul2_0_1_n12), .ZN(
        s4_concat[6]) );
  NAND2_X1 s4_mul2_0_1_U3 ( .A1(s4_inv_out_1__0_), .A2(stage3Out[4]), .ZN(
        s4_mul2_0_1_n12) );
  AOI221_X1 s4_mul2_0_1_U2 ( .B1(s4_inv_out_1__0_), .B2(s4_inv_out_1__1_), 
        .C1(stage3Out[5]), .C2(stage3Out[4]), .A(s4_mul2_0_1_n11), .ZN(
        s4_mul2_0_1_n13) );
  OAI22_X1 s4_mul2_0_1_U1 ( .A1(s4_inv_out_1__0_), .A2(s4_inv_out_1__1_), .B1(
        stage3Out[4]), .B2(stage3Out[5]), .ZN(s4_mul2_0_1_n11) );
  XNOR2_X1 s4_mul2_0_0_U6 ( .A(s4_mul2_0_0_n14), .B(s4_mul2_0_0_n13), .ZN(
        s4_concat[3]) );
  NAND2_X1 s4_mul2_0_0_U5 ( .A1(stage3Out[5]), .A2(s4_inv_out_0__1_), .ZN(
        s4_mul2_0_0_n14) );
  XNOR2_X1 s4_mul2_0_0_U4 ( .A(s4_mul2_0_0_n13), .B(s4_mul2_0_0_n12), .ZN(
        s4_concat[2]) );
  NAND2_X1 s4_mul2_0_0_U3 ( .A1(s4_inv_out_0__0_), .A2(stage3Out[4]), .ZN(
        s4_mul2_0_0_n12) );
  AOI221_X1 s4_mul2_0_0_U2 ( .B1(s4_inv_out_0__0_), .B2(s4_inv_out_0__1_), 
        .C1(stage3Out[5]), .C2(stage3Out[4]), .A(s4_mul2_0_0_n11), .ZN(
        s4_mul2_0_0_n13) );
  OAI22_X1 s4_mul2_0_0_U1 ( .A1(s4_inv_out_0__0_), .A2(s4_inv_out_0__1_), .B1(
        stage3Out[4]), .B2(stage3Out[5]), .ZN(s4_mul2_0_0_n11) );
  XOR2_X1 s4_compr_0_0_U4 ( .A(s4_regOut_0__1__3_), .B(s4_regOut_0__2__3_), 
        .Z(s4_chain_0__1__3_) );
  XOR2_X1 s4_compr_0_0_U3 ( .A(s4_regOut_0__1__2_), .B(s4_regOut_0__2__2_), 
        .Z(s4_chain_0__1__2_) );
  XOR2_X1 s4_compr_0_0_U2 ( .A(s4_regOut_0__1__1_), .B(s4_regOut_0__2__1_), 
        .Z(s4_chain_0__1__1_) );
  XOR2_X1 s4_compr_0_0_U1 ( .A(s4_regOut_0__1__0_), .B(s4_regOut_0__2__0_), 
        .Z(s4_chain_0__1__0_) );
  XOR2_X1 s4_compr_0_1_U4 ( .A(s4_chain_0__1__3_), .B(s4_regOut_0__3__3_), .Z(
        stage4Out[7]) );
  XOR2_X1 s4_compr_0_1_U3 ( .A(s4_chain_0__1__2_), .B(s4_regOut_0__3__2_), .Z(
        stage4Out[6]) );
  XOR2_X1 s4_compr_0_1_U2 ( .A(s4_chain_0__1__1_), .B(s4_regOut_0__3__1_), .Z(
        stage4Out[5]) );
  XOR2_X1 s4_compr_0_1_U1 ( .A(s4_chain_0__1__0_), .B(s4_regOut_0__3__0_), .Z(
        stage4Out[4]) );
  XOR2_X1 s4_compr_1_0_U4 ( .A(s4_regOut_1__1__3_), .B(s4_regOut_1__2__3_), 
        .Z(s4_chain_1__1__3_) );
  XOR2_X1 s4_compr_1_0_U3 ( .A(s4_regOut_1__1__2_), .B(s4_regOut_1__2__2_), 
        .Z(s4_chain_1__1__2_) );
  XOR2_X1 s4_compr_1_0_U2 ( .A(s4_regOut_1__1__1_), .B(s4_regOut_1__2__1_), 
        .Z(s4_chain_1__1__1_) );
  XOR2_X1 s4_compr_1_0_U1 ( .A(s4_regOut_1__1__0_), .B(s4_regOut_1__2__0_), 
        .Z(s4_chain_1__1__0_) );
  XOR2_X1 s4_compr_1_1_U4 ( .A(s4_chain_1__1__3_), .B(s4_regOut_1__3__3_), .Z(
        stage4Out[19]) );
  XOR2_X1 s4_compr_1_1_U3 ( .A(s4_chain_1__1__2_), .B(s4_regOut_1__3__2_), .Z(
        stage4Out[18]) );
  XOR2_X1 s4_compr_1_1_U2 ( .A(s4_chain_1__1__1_), .B(s4_regOut_1__3__1_), .Z(
        stage4Out[17]) );
  XOR2_X1 s4_compr_1_1_U1 ( .A(s4_chain_1__1__0_), .B(s4_regOut_1__3__0_), .Z(
        stage4Out[16]) );
  XOR2_X1 s4_compr_2_0_U4 ( .A(s4_regOut_2__1__3_), .B(s4_regOut_2__2__3_), 
        .Z(s4_chain_2__1__3_) );
  XOR2_X1 s4_compr_2_0_U3 ( .A(s4_regOut_2__1__2_), .B(s4_regOut_2__2__2_), 
        .Z(s4_chain_2__1__2_) );
  XOR2_X1 s4_compr_2_0_U2 ( .A(s4_regOut_2__1__1_), .B(s4_regOut_2__2__1_), 
        .Z(s4_chain_2__1__1_) );
  XOR2_X1 s4_compr_2_0_U1 ( .A(s4_regOut_2__1__0_), .B(s4_regOut_2__2__0_), 
        .Z(s4_chain_2__1__0_) );
  XOR2_X1 s4_compr_2_1_U4 ( .A(s4_chain_2__1__3_), .B(s4_regOut_2__3__3_), .Z(
        stage4Out[31]) );
  XOR2_X1 s4_compr_2_1_U3 ( .A(s4_chain_2__1__2_), .B(s4_regOut_2__3__2_), .Z(
        stage4Out[30]) );
  XOR2_X1 s4_compr_2_1_U2 ( .A(s4_chain_2__1__1_), .B(s4_regOut_2__3__1_), .Z(
        stage4Out[29]) );
  XOR2_X1 s4_compr_2_1_U1 ( .A(s4_chain_2__1__0_), .B(s4_regOut_2__3__0_), .Z(
        stage4Out[28]) );
  XNOR2_X1 s5_U158 ( .A(s5_n84), .B(s5_concat[71]), .ZN(s5_refreshed[71]) );
  XNOR2_X1 s5_U157 ( .A(randomS5[7]), .B(randomS5[15]), .ZN(s5_n84) );
  XNOR2_X1 s5_U156 ( .A(s5_n83), .B(s5_concat[70]), .ZN(s5_refreshed[70]) );
  XNOR2_X1 s5_U155 ( .A(randomS5[6]), .B(randomS5[14]), .ZN(s5_n83) );
  XNOR2_X1 s5_U154 ( .A(s5_n82), .B(s5_concat[69]), .ZN(s5_refreshed[69]) );
  XNOR2_X1 s5_U153 ( .A(randomS5[5]), .B(randomS5[13]), .ZN(s5_n82) );
  XNOR2_X1 s5_U152 ( .A(s5_n81), .B(s5_concat[68]), .ZN(s5_refreshed[68]) );
  XNOR2_X1 s5_U151 ( .A(randomS5[4]), .B(randomS5[12]), .ZN(s5_n81) );
  XNOR2_X1 s5_U150 ( .A(s5_n80), .B(s5_concat[67]), .ZN(s5_refreshed[67]) );
  XNOR2_X1 s5_U149 ( .A(randomS5[3]), .B(randomS5[11]), .ZN(s5_n80) );
  XNOR2_X1 s5_U148 ( .A(s5_n79), .B(s5_concat[66]), .ZN(s5_refreshed[66]) );
  XNOR2_X1 s5_U147 ( .A(randomS5[2]), .B(randomS5[10]), .ZN(s5_n79) );
  XNOR2_X1 s5_U146 ( .A(s5_n78), .B(s5_concat[65]), .ZN(s5_refreshed[65]) );
  XNOR2_X1 s5_U145 ( .A(randomS5[1]), .B(randomS5[9]), .ZN(s5_n78) );
  XNOR2_X1 s5_U144 ( .A(s5_n77), .B(s5_concat[64]), .ZN(s5_refreshed[64]) );
  XNOR2_X1 s5_U143 ( .A(randomS5[0]), .B(randomS5[8]), .ZN(s5_n77) );
  XNOR2_X1 s5_U142 ( .A(s5_n76), .B(s5_concat[63]), .ZN(s5_refreshed[63]) );
  XNOR2_X1 s5_U141 ( .A(randomS5[23]), .B(randomS5[15]), .ZN(s5_n76) );
  XNOR2_X1 s5_U140 ( .A(s5_n75), .B(s5_concat[62]), .ZN(s5_refreshed[62]) );
  XNOR2_X1 s5_U139 ( .A(randomS5[22]), .B(randomS5[14]), .ZN(s5_n75) );
  XNOR2_X1 s5_U138 ( .A(s5_n74), .B(s5_concat[61]), .ZN(s5_refreshed[61]) );
  XNOR2_X1 s5_U137 ( .A(randomS5[21]), .B(randomS5[13]), .ZN(s5_n74) );
  XNOR2_X1 s5_U136 ( .A(s5_n73), .B(s5_concat[60]), .ZN(s5_refreshed[60]) );
  XNOR2_X1 s5_U135 ( .A(randomS5[20]), .B(randomS5[12]), .ZN(s5_n73) );
  XNOR2_X1 s5_U134 ( .A(s5_n72), .B(s5_concat[59]), .ZN(s5_refreshed[59]) );
  XNOR2_X1 s5_U133 ( .A(randomS5[19]), .B(randomS5[11]), .ZN(s5_n72) );
  XNOR2_X1 s5_U132 ( .A(s5_n71), .B(s5_concat[58]), .ZN(s5_refreshed[58]) );
  XNOR2_X1 s5_U131 ( .A(randomS5[18]), .B(randomS5[10]), .ZN(s5_n71) );
  XNOR2_X1 s5_U130 ( .A(s5_n70), .B(s5_concat[57]), .ZN(s5_refreshed[57]) );
  XNOR2_X1 s5_U129 ( .A(randomS5[17]), .B(randomS5[9]), .ZN(s5_n70) );
  XNOR2_X1 s5_U128 ( .A(s5_n69), .B(s5_concat[56]), .ZN(s5_refreshed[56]) );
  XNOR2_X1 s5_U127 ( .A(randomS5[16]), .B(randomS5[8]), .ZN(s5_n69) );
  XNOR2_X1 s5_U126 ( .A(s5_n68), .B(s5_concat[55]), .ZN(s5_refreshed[55]) );
  XNOR2_X1 s5_U125 ( .A(randomS5[31]), .B(randomS5[23]), .ZN(s5_n68) );
  XNOR2_X1 s5_U124 ( .A(s5_n67), .B(s5_concat[54]), .ZN(s5_refreshed[54]) );
  XNOR2_X1 s5_U123 ( .A(randomS5[30]), .B(randomS5[22]), .ZN(s5_n67) );
  XNOR2_X1 s5_U122 ( .A(s5_n66), .B(s5_concat[53]), .ZN(s5_refreshed[53]) );
  XNOR2_X1 s5_U121 ( .A(randomS5[29]), .B(randomS5[21]), .ZN(s5_n66) );
  XNOR2_X1 s5_U120 ( .A(s5_n65), .B(s5_concat[52]), .ZN(s5_refreshed[52]) );
  XNOR2_X1 s5_U119 ( .A(randomS5[28]), .B(randomS5[20]), .ZN(s5_n65) );
  XNOR2_X1 s5_U118 ( .A(s5_n64), .B(s5_concat[51]), .ZN(s5_refreshed[51]) );
  XNOR2_X1 s5_U117 ( .A(randomS5[27]), .B(randomS5[19]), .ZN(s5_n64) );
  XNOR2_X1 s5_U116 ( .A(s5_n63), .B(s5_concat[50]), .ZN(s5_refreshed[50]) );
  XNOR2_X1 s5_U115 ( .A(randomS5[26]), .B(randomS5[18]), .ZN(s5_n63) );
  XNOR2_X1 s5_U114 ( .A(s5_n62), .B(s5_concat[49]), .ZN(s5_refreshed[49]) );
  XNOR2_X1 s5_U113 ( .A(randomS5[25]), .B(randomS5[17]), .ZN(s5_n62) );
  XNOR2_X1 s5_U112 ( .A(s5_n61), .B(s5_concat[48]), .ZN(s5_refreshed[48]) );
  XNOR2_X1 s5_U111 ( .A(randomS5[24]), .B(randomS5[16]), .ZN(s5_n61) );
  XNOR2_X1 s5_U110 ( .A(s5_n60), .B(s5_concat[47]), .ZN(s5_refreshed[47]) );
  XNOR2_X1 s5_U109 ( .A(randomS5[39]), .B(randomS5[31]), .ZN(s5_n60) );
  XNOR2_X1 s5_U108 ( .A(s5_n59), .B(s5_concat[46]), .ZN(s5_refreshed[46]) );
  XNOR2_X1 s5_U107 ( .A(randomS5[38]), .B(randomS5[30]), .ZN(s5_n59) );
  XNOR2_X1 s5_U106 ( .A(s5_n58), .B(s5_concat[45]), .ZN(s5_refreshed[45]) );
  XNOR2_X1 s5_U105 ( .A(randomS5[37]), .B(randomS5[29]), .ZN(s5_n58) );
  XNOR2_X1 s5_U104 ( .A(s5_n57), .B(s5_concat[44]), .ZN(s5_refreshed[44]) );
  XNOR2_X1 s5_U103 ( .A(randomS5[36]), .B(randomS5[28]), .ZN(s5_n57) );
  XNOR2_X1 s5_U102 ( .A(s5_n56), .B(s5_concat[43]), .ZN(s5_refreshed[43]) );
  XNOR2_X1 s5_U101 ( .A(randomS5[35]), .B(randomS5[27]), .ZN(s5_n56) );
  XNOR2_X1 s5_U100 ( .A(s5_n55), .B(s5_concat[42]), .ZN(s5_refreshed[42]) );
  XNOR2_X1 s5_U99 ( .A(randomS5[34]), .B(randomS5[26]), .ZN(s5_n55) );
  XNOR2_X1 s5_U98 ( .A(s5_n54), .B(s5_concat[41]), .ZN(s5_refreshed[41]) );
  XNOR2_X1 s5_U97 ( .A(randomS5[33]), .B(randomS5[25]), .ZN(s5_n54) );
  XNOR2_X1 s5_U96 ( .A(s5_n53), .B(s5_concat[40]), .ZN(s5_refreshed[40]) );
  XNOR2_X1 s5_U95 ( .A(randomS5[32]), .B(randomS5[24]), .ZN(s5_n53) );
  XNOR2_X1 s5_U94 ( .A(s5_n52), .B(s5_concat[39]), .ZN(s5_refreshed[39]) );
  XNOR2_X1 s5_U93 ( .A(randomS5[47]), .B(randomS5[39]), .ZN(s5_n52) );
  XNOR2_X1 s5_U92 ( .A(s5_n51), .B(s5_concat[38]), .ZN(s5_refreshed[38]) );
  XNOR2_X1 s5_U91 ( .A(randomS5[46]), .B(randomS5[38]), .ZN(s5_n51) );
  XNOR2_X1 s5_U90 ( .A(s5_n50), .B(s5_concat[37]), .ZN(s5_refreshed[37]) );
  XNOR2_X1 s5_U89 ( .A(randomS5[45]), .B(randomS5[37]), .ZN(s5_n50) );
  XNOR2_X1 s5_U88 ( .A(s5_n49), .B(s5_concat[36]), .ZN(s5_refreshed[36]) );
  XNOR2_X1 s5_U87 ( .A(randomS5[44]), .B(randomS5[36]), .ZN(s5_n49) );
  XNOR2_X1 s5_U86 ( .A(s5_n48), .B(s5_concat[35]), .ZN(s5_refreshed[35]) );
  XNOR2_X1 s5_U85 ( .A(randomS5[43]), .B(randomS5[35]), .ZN(s5_n48) );
  XNOR2_X1 s5_U84 ( .A(s5_n47), .B(s5_concat[34]), .ZN(s5_refreshed[34]) );
  XNOR2_X1 s5_U83 ( .A(randomS5[42]), .B(randomS5[34]), .ZN(s5_n47) );
  XNOR2_X1 s5_U82 ( .A(s5_n46), .B(s5_concat[33]), .ZN(s5_refreshed[33]) );
  XNOR2_X1 s5_U81 ( .A(randomS5[41]), .B(randomS5[33]), .ZN(s5_n46) );
  XNOR2_X1 s5_U80 ( .A(s5_n45), .B(s5_concat[32]), .ZN(s5_refreshed[32]) );
  XNOR2_X1 s5_U79 ( .A(randomS5[40]), .B(randomS5[32]), .ZN(s5_n45) );
  XNOR2_X1 s5_U78 ( .A(s5_n44), .B(s5_concat[31]), .ZN(s5_refreshed[31]) );
  XNOR2_X1 s5_U77 ( .A(randomS5[55]), .B(randomS5[47]), .ZN(s5_n44) );
  XNOR2_X1 s5_U76 ( .A(s5_n43), .B(s5_concat[30]), .ZN(s5_refreshed[30]) );
  XNOR2_X1 s5_U75 ( .A(randomS5[54]), .B(randomS5[46]), .ZN(s5_n43) );
  XNOR2_X1 s5_U74 ( .A(s5_n42), .B(s5_concat[29]), .ZN(s5_refreshed[29]) );
  XNOR2_X1 s5_U73 ( .A(randomS5[53]), .B(randomS5[45]), .ZN(s5_n42) );
  XNOR2_X1 s5_U72 ( .A(s5_n41), .B(s5_concat[28]), .ZN(s5_refreshed[28]) );
  XNOR2_X1 s5_U71 ( .A(randomS5[52]), .B(randomS5[44]), .ZN(s5_n41) );
  XNOR2_X1 s5_U70 ( .A(s5_n40), .B(s5_concat[27]), .ZN(s5_refreshed[27]) );
  XNOR2_X1 s5_U69 ( .A(randomS5[51]), .B(randomS5[43]), .ZN(s5_n40) );
  XNOR2_X1 s5_U68 ( .A(s5_n39), .B(s5_concat[26]), .ZN(s5_refreshed[26]) );
  XNOR2_X1 s5_U67 ( .A(randomS5[50]), .B(randomS5[42]), .ZN(s5_n39) );
  XNOR2_X1 s5_U66 ( .A(s5_n38), .B(s5_concat[25]), .ZN(s5_refreshed[25]) );
  XNOR2_X1 s5_U65 ( .A(randomS5[49]), .B(randomS5[41]), .ZN(s5_n38) );
  XNOR2_X1 s5_U64 ( .A(s5_n37), .B(s5_concat[24]), .ZN(s5_refreshed[24]) );
  XNOR2_X1 s5_U63 ( .A(randomS5[48]), .B(randomS5[40]), .ZN(s5_n37) );
  XNOR2_X1 s5_U62 ( .A(s5_n36), .B(s5_concat[23]), .ZN(s5_refreshed[23]) );
  XNOR2_X1 s5_U61 ( .A(randomS5[63]), .B(randomS5[55]), .ZN(s5_n36) );
  XNOR2_X1 s5_U60 ( .A(s5_n35), .B(s5_concat[22]), .ZN(s5_refreshed[22]) );
  XNOR2_X1 s5_U59 ( .A(randomS5[62]), .B(randomS5[54]), .ZN(s5_n35) );
  XNOR2_X1 s5_U58 ( .A(s5_n34), .B(s5_concat[21]), .ZN(s5_refreshed[21]) );
  XNOR2_X1 s5_U57 ( .A(randomS5[61]), .B(randomS5[53]), .ZN(s5_n34) );
  XNOR2_X1 s5_U56 ( .A(s5_n33), .B(s5_concat[20]), .ZN(s5_refreshed[20]) );
  XNOR2_X1 s5_U55 ( .A(randomS5[60]), .B(randomS5[52]), .ZN(s5_n33) );
  XNOR2_X1 s5_U54 ( .A(s5_n32), .B(s5_concat[19]), .ZN(s5_refreshed[19]) );
  XNOR2_X1 s5_U53 ( .A(randomS5[59]), .B(randomS5[51]), .ZN(s5_n32) );
  XNOR2_X1 s5_U52 ( .A(s5_n31), .B(s5_concat[18]), .ZN(s5_refreshed[18]) );
  XNOR2_X1 s5_U51 ( .A(randomS5[58]), .B(randomS5[50]), .ZN(s5_n31) );
  XNOR2_X1 s5_U50 ( .A(s5_n30), .B(s5_concat[17]), .ZN(s5_refreshed[17]) );
  XNOR2_X1 s5_U49 ( .A(randomS5[57]), .B(randomS5[49]), .ZN(s5_n30) );
  XNOR2_X1 s5_U48 ( .A(s5_n29), .B(s5_concat[16]), .ZN(s5_refreshed[16]) );
  XNOR2_X1 s5_U47 ( .A(randomS5[56]), .B(randomS5[48]), .ZN(s5_n29) );
  XNOR2_X1 s5_U46 ( .A(s5_n28), .B(s5_concat[15]), .ZN(s5_refreshed[15]) );
  XNOR2_X1 s5_U45 ( .A(randomS5[71]), .B(randomS5[63]), .ZN(s5_n28) );
  XNOR2_X1 s5_U44 ( .A(s5_n27), .B(s5_concat[14]), .ZN(s5_refreshed[14]) );
  XNOR2_X1 s5_U43 ( .A(randomS5[70]), .B(randomS5[62]), .ZN(s5_n27) );
  XNOR2_X1 s5_U42 ( .A(s5_n26), .B(s5_concat[13]), .ZN(s5_refreshed[13]) );
  XNOR2_X1 s5_U41 ( .A(randomS5[69]), .B(randomS5[61]), .ZN(s5_n26) );
  XNOR2_X1 s5_U40 ( .A(s5_n25), .B(s5_concat[12]), .ZN(s5_refreshed[12]) );
  XNOR2_X1 s5_U39 ( .A(randomS5[68]), .B(randomS5[60]), .ZN(s5_n25) );
  XNOR2_X1 s5_U38 ( .A(s5_n24), .B(s5_concat[11]), .ZN(s5_refreshed[11]) );
  XNOR2_X1 s5_U37 ( .A(randomS5[67]), .B(randomS5[59]), .ZN(s5_n24) );
  XNOR2_X1 s5_U36 ( .A(s5_n23), .B(s5_concat[10]), .ZN(s5_refreshed[10]) );
  XNOR2_X1 s5_U35 ( .A(randomS5[66]), .B(randomS5[58]), .ZN(s5_n23) );
  XNOR2_X1 s5_U34 ( .A(s5_n22), .B(s5_concat[9]), .ZN(s5_refreshed[9]) );
  XNOR2_X1 s5_U33 ( .A(randomS5[65]), .B(randomS5[57]), .ZN(s5_n22) );
  XNOR2_X1 s5_U32 ( .A(s5_n21), .B(s5_concat[8]), .ZN(s5_refreshed[8]) );
  XNOR2_X1 s5_U31 ( .A(randomS5[64]), .B(randomS5[56]), .ZN(s5_n21) );
  XNOR2_X1 s5_U30 ( .A(s5_n20), .B(s5_concat[7]), .ZN(s5_refreshed[7]) );
  XNOR2_X1 s5_U29 ( .A(randomS5[7]), .B(randomS5[71]), .ZN(s5_n20) );
  XNOR2_X1 s5_U28 ( .A(s5_n19), .B(s5_concat[6]), .ZN(s5_refreshed[6]) );
  XNOR2_X1 s5_U27 ( .A(randomS5[6]), .B(randomS5[70]), .ZN(s5_n19) );
  XNOR2_X1 s5_U26 ( .A(s5_n18), .B(s5_concat[5]), .ZN(s5_refreshed[5]) );
  XNOR2_X1 s5_U25 ( .A(randomS5[5]), .B(randomS5[69]), .ZN(s5_n18) );
  XNOR2_X1 s5_U24 ( .A(s5_n17), .B(s5_concat[4]), .ZN(s5_refreshed[4]) );
  XNOR2_X1 s5_U23 ( .A(randomS5[4]), .B(randomS5[68]), .ZN(s5_n17) );
  XNOR2_X1 s5_U22 ( .A(s5_n16), .B(s5_concat[3]), .ZN(s5_refreshed[3]) );
  XNOR2_X1 s5_U21 ( .A(randomS5[3]), .B(randomS5[67]), .ZN(s5_n16) );
  XNOR2_X1 s5_U20 ( .A(s5_n15), .B(s5_concat[2]), .ZN(s5_refreshed[2]) );
  XNOR2_X1 s5_U19 ( .A(randomS5[2]), .B(randomS5[66]), .ZN(s5_n15) );
  XNOR2_X1 s5_U18 ( .A(s5_n14), .B(s5_concat[1]), .ZN(s5_refreshed[1]) );
  XNOR2_X1 s5_U17 ( .A(randomS5[1]), .B(randomS5[65]), .ZN(s5_n14) );
  XNOR2_X1 s5_U16 ( .A(s5_n13), .B(s5_concat[0]), .ZN(s5_refreshed[0]) );
  XNOR2_X1 s5_U15 ( .A(randomS5[0]), .B(randomS5[64]), .ZN(s5_n13) );
  BUF_X2 s5_U14 ( .A(stage4Out[6]), .Z(s5_n3) );
  BUF_X2 s5_U13 ( .A(stage4Out[18]), .Z(s5_n7) );
  BUF_X2 s5_U12 ( .A(stage4Out[30]), .Z(s5_n11) );
  BUF_X2 s5_U11 ( .A(stage4Out[5]), .Z(s5_n2) );
  BUF_X2 s5_U10 ( .A(stage4Out[17]), .Z(s5_n6) );
  BUF_X2 s5_U9 ( .A(stage4Out[29]), .Z(s5_n10) );
  BUF_X2 s5_U8 ( .A(stage4Out[19]), .Z(s5_n8) );
  BUF_X2 s5_U7 ( .A(stage4Out[7]), .Z(s5_n4) );
  BUF_X2 s5_U6 ( .A(stage4Out[31]), .Z(s5_n12) );
  BUF_X2 s5_U5 ( .A(stage4Out[16]), .Z(s5_n5) );
  BUF_X2 s5_U4 ( .A(stage4Out[4]), .Z(s5_n1) );
  BUF_X2 s5_U3 ( .A(stage4Out[28]), .Z(s5_n9) );
  DFF_X1 s5_regOut_reg_0__0__0_ ( .D(s5_refreshed[0]), .CK(clk), .Q(
        s5_regOut[0]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__1_ ( .D(s5_refreshed[1]), .CK(clk), .Q(
        s5_regOut[1]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__2_ ( .D(s5_refreshed[2]), .CK(clk), .Q(
        s5_regOut[2]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__3_ ( .D(s5_refreshed[3]), .CK(clk), .Q(
        s5_regOut[3]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__4_ ( .D(s5_refreshed[4]), .CK(clk), .Q(
        s5_regOut[4]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__5_ ( .D(s5_refreshed[5]), .CK(clk), .Q(
        s5_regOut[5]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__6_ ( .D(s5_refreshed[6]), .CK(clk), .Q(
        s5_regOut[6]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__7_ ( .D(s5_refreshed[7]), .CK(clk), .Q(
        s5_regOut[7]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__0_ ( .D(s5_refreshed[8]), .CK(clk), .Q(
        s5_regOut[8]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__1_ ( .D(s5_refreshed[9]), .CK(clk), .Q(
        s5_regOut[9]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__2_ ( .D(s5_refreshed[10]), .CK(clk), .Q(
        s5_regOut[10]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__3_ ( .D(s5_refreshed[11]), .CK(clk), .Q(
        s5_regOut[11]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__4_ ( .D(s5_refreshed[12]), .CK(clk), .Q(
        s5_regOut[12]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__5_ ( .D(s5_refreshed[13]), .CK(clk), .Q(
        s5_regOut[13]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__6_ ( .D(s5_refreshed[14]), .CK(clk), .Q(
        s5_regOut[14]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__7_ ( .D(s5_refreshed[15]), .CK(clk), .Q(
        s5_regOut[15]), .QN() );
  DFF_X1 s5_regOut_reg_0__2__0_ ( .D(s5_refreshed[16]), .CK(clk), .Q(
        s5_regOut[16]), .QN() );
  DFF_X1 s5_regOut_reg_0__2__1_ ( .D(s5_refreshed[17]), .CK(clk), .Q(
        s5_regOut[17]), .QN() );
  DFF_X1 s5_regOut_reg_0__2__2_ ( .D(s5_refreshed[18]), .CK(clk), .Q(
        s5_regOut[18]), .QN() );
  DFF_X1 s5_regOut_reg_0__2__3_ ( .D(s5_refreshed[19]), .CK(clk), .Q(
        s5_regOut[19]), .QN() );
  DFF_X1 s5_regOut_reg_0__2__4_ ( .D(s5_refreshed[20]), .CK(clk), .Q(
        s5_regOut[20]), .QN() );
  DFF_X1 s5_regOut_reg_0__2__5_ ( .D(s5_refreshed[21]), .CK(clk), .Q(
        s5_regOut[21]), .QN() );
  DFF_X1 s5_regOut_reg_0__2__6_ ( .D(s5_refreshed[22]), .CK(clk), .Q(
        s5_regOut[22]), .QN() );
  DFF_X1 s5_regOut_reg_0__2__7_ ( .D(s5_refreshed[23]), .CK(clk), .Q(
        s5_regOut[23]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__0_ ( .D(s5_refreshed[24]), .CK(clk), .Q(
        s5_regOut[24]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__1_ ( .D(s5_refreshed[25]), .CK(clk), .Q(
        s5_regOut[25]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__2_ ( .D(s5_refreshed[26]), .CK(clk), .Q(
        s5_regOut[26]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__3_ ( .D(s5_refreshed[27]), .CK(clk), .Q(
        s5_regOut[27]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__4_ ( .D(s5_refreshed[28]), .CK(clk), .Q(
        s5_regOut[28]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__5_ ( .D(s5_refreshed[29]), .CK(clk), .Q(
        s5_regOut[29]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__6_ ( .D(s5_refreshed[30]), .CK(clk), .Q(
        s5_regOut[30]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__7_ ( .D(s5_refreshed[31]), .CK(clk), .Q(
        s5_regOut[31]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__0_ ( .D(s5_refreshed[32]), .CK(clk), .Q(
        s5_regOut[32]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__1_ ( .D(s5_refreshed[33]), .CK(clk), .Q(
        s5_regOut[33]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__2_ ( .D(s5_refreshed[34]), .CK(clk), .Q(
        s5_regOut[34]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__3_ ( .D(s5_refreshed[35]), .CK(clk), .Q(
        s5_regOut[35]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__4_ ( .D(s5_refreshed[36]), .CK(clk), .Q(
        s5_regOut[36]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__5_ ( .D(s5_refreshed[37]), .CK(clk), .Q(
        s5_regOut[37]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__6_ ( .D(s5_refreshed[38]), .CK(clk), .Q(
        s5_regOut[38]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__7_ ( .D(s5_refreshed[39]), .CK(clk), .Q(
        s5_regOut[39]), .QN() );
  DFF_X1 s5_regOut_reg_1__2__0_ ( .D(s5_refreshed[40]), .CK(clk), .Q(
        s5_regOut[40]), .QN() );
  DFF_X1 s5_regOut_reg_1__2__1_ ( .D(s5_refreshed[41]), .CK(clk), .Q(
        s5_regOut[41]), .QN() );
  DFF_X1 s5_regOut_reg_1__2__2_ ( .D(s5_refreshed[42]), .CK(clk), .Q(
        s5_regOut[42]), .QN() );
  DFF_X1 s5_regOut_reg_1__2__3_ ( .D(s5_refreshed[43]), .CK(clk), .Q(
        s5_regOut[43]), .QN() );
  DFF_X1 s5_regOut_reg_1__2__4_ ( .D(s5_refreshed[44]), .CK(clk), .Q(
        s5_regOut[44]), .QN() );
  DFF_X1 s5_regOut_reg_1__2__5_ ( .D(s5_refreshed[45]), .CK(clk), .Q(
        s5_regOut[45]), .QN() );
  DFF_X1 s5_regOut_reg_1__2__6_ ( .D(s5_refreshed[46]), .CK(clk), .Q(
        s5_regOut[46]), .QN() );
  DFF_X1 s5_regOut_reg_1__2__7_ ( .D(s5_refreshed[47]), .CK(clk), .Q(
        s5_regOut[47]), .QN() );
  DFF_X1 s5_regOut_reg_2__0__0_ ( .D(s5_refreshed[48]), .CK(clk), .Q(
        s5_regOut[48]), .QN() );
  DFF_X1 s5_regOut_reg_2__0__1_ ( .D(s5_refreshed[49]), .CK(clk), .Q(
        s5_regOut[49]), .QN() );
  DFF_X1 s5_regOut_reg_2__0__2_ ( .D(s5_refreshed[50]), .CK(clk), .Q(
        s5_regOut[50]), .QN() );
  DFF_X1 s5_regOut_reg_2__0__3_ ( .D(s5_refreshed[51]), .CK(clk), .Q(
        s5_regOut[51]), .QN() );
  DFF_X1 s5_regOut_reg_2__0__4_ ( .D(s5_refreshed[52]), .CK(clk), .Q(
        s5_regOut[52]), .QN() );
  DFF_X1 s5_regOut_reg_2__0__5_ ( .D(s5_refreshed[53]), .CK(clk), .Q(
        s5_regOut[53]), .QN() );
  DFF_X1 s5_regOut_reg_2__0__6_ ( .D(s5_refreshed[54]), .CK(clk), .Q(
        s5_regOut[54]), .QN() );
  DFF_X1 s5_regOut_reg_2__0__7_ ( .D(s5_refreshed[55]), .CK(clk), .Q(
        s5_regOut[55]), .QN() );
  DFF_X1 s5_regOut_reg_2__1__0_ ( .D(s5_refreshed[56]), .CK(clk), .Q(
        s5_regOut[56]), .QN() );
  DFF_X1 s5_regOut_reg_2__1__1_ ( .D(s5_refreshed[57]), .CK(clk), .Q(
        s5_regOut[57]), .QN() );
  DFF_X1 s5_regOut_reg_2__1__2_ ( .D(s5_refreshed[58]), .CK(clk), .Q(
        s5_regOut[58]), .QN() );
  DFF_X1 s5_regOut_reg_2__1__3_ ( .D(s5_refreshed[59]), .CK(clk), .Q(
        s5_regOut[59]), .QN() );
  DFF_X1 s5_regOut_reg_2__1__4_ ( .D(s5_refreshed[60]), .CK(clk), .Q(
        s5_regOut[60]), .QN() );
  DFF_X1 s5_regOut_reg_2__1__5_ ( .D(s5_refreshed[61]), .CK(clk), .Q(
        s5_regOut[61]), .QN() );
  DFF_X1 s5_regOut_reg_2__1__6_ ( .D(s5_refreshed[62]), .CK(clk), .Q(
        s5_regOut[62]), .QN() );
  DFF_X1 s5_regOut_reg_2__1__7_ ( .D(s5_refreshed[63]), .CK(clk), .Q(
        s5_regOut[63]), .QN() );
  DFF_X1 s5_regOut_reg_2__2__0_ ( .D(s5_refreshed[64]), .CK(clk), .Q(
        s5_regOut[64]), .QN() );
  DFF_X1 s5_regOut_reg_2__2__1_ ( .D(s5_refreshed[65]), .CK(clk), .Q(
        s5_regOut[65]), .QN() );
  DFF_X1 s5_regOut_reg_2__2__2_ ( .D(s5_refreshed[66]), .CK(clk), .Q(
        s5_regOut[66]), .QN() );
  DFF_X1 s5_regOut_reg_2__2__3_ ( .D(s5_refreshed[67]), .CK(clk), .Q(
        s5_regOut[67]), .QN() );
  DFF_X1 s5_regOut_reg_2__2__4_ ( .D(s5_refreshed[68]), .CK(clk), .Q(
        s5_regOut[68]), .QN() );
  DFF_X1 s5_regOut_reg_2__2__5_ ( .D(s5_refreshed[69]), .CK(clk), .Q(
        s5_regOut[69]), .QN() );
  DFF_X1 s5_regOut_reg_2__2__6_ ( .D(s5_refreshed[70]), .CK(clk), .Q(
        s5_regOut[70]), .QN() );
  DFF_X1 s5_regOut_reg_2__2__7_ ( .D(s5_refreshed[71]), .CK(clk), .Q(
        s5_regOut[71]), .QN() );
  XNOR2_X1 s5_mul1_2_2_U28 ( .A(s5_mul1_2_2_n76), .B(s5_mul1_2_2_n75), .ZN(
        s5_concat[67]) );
  NAND2_X1 s5_mul1_2_2_U27 ( .A1(s5_n12), .A2(stage4Out[35]), .ZN(
        s5_mul1_2_2_n75) );
  XOR2_X1 s5_mul1_2_2_U26 ( .A(s5_mul1_2_2_n74), .B(s5_mul1_2_2_n73), .Z(
        s5_mul1_2_2_n76) );
  XNOR2_X1 s5_mul1_2_2_U25 ( .A(s5_mul1_2_2_n72), .B(s5_mul1_2_2_n71), .ZN(
        s5_concat[66]) );
  NAND2_X1 s5_mul1_2_2_U24 ( .A1(stage4Out[34]), .A2(s5_n11), .ZN(
        s5_mul1_2_2_n71) );
  XOR2_X1 s5_mul1_2_2_U23 ( .A(s5_mul1_2_2_n73), .B(s5_mul1_2_2_n70), .Z(
        s5_mul1_2_2_n72) );
  AOI221_X1 s5_mul1_2_2_U22 ( .B1(s5_n11), .B2(s5_n12), .C1(stage4Out[34]), 
        .C2(stage4Out[35]), .A(s5_mul1_2_2_n69), .ZN(s5_mul1_2_2_n73) );
  OAI22_X1 s5_mul1_2_2_U21 ( .A1(s5_n11), .A2(s5_n12), .B1(stage4Out[35]), 
        .B2(stage4Out[34]), .ZN(s5_mul1_2_2_n69) );
  XNOR2_X1 s5_mul1_2_2_U20 ( .A(s5_mul1_2_2_n68), .B(s5_mul1_2_2_n67), .ZN(
        s5_concat[65]) );
  NAND2_X1 s5_mul1_2_2_U19 ( .A1(s5_n10), .A2(stage4Out[33]), .ZN(
        s5_mul1_2_2_n67) );
  XOR2_X1 s5_mul1_2_2_U18 ( .A(s5_mul1_2_2_n74), .B(s5_mul1_2_2_n66), .Z(
        s5_mul1_2_2_n68) );
  OAI22_X1 s5_mul1_2_2_U17 ( .A1(s5_mul1_2_2_n65), .A2(s5_mul1_2_2_n64), .B1(
        s5_mul1_2_2_n63), .B2(s5_mul1_2_2_n62), .ZN(s5_mul1_2_2_n74) );
  NAND2_X1 s5_mul1_2_2_U16 ( .A1(s5_mul1_2_2_n61), .A2(s5_mul1_2_2_n65), .ZN(
        s5_mul1_2_2_n62) );
  XNOR2_X1 s5_mul1_2_2_U15 ( .A(s5_mul1_2_2_n60), .B(s5_mul1_2_2_n59), .ZN(
        s5_mul1_2_2_n64) );
  NAND2_X1 s5_mul1_2_2_U14 ( .A1(s5_mul1_2_2_n61), .A2(s5_mul1_2_2_n63), .ZN(
        s5_mul1_2_2_n59) );
  INV_X1 s5_mul1_2_2_U13 ( .A(s5_mul1_2_2_n58), .ZN(s5_mul1_2_2_n65) );
  XNOR2_X1 s5_mul1_2_2_U12 ( .A(s5_mul1_2_2_n57), .B(s5_mul1_2_2_n56), .ZN(
        s5_concat[64]) );
  NAND2_X1 s5_mul1_2_2_U11 ( .A1(stage4Out[32]), .A2(s5_n9), .ZN(
        s5_mul1_2_2_n56) );
  XOR2_X1 s5_mul1_2_2_U10 ( .A(s5_mul1_2_2_n66), .B(s5_mul1_2_2_n70), .Z(
        s5_mul1_2_2_n57) );
  XNOR2_X1 s5_mul1_2_2_U9 ( .A(s5_mul1_2_2_n55), .B(s5_mul1_2_2_n54), .ZN(
        s5_mul1_2_2_n70) );
  NAND2_X1 s5_mul1_2_2_U8 ( .A1(s5_mul1_2_2_n61), .A2(s5_mul1_2_2_n58), .ZN(
        s5_mul1_2_2_n54) );
  XOR2_X1 s5_mul1_2_2_U7 ( .A(s5_n10), .B(s5_n12), .Z(s5_mul1_2_2_n58) );
  XOR2_X1 s5_mul1_2_2_U6 ( .A(stage4Out[33]), .B(stage4Out[35]), .Z(
        s5_mul1_2_2_n61) );
  NOR2_X1 s5_mul1_2_2_U5 ( .A1(s5_mul1_2_2_n63), .A2(s5_mul1_2_2_n60), .ZN(
        s5_mul1_2_2_n55) );
  XNOR2_X1 s5_mul1_2_2_U4 ( .A(stage4Out[32]), .B(stage4Out[34]), .ZN(
        s5_mul1_2_2_n60) );
  XNOR2_X1 s5_mul1_2_2_U3 ( .A(s5_n9), .B(s5_n11), .ZN(s5_mul1_2_2_n63) );
  AOI221_X1 s5_mul1_2_2_U2 ( .B1(s5_n9), .B2(s5_n10), .C1(stage4Out[32]), .C2(
        stage4Out[33]), .A(s5_mul1_2_2_n53), .ZN(s5_mul1_2_2_n66) );
  OAI22_X1 s5_mul1_2_2_U1 ( .A1(s5_n9), .A2(s5_n10), .B1(stage4Out[33]), .B2(
        stage4Out[32]), .ZN(s5_mul1_2_2_n53) );
  XNOR2_X1 s5_mul1_2_1_U28 ( .A(s5_mul1_2_1_n76), .B(s5_mul1_2_1_n75), .ZN(
        s5_concat[59]) );
  NAND2_X1 s5_mul1_2_1_U27 ( .A1(s5_n8), .A2(stage4Out[35]), .ZN(
        s5_mul1_2_1_n75) );
  XOR2_X1 s5_mul1_2_1_U26 ( .A(s5_mul1_2_1_n74), .B(s5_mul1_2_1_n73), .Z(
        s5_mul1_2_1_n76) );
  XNOR2_X1 s5_mul1_2_1_U25 ( .A(s5_mul1_2_1_n72), .B(s5_mul1_2_1_n71), .ZN(
        s5_concat[58]) );
  NAND2_X1 s5_mul1_2_1_U24 ( .A1(stage4Out[34]), .A2(s5_n7), .ZN(
        s5_mul1_2_1_n71) );
  XOR2_X1 s5_mul1_2_1_U23 ( .A(s5_mul1_2_1_n73), .B(s5_mul1_2_1_n70), .Z(
        s5_mul1_2_1_n72) );
  AOI221_X1 s5_mul1_2_1_U22 ( .B1(s5_n7), .B2(s5_n8), .C1(stage4Out[34]), .C2(
        stage4Out[35]), .A(s5_mul1_2_1_n69), .ZN(s5_mul1_2_1_n73) );
  OAI22_X1 s5_mul1_2_1_U21 ( .A1(s5_n7), .A2(s5_n8), .B1(stage4Out[35]), .B2(
        stage4Out[34]), .ZN(s5_mul1_2_1_n69) );
  XNOR2_X1 s5_mul1_2_1_U20 ( .A(s5_mul1_2_1_n68), .B(s5_mul1_2_1_n67), .ZN(
        s5_concat[57]) );
  NAND2_X1 s5_mul1_2_1_U19 ( .A1(s5_n6), .A2(stage4Out[33]), .ZN(
        s5_mul1_2_1_n67) );
  XOR2_X1 s5_mul1_2_1_U18 ( .A(s5_mul1_2_1_n74), .B(s5_mul1_2_1_n66), .Z(
        s5_mul1_2_1_n68) );
  OAI22_X1 s5_mul1_2_1_U17 ( .A1(s5_mul1_2_1_n65), .A2(s5_mul1_2_1_n64), .B1(
        s5_mul1_2_1_n63), .B2(s5_mul1_2_1_n62), .ZN(s5_mul1_2_1_n74) );
  NAND2_X1 s5_mul1_2_1_U16 ( .A1(s5_mul1_2_1_n61), .A2(s5_mul1_2_1_n65), .ZN(
        s5_mul1_2_1_n62) );
  XNOR2_X1 s5_mul1_2_1_U15 ( .A(s5_mul1_2_1_n60), .B(s5_mul1_2_1_n59), .ZN(
        s5_mul1_2_1_n64) );
  NAND2_X1 s5_mul1_2_1_U14 ( .A1(s5_mul1_2_1_n61), .A2(s5_mul1_2_1_n63), .ZN(
        s5_mul1_2_1_n59) );
  INV_X1 s5_mul1_2_1_U13 ( .A(s5_mul1_2_1_n58), .ZN(s5_mul1_2_1_n65) );
  XNOR2_X1 s5_mul1_2_1_U12 ( .A(s5_mul1_2_1_n57), .B(s5_mul1_2_1_n56), .ZN(
        s5_concat[56]) );
  NAND2_X1 s5_mul1_2_1_U11 ( .A1(stage4Out[32]), .A2(s5_n5), .ZN(
        s5_mul1_2_1_n56) );
  XOR2_X1 s5_mul1_2_1_U10 ( .A(s5_mul1_2_1_n66), .B(s5_mul1_2_1_n70), .Z(
        s5_mul1_2_1_n57) );
  XNOR2_X1 s5_mul1_2_1_U9 ( .A(s5_mul1_2_1_n55), .B(s5_mul1_2_1_n54), .ZN(
        s5_mul1_2_1_n70) );
  NAND2_X1 s5_mul1_2_1_U8 ( .A1(s5_mul1_2_1_n61), .A2(s5_mul1_2_1_n58), .ZN(
        s5_mul1_2_1_n54) );
  XOR2_X1 s5_mul1_2_1_U7 ( .A(s5_n6), .B(s5_n8), .Z(s5_mul1_2_1_n58) );
  XOR2_X1 s5_mul1_2_1_U6 ( .A(stage4Out[33]), .B(stage4Out[35]), .Z(
        s5_mul1_2_1_n61) );
  NOR2_X1 s5_mul1_2_1_U5 ( .A1(s5_mul1_2_1_n63), .A2(s5_mul1_2_1_n60), .ZN(
        s5_mul1_2_1_n55) );
  XNOR2_X1 s5_mul1_2_1_U4 ( .A(stage4Out[32]), .B(stage4Out[34]), .ZN(
        s5_mul1_2_1_n60) );
  XNOR2_X1 s5_mul1_2_1_U3 ( .A(s5_n5), .B(s5_n7), .ZN(s5_mul1_2_1_n63) );
  AOI221_X1 s5_mul1_2_1_U2 ( .B1(s5_n5), .B2(s5_n6), .C1(stage4Out[32]), .C2(
        stage4Out[33]), .A(s5_mul1_2_1_n53), .ZN(s5_mul1_2_1_n66) );
  OAI22_X1 s5_mul1_2_1_U1 ( .A1(s5_n5), .A2(s5_n6), .B1(stage4Out[33]), .B2(
        stage4Out[32]), .ZN(s5_mul1_2_1_n53) );
  XNOR2_X1 s5_mul1_2_0_U28 ( .A(s5_mul1_2_0_n76), .B(s5_mul1_2_0_n75), .ZN(
        s5_concat[51]) );
  NAND2_X1 s5_mul1_2_0_U27 ( .A1(s5_n4), .A2(stage4Out[35]), .ZN(
        s5_mul1_2_0_n75) );
  XOR2_X1 s5_mul1_2_0_U26 ( .A(s5_mul1_2_0_n74), .B(s5_mul1_2_0_n73), .Z(
        s5_mul1_2_0_n76) );
  XNOR2_X1 s5_mul1_2_0_U25 ( .A(s5_mul1_2_0_n72), .B(s5_mul1_2_0_n71), .ZN(
        s5_concat[50]) );
  NAND2_X1 s5_mul1_2_0_U24 ( .A1(stage4Out[34]), .A2(s5_n3), .ZN(
        s5_mul1_2_0_n71) );
  XOR2_X1 s5_mul1_2_0_U23 ( .A(s5_mul1_2_0_n73), .B(s5_mul1_2_0_n70), .Z(
        s5_mul1_2_0_n72) );
  AOI221_X1 s5_mul1_2_0_U22 ( .B1(s5_n3), .B2(s5_n4), .C1(stage4Out[34]), .C2(
        stage4Out[35]), .A(s5_mul1_2_0_n69), .ZN(s5_mul1_2_0_n73) );
  OAI22_X1 s5_mul1_2_0_U21 ( .A1(s5_n3), .A2(s5_n4), .B1(stage4Out[35]), .B2(
        stage4Out[34]), .ZN(s5_mul1_2_0_n69) );
  XNOR2_X1 s5_mul1_2_0_U20 ( .A(s5_mul1_2_0_n68), .B(s5_mul1_2_0_n67), .ZN(
        s5_concat[49]) );
  NAND2_X1 s5_mul1_2_0_U19 ( .A1(s5_n2), .A2(stage4Out[33]), .ZN(
        s5_mul1_2_0_n67) );
  XOR2_X1 s5_mul1_2_0_U18 ( .A(s5_mul1_2_0_n74), .B(s5_mul1_2_0_n66), .Z(
        s5_mul1_2_0_n68) );
  OAI22_X1 s5_mul1_2_0_U17 ( .A1(s5_mul1_2_0_n65), .A2(s5_mul1_2_0_n64), .B1(
        s5_mul1_2_0_n63), .B2(s5_mul1_2_0_n62), .ZN(s5_mul1_2_0_n74) );
  NAND2_X1 s5_mul1_2_0_U16 ( .A1(s5_mul1_2_0_n61), .A2(s5_mul1_2_0_n65), .ZN(
        s5_mul1_2_0_n62) );
  XNOR2_X1 s5_mul1_2_0_U15 ( .A(s5_mul1_2_0_n60), .B(s5_mul1_2_0_n59), .ZN(
        s5_mul1_2_0_n64) );
  NAND2_X1 s5_mul1_2_0_U14 ( .A1(s5_mul1_2_0_n61), .A2(s5_mul1_2_0_n63), .ZN(
        s5_mul1_2_0_n59) );
  INV_X1 s5_mul1_2_0_U13 ( .A(s5_mul1_2_0_n58), .ZN(s5_mul1_2_0_n65) );
  XNOR2_X1 s5_mul1_2_0_U12 ( .A(s5_mul1_2_0_n57), .B(s5_mul1_2_0_n56), .ZN(
        s5_concat[48]) );
  NAND2_X1 s5_mul1_2_0_U11 ( .A1(stage4Out[32]), .A2(s5_n1), .ZN(
        s5_mul1_2_0_n56) );
  XOR2_X1 s5_mul1_2_0_U10 ( .A(s5_mul1_2_0_n66), .B(s5_mul1_2_0_n70), .Z(
        s5_mul1_2_0_n57) );
  XNOR2_X1 s5_mul1_2_0_U9 ( .A(s5_mul1_2_0_n55), .B(s5_mul1_2_0_n54), .ZN(
        s5_mul1_2_0_n70) );
  NAND2_X1 s5_mul1_2_0_U8 ( .A1(s5_mul1_2_0_n61), .A2(s5_mul1_2_0_n58), .ZN(
        s5_mul1_2_0_n54) );
  XOR2_X1 s5_mul1_2_0_U7 ( .A(s5_n2), .B(s5_n4), .Z(s5_mul1_2_0_n58) );
  XOR2_X1 s5_mul1_2_0_U6 ( .A(stage4Out[33]), .B(stage4Out[35]), .Z(
        s5_mul1_2_0_n61) );
  NOR2_X1 s5_mul1_2_0_U5 ( .A1(s5_mul1_2_0_n63), .A2(s5_mul1_2_0_n60), .ZN(
        s5_mul1_2_0_n55) );
  XNOR2_X1 s5_mul1_2_0_U4 ( .A(stage4Out[32]), .B(stage4Out[34]), .ZN(
        s5_mul1_2_0_n60) );
  XNOR2_X1 s5_mul1_2_0_U3 ( .A(s5_n1), .B(s5_n3), .ZN(s5_mul1_2_0_n63) );
  AOI221_X1 s5_mul1_2_0_U2 ( .B1(s5_n1), .B2(s5_n2), .C1(stage4Out[32]), .C2(
        stage4Out[33]), .A(s5_mul1_2_0_n53), .ZN(s5_mul1_2_0_n66) );
  OAI22_X1 s5_mul1_2_0_U1 ( .A1(s5_n1), .A2(s5_n2), .B1(stage4Out[33]), .B2(
        stage4Out[32]), .ZN(s5_mul1_2_0_n53) );
  XNOR2_X1 s5_mul1_1_2_U28 ( .A(s5_mul1_1_2_n76), .B(s5_mul1_1_2_n75), .ZN(
        s5_concat[43]) );
  NAND2_X1 s5_mul1_1_2_U27 ( .A1(s5_n12), .A2(stage4Out[23]), .ZN(
        s5_mul1_1_2_n75) );
  XOR2_X1 s5_mul1_1_2_U26 ( .A(s5_mul1_1_2_n74), .B(s5_mul1_1_2_n73), .Z(
        s5_mul1_1_2_n76) );
  XNOR2_X1 s5_mul1_1_2_U25 ( .A(s5_mul1_1_2_n72), .B(s5_mul1_1_2_n71), .ZN(
        s5_concat[42]) );
  NAND2_X1 s5_mul1_1_2_U24 ( .A1(stage4Out[22]), .A2(s5_n11), .ZN(
        s5_mul1_1_2_n71) );
  XOR2_X1 s5_mul1_1_2_U23 ( .A(s5_mul1_1_2_n73), .B(s5_mul1_1_2_n70), .Z(
        s5_mul1_1_2_n72) );
  AOI221_X1 s5_mul1_1_2_U22 ( .B1(s5_n11), .B2(s5_n12), .C1(stage4Out[22]), 
        .C2(stage4Out[23]), .A(s5_mul1_1_2_n69), .ZN(s5_mul1_1_2_n73) );
  OAI22_X1 s5_mul1_1_2_U21 ( .A1(s5_n11), .A2(s5_n12), .B1(stage4Out[23]), 
        .B2(stage4Out[22]), .ZN(s5_mul1_1_2_n69) );
  XNOR2_X1 s5_mul1_1_2_U20 ( .A(s5_mul1_1_2_n68), .B(s5_mul1_1_2_n67), .ZN(
        s5_concat[41]) );
  NAND2_X1 s5_mul1_1_2_U19 ( .A1(s5_n10), .A2(stage4Out[21]), .ZN(
        s5_mul1_1_2_n67) );
  XOR2_X1 s5_mul1_1_2_U18 ( .A(s5_mul1_1_2_n74), .B(s5_mul1_1_2_n66), .Z(
        s5_mul1_1_2_n68) );
  OAI22_X1 s5_mul1_1_2_U17 ( .A1(s5_mul1_1_2_n65), .A2(s5_mul1_1_2_n64), .B1(
        s5_mul1_1_2_n63), .B2(s5_mul1_1_2_n62), .ZN(s5_mul1_1_2_n74) );
  NAND2_X1 s5_mul1_1_2_U16 ( .A1(s5_mul1_1_2_n61), .A2(s5_mul1_1_2_n65), .ZN(
        s5_mul1_1_2_n62) );
  XNOR2_X1 s5_mul1_1_2_U15 ( .A(s5_mul1_1_2_n60), .B(s5_mul1_1_2_n59), .ZN(
        s5_mul1_1_2_n64) );
  NAND2_X1 s5_mul1_1_2_U14 ( .A1(s5_mul1_1_2_n61), .A2(s5_mul1_1_2_n63), .ZN(
        s5_mul1_1_2_n59) );
  INV_X1 s5_mul1_1_2_U13 ( .A(s5_mul1_1_2_n58), .ZN(s5_mul1_1_2_n65) );
  XNOR2_X1 s5_mul1_1_2_U12 ( .A(s5_mul1_1_2_n57), .B(s5_mul1_1_2_n56), .ZN(
        s5_concat[40]) );
  NAND2_X1 s5_mul1_1_2_U11 ( .A1(stage4Out[20]), .A2(s5_n9), .ZN(
        s5_mul1_1_2_n56) );
  XOR2_X1 s5_mul1_1_2_U10 ( .A(s5_mul1_1_2_n66), .B(s5_mul1_1_2_n70), .Z(
        s5_mul1_1_2_n57) );
  XNOR2_X1 s5_mul1_1_2_U9 ( .A(s5_mul1_1_2_n55), .B(s5_mul1_1_2_n54), .ZN(
        s5_mul1_1_2_n70) );
  NAND2_X1 s5_mul1_1_2_U8 ( .A1(s5_mul1_1_2_n61), .A2(s5_mul1_1_2_n58), .ZN(
        s5_mul1_1_2_n54) );
  XOR2_X1 s5_mul1_1_2_U7 ( .A(s5_n10), .B(s5_n12), .Z(s5_mul1_1_2_n58) );
  XOR2_X1 s5_mul1_1_2_U6 ( .A(stage4Out[21]), .B(stage4Out[23]), .Z(
        s5_mul1_1_2_n61) );
  NOR2_X1 s5_mul1_1_2_U5 ( .A1(s5_mul1_1_2_n63), .A2(s5_mul1_1_2_n60), .ZN(
        s5_mul1_1_2_n55) );
  XNOR2_X1 s5_mul1_1_2_U4 ( .A(stage4Out[20]), .B(stage4Out[22]), .ZN(
        s5_mul1_1_2_n60) );
  XNOR2_X1 s5_mul1_1_2_U3 ( .A(s5_n9), .B(s5_n11), .ZN(s5_mul1_1_2_n63) );
  AOI221_X1 s5_mul1_1_2_U2 ( .B1(s5_n9), .B2(s5_n10), .C1(stage4Out[20]), .C2(
        stage4Out[21]), .A(s5_mul1_1_2_n53), .ZN(s5_mul1_1_2_n66) );
  OAI22_X1 s5_mul1_1_2_U1 ( .A1(s5_n9), .A2(s5_n10), .B1(stage4Out[21]), .B2(
        stage4Out[20]), .ZN(s5_mul1_1_2_n53) );
  XNOR2_X1 s5_mul1_1_1_U28 ( .A(s5_mul1_1_1_n76), .B(s5_mul1_1_1_n75), .ZN(
        s5_concat[35]) );
  NAND2_X1 s5_mul1_1_1_U27 ( .A1(s5_n8), .A2(stage4Out[23]), .ZN(
        s5_mul1_1_1_n75) );
  XOR2_X1 s5_mul1_1_1_U26 ( .A(s5_mul1_1_1_n74), .B(s5_mul1_1_1_n73), .Z(
        s5_mul1_1_1_n76) );
  XNOR2_X1 s5_mul1_1_1_U25 ( .A(s5_mul1_1_1_n72), .B(s5_mul1_1_1_n71), .ZN(
        s5_concat[34]) );
  NAND2_X1 s5_mul1_1_1_U24 ( .A1(stage4Out[22]), .A2(s5_n7), .ZN(
        s5_mul1_1_1_n71) );
  XOR2_X1 s5_mul1_1_1_U23 ( .A(s5_mul1_1_1_n73), .B(s5_mul1_1_1_n70), .Z(
        s5_mul1_1_1_n72) );
  AOI221_X1 s5_mul1_1_1_U22 ( .B1(s5_n7), .B2(s5_n8), .C1(stage4Out[22]), .C2(
        stage4Out[23]), .A(s5_mul1_1_1_n69), .ZN(s5_mul1_1_1_n73) );
  OAI22_X1 s5_mul1_1_1_U21 ( .A1(s5_n7), .A2(s5_n8), .B1(stage4Out[23]), .B2(
        stage4Out[22]), .ZN(s5_mul1_1_1_n69) );
  XNOR2_X1 s5_mul1_1_1_U20 ( .A(s5_mul1_1_1_n68), .B(s5_mul1_1_1_n67), .ZN(
        s5_concat[33]) );
  NAND2_X1 s5_mul1_1_1_U19 ( .A1(s5_n6), .A2(stage4Out[21]), .ZN(
        s5_mul1_1_1_n67) );
  XOR2_X1 s5_mul1_1_1_U18 ( .A(s5_mul1_1_1_n74), .B(s5_mul1_1_1_n66), .Z(
        s5_mul1_1_1_n68) );
  OAI22_X1 s5_mul1_1_1_U17 ( .A1(s5_mul1_1_1_n65), .A2(s5_mul1_1_1_n64), .B1(
        s5_mul1_1_1_n63), .B2(s5_mul1_1_1_n62), .ZN(s5_mul1_1_1_n74) );
  NAND2_X1 s5_mul1_1_1_U16 ( .A1(s5_mul1_1_1_n61), .A2(s5_mul1_1_1_n65), .ZN(
        s5_mul1_1_1_n62) );
  XNOR2_X1 s5_mul1_1_1_U15 ( .A(s5_mul1_1_1_n60), .B(s5_mul1_1_1_n59), .ZN(
        s5_mul1_1_1_n64) );
  NAND2_X1 s5_mul1_1_1_U14 ( .A1(s5_mul1_1_1_n61), .A2(s5_mul1_1_1_n63), .ZN(
        s5_mul1_1_1_n59) );
  INV_X1 s5_mul1_1_1_U13 ( .A(s5_mul1_1_1_n58), .ZN(s5_mul1_1_1_n65) );
  XNOR2_X1 s5_mul1_1_1_U12 ( .A(s5_mul1_1_1_n57), .B(s5_mul1_1_1_n56), .ZN(
        s5_concat[32]) );
  NAND2_X1 s5_mul1_1_1_U11 ( .A1(stage4Out[20]), .A2(s5_n5), .ZN(
        s5_mul1_1_1_n56) );
  XOR2_X1 s5_mul1_1_1_U10 ( .A(s5_mul1_1_1_n66), .B(s5_mul1_1_1_n70), .Z(
        s5_mul1_1_1_n57) );
  XNOR2_X1 s5_mul1_1_1_U9 ( .A(s5_mul1_1_1_n55), .B(s5_mul1_1_1_n54), .ZN(
        s5_mul1_1_1_n70) );
  NAND2_X1 s5_mul1_1_1_U8 ( .A1(s5_mul1_1_1_n61), .A2(s5_mul1_1_1_n58), .ZN(
        s5_mul1_1_1_n54) );
  XOR2_X1 s5_mul1_1_1_U7 ( .A(s5_n6), .B(s5_n8), .Z(s5_mul1_1_1_n58) );
  XOR2_X1 s5_mul1_1_1_U6 ( .A(stage4Out[21]), .B(stage4Out[23]), .Z(
        s5_mul1_1_1_n61) );
  NOR2_X1 s5_mul1_1_1_U5 ( .A1(s5_mul1_1_1_n63), .A2(s5_mul1_1_1_n60), .ZN(
        s5_mul1_1_1_n55) );
  XNOR2_X1 s5_mul1_1_1_U4 ( .A(stage4Out[20]), .B(stage4Out[22]), .ZN(
        s5_mul1_1_1_n60) );
  XNOR2_X1 s5_mul1_1_1_U3 ( .A(s5_n5), .B(s5_n7), .ZN(s5_mul1_1_1_n63) );
  AOI221_X1 s5_mul1_1_1_U2 ( .B1(s5_n5), .B2(s5_n6), .C1(stage4Out[20]), .C2(
        stage4Out[21]), .A(s5_mul1_1_1_n53), .ZN(s5_mul1_1_1_n66) );
  OAI22_X1 s5_mul1_1_1_U1 ( .A1(s5_n5), .A2(s5_n6), .B1(stage4Out[21]), .B2(
        stage4Out[20]), .ZN(s5_mul1_1_1_n53) );
  XNOR2_X1 s5_mul1_1_0_U28 ( .A(s5_mul1_1_0_n76), .B(s5_mul1_1_0_n75), .ZN(
        s5_concat[27]) );
  NAND2_X1 s5_mul1_1_0_U27 ( .A1(s5_n4), .A2(stage4Out[23]), .ZN(
        s5_mul1_1_0_n75) );
  XOR2_X1 s5_mul1_1_0_U26 ( .A(s5_mul1_1_0_n74), .B(s5_mul1_1_0_n73), .Z(
        s5_mul1_1_0_n76) );
  XNOR2_X1 s5_mul1_1_0_U25 ( .A(s5_mul1_1_0_n72), .B(s5_mul1_1_0_n71), .ZN(
        s5_concat[26]) );
  NAND2_X1 s5_mul1_1_0_U24 ( .A1(stage4Out[22]), .A2(s5_n3), .ZN(
        s5_mul1_1_0_n71) );
  XOR2_X1 s5_mul1_1_0_U23 ( .A(s5_mul1_1_0_n73), .B(s5_mul1_1_0_n70), .Z(
        s5_mul1_1_0_n72) );
  AOI221_X1 s5_mul1_1_0_U22 ( .B1(s5_n3), .B2(s5_n4), .C1(stage4Out[22]), .C2(
        stage4Out[23]), .A(s5_mul1_1_0_n69), .ZN(s5_mul1_1_0_n73) );
  OAI22_X1 s5_mul1_1_0_U21 ( .A1(s5_n3), .A2(s5_n4), .B1(stage4Out[23]), .B2(
        stage4Out[22]), .ZN(s5_mul1_1_0_n69) );
  XNOR2_X1 s5_mul1_1_0_U20 ( .A(s5_mul1_1_0_n68), .B(s5_mul1_1_0_n67), .ZN(
        s5_concat[25]) );
  NAND2_X1 s5_mul1_1_0_U19 ( .A1(s5_n2), .A2(stage4Out[21]), .ZN(
        s5_mul1_1_0_n67) );
  XOR2_X1 s5_mul1_1_0_U18 ( .A(s5_mul1_1_0_n74), .B(s5_mul1_1_0_n66), .Z(
        s5_mul1_1_0_n68) );
  OAI22_X1 s5_mul1_1_0_U17 ( .A1(s5_mul1_1_0_n65), .A2(s5_mul1_1_0_n64), .B1(
        s5_mul1_1_0_n63), .B2(s5_mul1_1_0_n62), .ZN(s5_mul1_1_0_n74) );
  NAND2_X1 s5_mul1_1_0_U16 ( .A1(s5_mul1_1_0_n61), .A2(s5_mul1_1_0_n65), .ZN(
        s5_mul1_1_0_n62) );
  XNOR2_X1 s5_mul1_1_0_U15 ( .A(s5_mul1_1_0_n60), .B(s5_mul1_1_0_n59), .ZN(
        s5_mul1_1_0_n64) );
  NAND2_X1 s5_mul1_1_0_U14 ( .A1(s5_mul1_1_0_n61), .A2(s5_mul1_1_0_n63), .ZN(
        s5_mul1_1_0_n59) );
  INV_X1 s5_mul1_1_0_U13 ( .A(s5_mul1_1_0_n58), .ZN(s5_mul1_1_0_n65) );
  XNOR2_X1 s5_mul1_1_0_U12 ( .A(s5_mul1_1_0_n57), .B(s5_mul1_1_0_n56), .ZN(
        s5_concat[24]) );
  NAND2_X1 s5_mul1_1_0_U11 ( .A1(stage4Out[20]), .A2(s5_n1), .ZN(
        s5_mul1_1_0_n56) );
  XOR2_X1 s5_mul1_1_0_U10 ( .A(s5_mul1_1_0_n66), .B(s5_mul1_1_0_n70), .Z(
        s5_mul1_1_0_n57) );
  XNOR2_X1 s5_mul1_1_0_U9 ( .A(s5_mul1_1_0_n55), .B(s5_mul1_1_0_n54), .ZN(
        s5_mul1_1_0_n70) );
  NAND2_X1 s5_mul1_1_0_U8 ( .A1(s5_mul1_1_0_n61), .A2(s5_mul1_1_0_n58), .ZN(
        s5_mul1_1_0_n54) );
  XOR2_X1 s5_mul1_1_0_U7 ( .A(s5_n2), .B(s5_n4), .Z(s5_mul1_1_0_n58) );
  XOR2_X1 s5_mul1_1_0_U6 ( .A(stage4Out[21]), .B(stage4Out[23]), .Z(
        s5_mul1_1_0_n61) );
  NOR2_X1 s5_mul1_1_0_U5 ( .A1(s5_mul1_1_0_n63), .A2(s5_mul1_1_0_n60), .ZN(
        s5_mul1_1_0_n55) );
  XNOR2_X1 s5_mul1_1_0_U4 ( .A(stage4Out[20]), .B(stage4Out[22]), .ZN(
        s5_mul1_1_0_n60) );
  XNOR2_X1 s5_mul1_1_0_U3 ( .A(s5_n1), .B(s5_n3), .ZN(s5_mul1_1_0_n63) );
  AOI221_X1 s5_mul1_1_0_U2 ( .B1(s5_n1), .B2(s5_n2), .C1(stage4Out[20]), .C2(
        stage4Out[21]), .A(s5_mul1_1_0_n53), .ZN(s5_mul1_1_0_n66) );
  OAI22_X1 s5_mul1_1_0_U1 ( .A1(s5_n1), .A2(s5_n2), .B1(stage4Out[21]), .B2(
        stage4Out[20]), .ZN(s5_mul1_1_0_n53) );
  XNOR2_X1 s5_mul1_0_2_U28 ( .A(s5_mul1_0_2_n76), .B(s5_mul1_0_2_n75), .ZN(
        s5_concat[19]) );
  NAND2_X1 s5_mul1_0_2_U27 ( .A1(s5_n12), .A2(stage4Out[11]), .ZN(
        s5_mul1_0_2_n75) );
  XOR2_X1 s5_mul1_0_2_U26 ( .A(s5_mul1_0_2_n74), .B(s5_mul1_0_2_n73), .Z(
        s5_mul1_0_2_n76) );
  XNOR2_X1 s5_mul1_0_2_U25 ( .A(s5_mul1_0_2_n72), .B(s5_mul1_0_2_n71), .ZN(
        s5_concat[18]) );
  NAND2_X1 s5_mul1_0_2_U24 ( .A1(stage4Out[10]), .A2(s5_n11), .ZN(
        s5_mul1_0_2_n71) );
  XOR2_X1 s5_mul1_0_2_U23 ( .A(s5_mul1_0_2_n73), .B(s5_mul1_0_2_n70), .Z(
        s5_mul1_0_2_n72) );
  AOI221_X1 s5_mul1_0_2_U22 ( .B1(s5_n11), .B2(s5_n12), .C1(stage4Out[10]), 
        .C2(stage4Out[11]), .A(s5_mul1_0_2_n69), .ZN(s5_mul1_0_2_n73) );
  OAI22_X1 s5_mul1_0_2_U21 ( .A1(s5_n11), .A2(s5_n12), .B1(stage4Out[11]), 
        .B2(stage4Out[10]), .ZN(s5_mul1_0_2_n69) );
  XNOR2_X1 s5_mul1_0_2_U20 ( .A(s5_mul1_0_2_n68), .B(s5_mul1_0_2_n67), .ZN(
        s5_concat[17]) );
  NAND2_X1 s5_mul1_0_2_U19 ( .A1(s5_n10), .A2(stage4Out[9]), .ZN(
        s5_mul1_0_2_n67) );
  XOR2_X1 s5_mul1_0_2_U18 ( .A(s5_mul1_0_2_n74), .B(s5_mul1_0_2_n66), .Z(
        s5_mul1_0_2_n68) );
  OAI22_X1 s5_mul1_0_2_U17 ( .A1(s5_mul1_0_2_n65), .A2(s5_mul1_0_2_n64), .B1(
        s5_mul1_0_2_n63), .B2(s5_mul1_0_2_n62), .ZN(s5_mul1_0_2_n74) );
  NAND2_X1 s5_mul1_0_2_U16 ( .A1(s5_mul1_0_2_n61), .A2(s5_mul1_0_2_n65), .ZN(
        s5_mul1_0_2_n62) );
  XNOR2_X1 s5_mul1_0_2_U15 ( .A(s5_mul1_0_2_n60), .B(s5_mul1_0_2_n59), .ZN(
        s5_mul1_0_2_n64) );
  NAND2_X1 s5_mul1_0_2_U14 ( .A1(s5_mul1_0_2_n61), .A2(s5_mul1_0_2_n63), .ZN(
        s5_mul1_0_2_n59) );
  INV_X1 s5_mul1_0_2_U13 ( .A(s5_mul1_0_2_n58), .ZN(s5_mul1_0_2_n65) );
  XNOR2_X1 s5_mul1_0_2_U12 ( .A(s5_mul1_0_2_n57), .B(s5_mul1_0_2_n56), .ZN(
        s5_concat[16]) );
  NAND2_X1 s5_mul1_0_2_U11 ( .A1(stage4Out[8]), .A2(s5_n9), .ZN(
        s5_mul1_0_2_n56) );
  XOR2_X1 s5_mul1_0_2_U10 ( .A(s5_mul1_0_2_n66), .B(s5_mul1_0_2_n70), .Z(
        s5_mul1_0_2_n57) );
  XNOR2_X1 s5_mul1_0_2_U9 ( .A(s5_mul1_0_2_n55), .B(s5_mul1_0_2_n54), .ZN(
        s5_mul1_0_2_n70) );
  NAND2_X1 s5_mul1_0_2_U8 ( .A1(s5_mul1_0_2_n61), .A2(s5_mul1_0_2_n58), .ZN(
        s5_mul1_0_2_n54) );
  XOR2_X1 s5_mul1_0_2_U7 ( .A(s5_n10), .B(s5_n12), .Z(s5_mul1_0_2_n58) );
  XOR2_X1 s5_mul1_0_2_U6 ( .A(stage4Out[9]), .B(stage4Out[11]), .Z(
        s5_mul1_0_2_n61) );
  NOR2_X1 s5_mul1_0_2_U5 ( .A1(s5_mul1_0_2_n63), .A2(s5_mul1_0_2_n60), .ZN(
        s5_mul1_0_2_n55) );
  XNOR2_X1 s5_mul1_0_2_U4 ( .A(stage4Out[8]), .B(stage4Out[10]), .ZN(
        s5_mul1_0_2_n60) );
  XNOR2_X1 s5_mul1_0_2_U3 ( .A(s5_n9), .B(s5_n11), .ZN(s5_mul1_0_2_n63) );
  AOI221_X1 s5_mul1_0_2_U2 ( .B1(s5_n9), .B2(s5_n10), .C1(stage4Out[8]), .C2(
        stage4Out[9]), .A(s5_mul1_0_2_n53), .ZN(s5_mul1_0_2_n66) );
  OAI22_X1 s5_mul1_0_2_U1 ( .A1(s5_n9), .A2(s5_n10), .B1(stage4Out[9]), .B2(
        stage4Out[8]), .ZN(s5_mul1_0_2_n53) );
  XNOR2_X1 s5_mul1_0_1_U28 ( .A(s5_mul1_0_1_n76), .B(s5_mul1_0_1_n75), .ZN(
        s5_concat[11]) );
  NAND2_X1 s5_mul1_0_1_U27 ( .A1(s5_n8), .A2(stage4Out[11]), .ZN(
        s5_mul1_0_1_n75) );
  XOR2_X1 s5_mul1_0_1_U26 ( .A(s5_mul1_0_1_n74), .B(s5_mul1_0_1_n73), .Z(
        s5_mul1_0_1_n76) );
  XNOR2_X1 s5_mul1_0_1_U25 ( .A(s5_mul1_0_1_n72), .B(s5_mul1_0_1_n71), .ZN(
        s5_concat[10]) );
  NAND2_X1 s5_mul1_0_1_U24 ( .A1(stage4Out[10]), .A2(s5_n7), .ZN(
        s5_mul1_0_1_n71) );
  XOR2_X1 s5_mul1_0_1_U23 ( .A(s5_mul1_0_1_n73), .B(s5_mul1_0_1_n70), .Z(
        s5_mul1_0_1_n72) );
  AOI221_X1 s5_mul1_0_1_U22 ( .B1(s5_n7), .B2(s5_n8), .C1(stage4Out[10]), .C2(
        stage4Out[11]), .A(s5_mul1_0_1_n69), .ZN(s5_mul1_0_1_n73) );
  OAI22_X1 s5_mul1_0_1_U21 ( .A1(s5_n7), .A2(s5_n8), .B1(stage4Out[11]), .B2(
        stage4Out[10]), .ZN(s5_mul1_0_1_n69) );
  XNOR2_X1 s5_mul1_0_1_U20 ( .A(s5_mul1_0_1_n68), .B(s5_mul1_0_1_n67), .ZN(
        s5_concat[9]) );
  NAND2_X1 s5_mul1_0_1_U19 ( .A1(s5_n6), .A2(stage4Out[9]), .ZN(
        s5_mul1_0_1_n67) );
  XOR2_X1 s5_mul1_0_1_U18 ( .A(s5_mul1_0_1_n74), .B(s5_mul1_0_1_n66), .Z(
        s5_mul1_0_1_n68) );
  OAI22_X1 s5_mul1_0_1_U17 ( .A1(s5_mul1_0_1_n65), .A2(s5_mul1_0_1_n64), .B1(
        s5_mul1_0_1_n63), .B2(s5_mul1_0_1_n62), .ZN(s5_mul1_0_1_n74) );
  NAND2_X1 s5_mul1_0_1_U16 ( .A1(s5_mul1_0_1_n61), .A2(s5_mul1_0_1_n65), .ZN(
        s5_mul1_0_1_n62) );
  XNOR2_X1 s5_mul1_0_1_U15 ( .A(s5_mul1_0_1_n60), .B(s5_mul1_0_1_n59), .ZN(
        s5_mul1_0_1_n64) );
  NAND2_X1 s5_mul1_0_1_U14 ( .A1(s5_mul1_0_1_n61), .A2(s5_mul1_0_1_n63), .ZN(
        s5_mul1_0_1_n59) );
  INV_X1 s5_mul1_0_1_U13 ( .A(s5_mul1_0_1_n58), .ZN(s5_mul1_0_1_n65) );
  XNOR2_X1 s5_mul1_0_1_U12 ( .A(s5_mul1_0_1_n57), .B(s5_mul1_0_1_n56), .ZN(
        s5_concat[8]) );
  NAND2_X1 s5_mul1_0_1_U11 ( .A1(stage4Out[8]), .A2(s5_n5), .ZN(
        s5_mul1_0_1_n56) );
  XOR2_X1 s5_mul1_0_1_U10 ( .A(s5_mul1_0_1_n66), .B(s5_mul1_0_1_n70), .Z(
        s5_mul1_0_1_n57) );
  XNOR2_X1 s5_mul1_0_1_U9 ( .A(s5_mul1_0_1_n55), .B(s5_mul1_0_1_n54), .ZN(
        s5_mul1_0_1_n70) );
  NAND2_X1 s5_mul1_0_1_U8 ( .A1(s5_mul1_0_1_n61), .A2(s5_mul1_0_1_n58), .ZN(
        s5_mul1_0_1_n54) );
  XOR2_X1 s5_mul1_0_1_U7 ( .A(s5_n6), .B(s5_n8), .Z(s5_mul1_0_1_n58) );
  XOR2_X1 s5_mul1_0_1_U6 ( .A(stage4Out[9]), .B(stage4Out[11]), .Z(
        s5_mul1_0_1_n61) );
  NOR2_X1 s5_mul1_0_1_U5 ( .A1(s5_mul1_0_1_n63), .A2(s5_mul1_0_1_n60), .ZN(
        s5_mul1_0_1_n55) );
  XNOR2_X1 s5_mul1_0_1_U4 ( .A(stage4Out[8]), .B(stage4Out[10]), .ZN(
        s5_mul1_0_1_n60) );
  XNOR2_X1 s5_mul1_0_1_U3 ( .A(s5_n5), .B(s5_n7), .ZN(s5_mul1_0_1_n63) );
  AOI221_X1 s5_mul1_0_1_U2 ( .B1(s5_n5), .B2(s5_n6), .C1(stage4Out[8]), .C2(
        stage4Out[9]), .A(s5_mul1_0_1_n53), .ZN(s5_mul1_0_1_n66) );
  OAI22_X1 s5_mul1_0_1_U1 ( .A1(s5_n5), .A2(s5_n6), .B1(stage4Out[9]), .B2(
        stage4Out[8]), .ZN(s5_mul1_0_1_n53) );
  XNOR2_X1 s5_mul1_0_0_U28 ( .A(s5_mul1_0_0_n76), .B(s5_mul1_0_0_n75), .ZN(
        s5_concat[3]) );
  NAND2_X1 s5_mul1_0_0_U27 ( .A1(s5_n4), .A2(stage4Out[11]), .ZN(
        s5_mul1_0_0_n75) );
  XOR2_X1 s5_mul1_0_0_U26 ( .A(s5_mul1_0_0_n74), .B(s5_mul1_0_0_n73), .Z(
        s5_mul1_0_0_n76) );
  XNOR2_X1 s5_mul1_0_0_U25 ( .A(s5_mul1_0_0_n72), .B(s5_mul1_0_0_n71), .ZN(
        s5_concat[2]) );
  NAND2_X1 s5_mul1_0_0_U24 ( .A1(stage4Out[10]), .A2(s5_n3), .ZN(
        s5_mul1_0_0_n71) );
  XOR2_X1 s5_mul1_0_0_U23 ( .A(s5_mul1_0_0_n73), .B(s5_mul1_0_0_n70), .Z(
        s5_mul1_0_0_n72) );
  AOI221_X1 s5_mul1_0_0_U22 ( .B1(s5_n3), .B2(s5_n4), .C1(stage4Out[10]), .C2(
        stage4Out[11]), .A(s5_mul1_0_0_n69), .ZN(s5_mul1_0_0_n73) );
  OAI22_X1 s5_mul1_0_0_U21 ( .A1(s5_n3), .A2(s5_n4), .B1(stage4Out[11]), .B2(
        stage4Out[10]), .ZN(s5_mul1_0_0_n69) );
  XNOR2_X1 s5_mul1_0_0_U20 ( .A(s5_mul1_0_0_n68), .B(s5_mul1_0_0_n67), .ZN(
        s5_concat[1]) );
  NAND2_X1 s5_mul1_0_0_U19 ( .A1(s5_n2), .A2(stage4Out[9]), .ZN(
        s5_mul1_0_0_n67) );
  XOR2_X1 s5_mul1_0_0_U18 ( .A(s5_mul1_0_0_n74), .B(s5_mul1_0_0_n66), .Z(
        s5_mul1_0_0_n68) );
  OAI22_X1 s5_mul1_0_0_U17 ( .A1(s5_mul1_0_0_n65), .A2(s5_mul1_0_0_n64), .B1(
        s5_mul1_0_0_n63), .B2(s5_mul1_0_0_n62), .ZN(s5_mul1_0_0_n74) );
  NAND2_X1 s5_mul1_0_0_U16 ( .A1(s5_mul1_0_0_n61), .A2(s5_mul1_0_0_n65), .ZN(
        s5_mul1_0_0_n62) );
  XNOR2_X1 s5_mul1_0_0_U15 ( .A(s5_mul1_0_0_n60), .B(s5_mul1_0_0_n59), .ZN(
        s5_mul1_0_0_n64) );
  NAND2_X1 s5_mul1_0_0_U14 ( .A1(s5_mul1_0_0_n61), .A2(s5_mul1_0_0_n63), .ZN(
        s5_mul1_0_0_n59) );
  INV_X1 s5_mul1_0_0_U13 ( .A(s5_mul1_0_0_n58), .ZN(s5_mul1_0_0_n65) );
  XNOR2_X1 s5_mul1_0_0_U12 ( .A(s5_mul1_0_0_n57), .B(s5_mul1_0_0_n56), .ZN(
        s5_concat[0]) );
  NAND2_X1 s5_mul1_0_0_U11 ( .A1(stage4Out[8]), .A2(s5_n1), .ZN(
        s5_mul1_0_0_n56) );
  XOR2_X1 s5_mul1_0_0_U10 ( .A(s5_mul1_0_0_n66), .B(s5_mul1_0_0_n70), .Z(
        s5_mul1_0_0_n57) );
  XNOR2_X1 s5_mul1_0_0_U9 ( .A(s5_mul1_0_0_n55), .B(s5_mul1_0_0_n54), .ZN(
        s5_mul1_0_0_n70) );
  NAND2_X1 s5_mul1_0_0_U8 ( .A1(s5_mul1_0_0_n61), .A2(s5_mul1_0_0_n58), .ZN(
        s5_mul1_0_0_n54) );
  XOR2_X1 s5_mul1_0_0_U7 ( .A(s5_n2), .B(s5_n4), .Z(s5_mul1_0_0_n58) );
  XOR2_X1 s5_mul1_0_0_U6 ( .A(stage4Out[9]), .B(stage4Out[11]), .Z(
        s5_mul1_0_0_n61) );
  NOR2_X1 s5_mul1_0_0_U5 ( .A1(s5_mul1_0_0_n63), .A2(s5_mul1_0_0_n60), .ZN(
        s5_mul1_0_0_n55) );
  XNOR2_X1 s5_mul1_0_0_U4 ( .A(stage4Out[8]), .B(stage4Out[10]), .ZN(
        s5_mul1_0_0_n60) );
  XNOR2_X1 s5_mul1_0_0_U3 ( .A(s5_n1), .B(s5_n3), .ZN(s5_mul1_0_0_n63) );
  AOI221_X1 s5_mul1_0_0_U2 ( .B1(s5_n1), .B2(s5_n2), .C1(stage4Out[8]), .C2(
        stage4Out[9]), .A(s5_mul1_0_0_n53), .ZN(s5_mul1_0_0_n66) );
  OAI22_X1 s5_mul1_0_0_U1 ( .A1(s5_n1), .A2(s5_n2), .B1(stage4Out[9]), .B2(
        stage4Out[8]), .ZN(s5_mul1_0_0_n53) );
  XNOR2_X1 s5_mul2_2_2_U28 ( .A(s5_mul2_2_2_n76), .B(s5_mul2_2_2_n75), .ZN(
        s5_concat[71]) );
  NAND2_X1 s5_mul2_2_2_U27 ( .A1(stage4Out[27]), .A2(s5_n12), .ZN(
        s5_mul2_2_2_n75) );
  XOR2_X1 s5_mul2_2_2_U26 ( .A(s5_mul2_2_2_n74), .B(s5_mul2_2_2_n73), .Z(
        s5_mul2_2_2_n76) );
  XNOR2_X1 s5_mul2_2_2_U25 ( .A(s5_mul2_2_2_n72), .B(s5_mul2_2_2_n71), .ZN(
        s5_concat[70]) );
  NAND2_X1 s5_mul2_2_2_U24 ( .A1(s5_n11), .A2(stage4Out[26]), .ZN(
        s5_mul2_2_2_n71) );
  XOR2_X1 s5_mul2_2_2_U23 ( .A(s5_mul2_2_2_n73), .B(s5_mul2_2_2_n70), .Z(
        s5_mul2_2_2_n72) );
  AOI221_X1 s5_mul2_2_2_U22 ( .B1(stage4Out[26]), .B2(stage4Out[27]), .C1(
        s5_n11), .C2(s5_n12), .A(s5_mul2_2_2_n69), .ZN(s5_mul2_2_2_n73) );
  OAI22_X1 s5_mul2_2_2_U21 ( .A1(stage4Out[26]), .A2(stage4Out[27]), .B1(
        s5_n12), .B2(s5_n11), .ZN(s5_mul2_2_2_n69) );
  XNOR2_X1 s5_mul2_2_2_U20 ( .A(s5_mul2_2_2_n68), .B(s5_mul2_2_2_n67), .ZN(
        s5_concat[69]) );
  NAND2_X1 s5_mul2_2_2_U19 ( .A1(stage4Out[25]), .A2(s5_n10), .ZN(
        s5_mul2_2_2_n67) );
  XOR2_X1 s5_mul2_2_2_U18 ( .A(s5_mul2_2_2_n74), .B(s5_mul2_2_2_n66), .Z(
        s5_mul2_2_2_n68) );
  OAI22_X1 s5_mul2_2_2_U17 ( .A1(s5_mul2_2_2_n65), .A2(s5_mul2_2_2_n64), .B1(
        s5_mul2_2_2_n63), .B2(s5_mul2_2_2_n62), .ZN(s5_mul2_2_2_n74) );
  NAND2_X1 s5_mul2_2_2_U16 ( .A1(s5_mul2_2_2_n61), .A2(s5_mul2_2_2_n65), .ZN(
        s5_mul2_2_2_n62) );
  XNOR2_X1 s5_mul2_2_2_U15 ( .A(s5_mul2_2_2_n60), .B(s5_mul2_2_2_n59), .ZN(
        s5_mul2_2_2_n64) );
  NAND2_X1 s5_mul2_2_2_U14 ( .A1(s5_mul2_2_2_n61), .A2(s5_mul2_2_2_n63), .ZN(
        s5_mul2_2_2_n59) );
  INV_X1 s5_mul2_2_2_U13 ( .A(s5_mul2_2_2_n58), .ZN(s5_mul2_2_2_n65) );
  XNOR2_X1 s5_mul2_2_2_U12 ( .A(s5_mul2_2_2_n57), .B(s5_mul2_2_2_n56), .ZN(
        s5_concat[68]) );
  NAND2_X1 s5_mul2_2_2_U11 ( .A1(s5_n9), .A2(stage4Out[24]), .ZN(
        s5_mul2_2_2_n56) );
  XOR2_X1 s5_mul2_2_2_U10 ( .A(s5_mul2_2_2_n66), .B(s5_mul2_2_2_n70), .Z(
        s5_mul2_2_2_n57) );
  XNOR2_X1 s5_mul2_2_2_U9 ( .A(s5_mul2_2_2_n55), .B(s5_mul2_2_2_n54), .ZN(
        s5_mul2_2_2_n70) );
  NAND2_X1 s5_mul2_2_2_U8 ( .A1(s5_mul2_2_2_n61), .A2(s5_mul2_2_2_n58), .ZN(
        s5_mul2_2_2_n54) );
  XOR2_X1 s5_mul2_2_2_U7 ( .A(stage4Out[25]), .B(stage4Out[27]), .Z(
        s5_mul2_2_2_n58) );
  XOR2_X1 s5_mul2_2_2_U6 ( .A(s5_n10), .B(s5_n12), .Z(s5_mul2_2_2_n61) );
  NOR2_X1 s5_mul2_2_2_U5 ( .A1(s5_mul2_2_2_n63), .A2(s5_mul2_2_2_n60), .ZN(
        s5_mul2_2_2_n55) );
  XNOR2_X1 s5_mul2_2_2_U4 ( .A(s5_n9), .B(s5_n11), .ZN(s5_mul2_2_2_n60) );
  XNOR2_X1 s5_mul2_2_2_U3 ( .A(stage4Out[24]), .B(stage4Out[26]), .ZN(
        s5_mul2_2_2_n63) );
  AOI221_X1 s5_mul2_2_2_U2 ( .B1(stage4Out[24]), .B2(stage4Out[25]), .C1(s5_n9), .C2(s5_n10), .A(s5_mul2_2_2_n53), .ZN(s5_mul2_2_2_n66) );
  OAI22_X1 s5_mul2_2_2_U1 ( .A1(stage4Out[24]), .A2(stage4Out[25]), .B1(s5_n10), .B2(s5_n9), .ZN(s5_mul2_2_2_n53) );
  XNOR2_X1 s5_mul2_2_1_U28 ( .A(s5_mul2_2_1_n76), .B(s5_mul2_2_1_n75), .ZN(
        s5_concat[63]) );
  NAND2_X1 s5_mul2_2_1_U27 ( .A1(stage4Out[15]), .A2(s5_n12), .ZN(
        s5_mul2_2_1_n75) );
  XOR2_X1 s5_mul2_2_1_U26 ( .A(s5_mul2_2_1_n74), .B(s5_mul2_2_1_n73), .Z(
        s5_mul2_2_1_n76) );
  XNOR2_X1 s5_mul2_2_1_U25 ( .A(s5_mul2_2_1_n72), .B(s5_mul2_2_1_n71), .ZN(
        s5_concat[62]) );
  NAND2_X1 s5_mul2_2_1_U24 ( .A1(s5_n11), .A2(stage4Out[14]), .ZN(
        s5_mul2_2_1_n71) );
  XOR2_X1 s5_mul2_2_1_U23 ( .A(s5_mul2_2_1_n73), .B(s5_mul2_2_1_n70), .Z(
        s5_mul2_2_1_n72) );
  AOI221_X1 s5_mul2_2_1_U22 ( .B1(stage4Out[14]), .B2(stage4Out[15]), .C1(
        s5_n11), .C2(s5_n12), .A(s5_mul2_2_1_n69), .ZN(s5_mul2_2_1_n73) );
  OAI22_X1 s5_mul2_2_1_U21 ( .A1(stage4Out[14]), .A2(stage4Out[15]), .B1(
        s5_n12), .B2(s5_n11), .ZN(s5_mul2_2_1_n69) );
  XNOR2_X1 s5_mul2_2_1_U20 ( .A(s5_mul2_2_1_n68), .B(s5_mul2_2_1_n67), .ZN(
        s5_concat[61]) );
  NAND2_X1 s5_mul2_2_1_U19 ( .A1(stage4Out[13]), .A2(s5_n10), .ZN(
        s5_mul2_2_1_n67) );
  XOR2_X1 s5_mul2_2_1_U18 ( .A(s5_mul2_2_1_n74), .B(s5_mul2_2_1_n66), .Z(
        s5_mul2_2_1_n68) );
  OAI22_X1 s5_mul2_2_1_U17 ( .A1(s5_mul2_2_1_n65), .A2(s5_mul2_2_1_n64), .B1(
        s5_mul2_2_1_n63), .B2(s5_mul2_2_1_n62), .ZN(s5_mul2_2_1_n74) );
  NAND2_X1 s5_mul2_2_1_U16 ( .A1(s5_mul2_2_1_n61), .A2(s5_mul2_2_1_n65), .ZN(
        s5_mul2_2_1_n62) );
  XNOR2_X1 s5_mul2_2_1_U15 ( .A(s5_mul2_2_1_n60), .B(s5_mul2_2_1_n59), .ZN(
        s5_mul2_2_1_n64) );
  NAND2_X1 s5_mul2_2_1_U14 ( .A1(s5_mul2_2_1_n61), .A2(s5_mul2_2_1_n63), .ZN(
        s5_mul2_2_1_n59) );
  INV_X1 s5_mul2_2_1_U13 ( .A(s5_mul2_2_1_n58), .ZN(s5_mul2_2_1_n65) );
  XNOR2_X1 s5_mul2_2_1_U12 ( .A(s5_mul2_2_1_n57), .B(s5_mul2_2_1_n56), .ZN(
        s5_concat[60]) );
  NAND2_X1 s5_mul2_2_1_U11 ( .A1(s5_n9), .A2(stage4Out[12]), .ZN(
        s5_mul2_2_1_n56) );
  XOR2_X1 s5_mul2_2_1_U10 ( .A(s5_mul2_2_1_n66), .B(s5_mul2_2_1_n70), .Z(
        s5_mul2_2_1_n57) );
  XNOR2_X1 s5_mul2_2_1_U9 ( .A(s5_mul2_2_1_n55), .B(s5_mul2_2_1_n54), .ZN(
        s5_mul2_2_1_n70) );
  NAND2_X1 s5_mul2_2_1_U8 ( .A1(s5_mul2_2_1_n61), .A2(s5_mul2_2_1_n58), .ZN(
        s5_mul2_2_1_n54) );
  XOR2_X1 s5_mul2_2_1_U7 ( .A(stage4Out[13]), .B(stage4Out[15]), .Z(
        s5_mul2_2_1_n58) );
  XOR2_X1 s5_mul2_2_1_U6 ( .A(s5_n10), .B(s5_n12), .Z(s5_mul2_2_1_n61) );
  NOR2_X1 s5_mul2_2_1_U5 ( .A1(s5_mul2_2_1_n63), .A2(s5_mul2_2_1_n60), .ZN(
        s5_mul2_2_1_n55) );
  XNOR2_X1 s5_mul2_2_1_U4 ( .A(s5_n9), .B(s5_n11), .ZN(s5_mul2_2_1_n60) );
  XNOR2_X1 s5_mul2_2_1_U3 ( .A(stage4Out[12]), .B(stage4Out[14]), .ZN(
        s5_mul2_2_1_n63) );
  AOI221_X1 s5_mul2_2_1_U2 ( .B1(stage4Out[12]), .B2(stage4Out[13]), .C1(s5_n9), .C2(s5_n10), .A(s5_mul2_2_1_n53), .ZN(s5_mul2_2_1_n66) );
  OAI22_X1 s5_mul2_2_1_U1 ( .A1(stage4Out[12]), .A2(stage4Out[13]), .B1(s5_n10), .B2(s5_n9), .ZN(s5_mul2_2_1_n53) );
  XNOR2_X1 s5_mul2_2_0_U28 ( .A(s5_mul2_2_0_n76), .B(s5_mul2_2_0_n75), .ZN(
        s5_concat[55]) );
  NAND2_X1 s5_mul2_2_0_U27 ( .A1(stage4Out[3]), .A2(s5_n12), .ZN(
        s5_mul2_2_0_n75) );
  XOR2_X1 s5_mul2_2_0_U26 ( .A(s5_mul2_2_0_n74), .B(s5_mul2_2_0_n73), .Z(
        s5_mul2_2_0_n76) );
  XNOR2_X1 s5_mul2_2_0_U25 ( .A(s5_mul2_2_0_n72), .B(s5_mul2_2_0_n71), .ZN(
        s5_concat[54]) );
  NAND2_X1 s5_mul2_2_0_U24 ( .A1(s5_n11), .A2(stage4Out[2]), .ZN(
        s5_mul2_2_0_n71) );
  XOR2_X1 s5_mul2_2_0_U23 ( .A(s5_mul2_2_0_n73), .B(s5_mul2_2_0_n70), .Z(
        s5_mul2_2_0_n72) );
  AOI221_X1 s5_mul2_2_0_U22 ( .B1(stage4Out[2]), .B2(stage4Out[3]), .C1(s5_n11), .C2(s5_n12), .A(s5_mul2_2_0_n69), .ZN(s5_mul2_2_0_n73) );
  OAI22_X1 s5_mul2_2_0_U21 ( .A1(stage4Out[2]), .A2(stage4Out[3]), .B1(s5_n12), 
        .B2(s5_n11), .ZN(s5_mul2_2_0_n69) );
  XNOR2_X1 s5_mul2_2_0_U20 ( .A(s5_mul2_2_0_n68), .B(s5_mul2_2_0_n67), .ZN(
        s5_concat[53]) );
  NAND2_X1 s5_mul2_2_0_U19 ( .A1(stage4Out[1]), .A2(s5_n10), .ZN(
        s5_mul2_2_0_n67) );
  XOR2_X1 s5_mul2_2_0_U18 ( .A(s5_mul2_2_0_n74), .B(s5_mul2_2_0_n66), .Z(
        s5_mul2_2_0_n68) );
  OAI22_X1 s5_mul2_2_0_U17 ( .A1(s5_mul2_2_0_n65), .A2(s5_mul2_2_0_n64), .B1(
        s5_mul2_2_0_n63), .B2(s5_mul2_2_0_n62), .ZN(s5_mul2_2_0_n74) );
  NAND2_X1 s5_mul2_2_0_U16 ( .A1(s5_mul2_2_0_n61), .A2(s5_mul2_2_0_n65), .ZN(
        s5_mul2_2_0_n62) );
  XNOR2_X1 s5_mul2_2_0_U15 ( .A(s5_mul2_2_0_n60), .B(s5_mul2_2_0_n59), .ZN(
        s5_mul2_2_0_n64) );
  NAND2_X1 s5_mul2_2_0_U14 ( .A1(s5_mul2_2_0_n61), .A2(s5_mul2_2_0_n63), .ZN(
        s5_mul2_2_0_n59) );
  INV_X1 s5_mul2_2_0_U13 ( .A(s5_mul2_2_0_n58), .ZN(s5_mul2_2_0_n65) );
  XNOR2_X1 s5_mul2_2_0_U12 ( .A(s5_mul2_2_0_n57), .B(s5_mul2_2_0_n56), .ZN(
        s5_concat[52]) );
  NAND2_X1 s5_mul2_2_0_U11 ( .A1(s5_n9), .A2(stage4Out[0]), .ZN(
        s5_mul2_2_0_n56) );
  XOR2_X1 s5_mul2_2_0_U10 ( .A(s5_mul2_2_0_n66), .B(s5_mul2_2_0_n70), .Z(
        s5_mul2_2_0_n57) );
  XNOR2_X1 s5_mul2_2_0_U9 ( .A(s5_mul2_2_0_n55), .B(s5_mul2_2_0_n54), .ZN(
        s5_mul2_2_0_n70) );
  NAND2_X1 s5_mul2_2_0_U8 ( .A1(s5_mul2_2_0_n61), .A2(s5_mul2_2_0_n58), .ZN(
        s5_mul2_2_0_n54) );
  XOR2_X1 s5_mul2_2_0_U7 ( .A(stage4Out[1]), .B(stage4Out[3]), .Z(
        s5_mul2_2_0_n58) );
  XOR2_X1 s5_mul2_2_0_U6 ( .A(s5_n10), .B(s5_n12), .Z(s5_mul2_2_0_n61) );
  NOR2_X1 s5_mul2_2_0_U5 ( .A1(s5_mul2_2_0_n63), .A2(s5_mul2_2_0_n60), .ZN(
        s5_mul2_2_0_n55) );
  XNOR2_X1 s5_mul2_2_0_U4 ( .A(s5_n9), .B(s5_n11), .ZN(s5_mul2_2_0_n60) );
  XNOR2_X1 s5_mul2_2_0_U3 ( .A(stage4Out[0]), .B(stage4Out[2]), .ZN(
        s5_mul2_2_0_n63) );
  AOI221_X1 s5_mul2_2_0_U2 ( .B1(stage4Out[0]), .B2(stage4Out[1]), .C1(s5_n9), 
        .C2(s5_n10), .A(s5_mul2_2_0_n53), .ZN(s5_mul2_2_0_n66) );
  OAI22_X1 s5_mul2_2_0_U1 ( .A1(stage4Out[0]), .A2(stage4Out[1]), .B1(s5_n10), 
        .B2(s5_n9), .ZN(s5_mul2_2_0_n53) );
  XNOR2_X1 s5_mul2_1_2_U28 ( .A(s5_mul2_1_2_n76), .B(s5_mul2_1_2_n75), .ZN(
        s5_concat[47]) );
  NAND2_X1 s5_mul2_1_2_U27 ( .A1(stage4Out[27]), .A2(s5_n8), .ZN(
        s5_mul2_1_2_n75) );
  XOR2_X1 s5_mul2_1_2_U26 ( .A(s5_mul2_1_2_n74), .B(s5_mul2_1_2_n73), .Z(
        s5_mul2_1_2_n76) );
  XNOR2_X1 s5_mul2_1_2_U25 ( .A(s5_mul2_1_2_n72), .B(s5_mul2_1_2_n71), .ZN(
        s5_concat[46]) );
  NAND2_X1 s5_mul2_1_2_U24 ( .A1(s5_n7), .A2(stage4Out[26]), .ZN(
        s5_mul2_1_2_n71) );
  XOR2_X1 s5_mul2_1_2_U23 ( .A(s5_mul2_1_2_n73), .B(s5_mul2_1_2_n70), .Z(
        s5_mul2_1_2_n72) );
  AOI221_X1 s5_mul2_1_2_U22 ( .B1(stage4Out[26]), .B2(stage4Out[27]), .C1(
        s5_n7), .C2(s5_n8), .A(s5_mul2_1_2_n69), .ZN(s5_mul2_1_2_n73) );
  OAI22_X1 s5_mul2_1_2_U21 ( .A1(stage4Out[26]), .A2(stage4Out[27]), .B1(s5_n8), .B2(s5_n7), .ZN(s5_mul2_1_2_n69) );
  XNOR2_X1 s5_mul2_1_2_U20 ( .A(s5_mul2_1_2_n68), .B(s5_mul2_1_2_n67), .ZN(
        s5_concat[45]) );
  NAND2_X1 s5_mul2_1_2_U19 ( .A1(stage4Out[25]), .A2(s5_n6), .ZN(
        s5_mul2_1_2_n67) );
  XOR2_X1 s5_mul2_1_2_U18 ( .A(s5_mul2_1_2_n74), .B(s5_mul2_1_2_n66), .Z(
        s5_mul2_1_2_n68) );
  OAI22_X1 s5_mul2_1_2_U17 ( .A1(s5_mul2_1_2_n65), .A2(s5_mul2_1_2_n64), .B1(
        s5_mul2_1_2_n63), .B2(s5_mul2_1_2_n62), .ZN(s5_mul2_1_2_n74) );
  NAND2_X1 s5_mul2_1_2_U16 ( .A1(s5_mul2_1_2_n61), .A2(s5_mul2_1_2_n65), .ZN(
        s5_mul2_1_2_n62) );
  XNOR2_X1 s5_mul2_1_2_U15 ( .A(s5_mul2_1_2_n60), .B(s5_mul2_1_2_n59), .ZN(
        s5_mul2_1_2_n64) );
  NAND2_X1 s5_mul2_1_2_U14 ( .A1(s5_mul2_1_2_n61), .A2(s5_mul2_1_2_n63), .ZN(
        s5_mul2_1_2_n59) );
  INV_X1 s5_mul2_1_2_U13 ( .A(s5_mul2_1_2_n58), .ZN(s5_mul2_1_2_n65) );
  XNOR2_X1 s5_mul2_1_2_U12 ( .A(s5_mul2_1_2_n57), .B(s5_mul2_1_2_n56), .ZN(
        s5_concat[44]) );
  NAND2_X1 s5_mul2_1_2_U11 ( .A1(s5_n5), .A2(stage4Out[24]), .ZN(
        s5_mul2_1_2_n56) );
  XOR2_X1 s5_mul2_1_2_U10 ( .A(s5_mul2_1_2_n66), .B(s5_mul2_1_2_n70), .Z(
        s5_mul2_1_2_n57) );
  XNOR2_X1 s5_mul2_1_2_U9 ( .A(s5_mul2_1_2_n55), .B(s5_mul2_1_2_n54), .ZN(
        s5_mul2_1_2_n70) );
  NAND2_X1 s5_mul2_1_2_U8 ( .A1(s5_mul2_1_2_n61), .A2(s5_mul2_1_2_n58), .ZN(
        s5_mul2_1_2_n54) );
  XOR2_X1 s5_mul2_1_2_U7 ( .A(stage4Out[25]), .B(stage4Out[27]), .Z(
        s5_mul2_1_2_n58) );
  XOR2_X1 s5_mul2_1_2_U6 ( .A(s5_n6), .B(s5_n8), .Z(s5_mul2_1_2_n61) );
  NOR2_X1 s5_mul2_1_2_U5 ( .A1(s5_mul2_1_2_n63), .A2(s5_mul2_1_2_n60), .ZN(
        s5_mul2_1_2_n55) );
  XNOR2_X1 s5_mul2_1_2_U4 ( .A(s5_n5), .B(s5_n7), .ZN(s5_mul2_1_2_n60) );
  XNOR2_X1 s5_mul2_1_2_U3 ( .A(stage4Out[24]), .B(stage4Out[26]), .ZN(
        s5_mul2_1_2_n63) );
  AOI221_X1 s5_mul2_1_2_U2 ( .B1(stage4Out[24]), .B2(stage4Out[25]), .C1(s5_n5), .C2(s5_n6), .A(s5_mul2_1_2_n53), .ZN(s5_mul2_1_2_n66) );
  OAI22_X1 s5_mul2_1_2_U1 ( .A1(stage4Out[24]), .A2(stage4Out[25]), .B1(s5_n6), 
        .B2(s5_n5), .ZN(s5_mul2_1_2_n53) );
  XNOR2_X1 s5_mul2_1_1_U28 ( .A(s5_mul2_1_1_n76), .B(s5_mul2_1_1_n75), .ZN(
        s5_concat[39]) );
  NAND2_X1 s5_mul2_1_1_U27 ( .A1(stage4Out[15]), .A2(s5_n8), .ZN(
        s5_mul2_1_1_n75) );
  XOR2_X1 s5_mul2_1_1_U26 ( .A(s5_mul2_1_1_n74), .B(s5_mul2_1_1_n73), .Z(
        s5_mul2_1_1_n76) );
  XNOR2_X1 s5_mul2_1_1_U25 ( .A(s5_mul2_1_1_n72), .B(s5_mul2_1_1_n71), .ZN(
        s5_concat[38]) );
  NAND2_X1 s5_mul2_1_1_U24 ( .A1(s5_n7), .A2(stage4Out[14]), .ZN(
        s5_mul2_1_1_n71) );
  XOR2_X1 s5_mul2_1_1_U23 ( .A(s5_mul2_1_1_n73), .B(s5_mul2_1_1_n70), .Z(
        s5_mul2_1_1_n72) );
  AOI221_X1 s5_mul2_1_1_U22 ( .B1(stage4Out[14]), .B2(stage4Out[15]), .C1(
        s5_n7), .C2(s5_n8), .A(s5_mul2_1_1_n69), .ZN(s5_mul2_1_1_n73) );
  OAI22_X1 s5_mul2_1_1_U21 ( .A1(stage4Out[14]), .A2(stage4Out[15]), .B1(s5_n8), .B2(s5_n7), .ZN(s5_mul2_1_1_n69) );
  XNOR2_X1 s5_mul2_1_1_U20 ( .A(s5_mul2_1_1_n68), .B(s5_mul2_1_1_n67), .ZN(
        s5_concat[37]) );
  NAND2_X1 s5_mul2_1_1_U19 ( .A1(stage4Out[13]), .A2(s5_n6), .ZN(
        s5_mul2_1_1_n67) );
  XOR2_X1 s5_mul2_1_1_U18 ( .A(s5_mul2_1_1_n74), .B(s5_mul2_1_1_n66), .Z(
        s5_mul2_1_1_n68) );
  OAI22_X1 s5_mul2_1_1_U17 ( .A1(s5_mul2_1_1_n65), .A2(s5_mul2_1_1_n64), .B1(
        s5_mul2_1_1_n63), .B2(s5_mul2_1_1_n62), .ZN(s5_mul2_1_1_n74) );
  NAND2_X1 s5_mul2_1_1_U16 ( .A1(s5_mul2_1_1_n61), .A2(s5_mul2_1_1_n65), .ZN(
        s5_mul2_1_1_n62) );
  XNOR2_X1 s5_mul2_1_1_U15 ( .A(s5_mul2_1_1_n60), .B(s5_mul2_1_1_n59), .ZN(
        s5_mul2_1_1_n64) );
  NAND2_X1 s5_mul2_1_1_U14 ( .A1(s5_mul2_1_1_n61), .A2(s5_mul2_1_1_n63), .ZN(
        s5_mul2_1_1_n59) );
  INV_X1 s5_mul2_1_1_U13 ( .A(s5_mul2_1_1_n58), .ZN(s5_mul2_1_1_n65) );
  XNOR2_X1 s5_mul2_1_1_U12 ( .A(s5_mul2_1_1_n57), .B(s5_mul2_1_1_n56), .ZN(
        s5_concat[36]) );
  NAND2_X1 s5_mul2_1_1_U11 ( .A1(s5_n5), .A2(stage4Out[12]), .ZN(
        s5_mul2_1_1_n56) );
  XOR2_X1 s5_mul2_1_1_U10 ( .A(s5_mul2_1_1_n66), .B(s5_mul2_1_1_n70), .Z(
        s5_mul2_1_1_n57) );
  XNOR2_X1 s5_mul2_1_1_U9 ( .A(s5_mul2_1_1_n55), .B(s5_mul2_1_1_n54), .ZN(
        s5_mul2_1_1_n70) );
  NAND2_X1 s5_mul2_1_1_U8 ( .A1(s5_mul2_1_1_n61), .A2(s5_mul2_1_1_n58), .ZN(
        s5_mul2_1_1_n54) );
  XOR2_X1 s5_mul2_1_1_U7 ( .A(stage4Out[13]), .B(stage4Out[15]), .Z(
        s5_mul2_1_1_n58) );
  XOR2_X1 s5_mul2_1_1_U6 ( .A(s5_n6), .B(s5_n8), .Z(s5_mul2_1_1_n61) );
  NOR2_X1 s5_mul2_1_1_U5 ( .A1(s5_mul2_1_1_n63), .A2(s5_mul2_1_1_n60), .ZN(
        s5_mul2_1_1_n55) );
  XNOR2_X1 s5_mul2_1_1_U4 ( .A(s5_n5), .B(s5_n7), .ZN(s5_mul2_1_1_n60) );
  XNOR2_X1 s5_mul2_1_1_U3 ( .A(stage4Out[12]), .B(stage4Out[14]), .ZN(
        s5_mul2_1_1_n63) );
  AOI221_X1 s5_mul2_1_1_U2 ( .B1(stage4Out[12]), .B2(stage4Out[13]), .C1(s5_n5), .C2(s5_n6), .A(s5_mul2_1_1_n53), .ZN(s5_mul2_1_1_n66) );
  OAI22_X1 s5_mul2_1_1_U1 ( .A1(stage4Out[12]), .A2(stage4Out[13]), .B1(s5_n6), 
        .B2(s5_n5), .ZN(s5_mul2_1_1_n53) );
  XNOR2_X1 s5_mul2_1_0_U28 ( .A(s5_mul2_1_0_n76), .B(s5_mul2_1_0_n75), .ZN(
        s5_concat[31]) );
  NAND2_X1 s5_mul2_1_0_U27 ( .A1(stage4Out[3]), .A2(s5_n8), .ZN(
        s5_mul2_1_0_n75) );
  XOR2_X1 s5_mul2_1_0_U26 ( .A(s5_mul2_1_0_n74), .B(s5_mul2_1_0_n73), .Z(
        s5_mul2_1_0_n76) );
  XNOR2_X1 s5_mul2_1_0_U25 ( .A(s5_mul2_1_0_n72), .B(s5_mul2_1_0_n71), .ZN(
        s5_concat[30]) );
  NAND2_X1 s5_mul2_1_0_U24 ( .A1(s5_n7), .A2(stage4Out[2]), .ZN(
        s5_mul2_1_0_n71) );
  XOR2_X1 s5_mul2_1_0_U23 ( .A(s5_mul2_1_0_n73), .B(s5_mul2_1_0_n70), .Z(
        s5_mul2_1_0_n72) );
  AOI221_X1 s5_mul2_1_0_U22 ( .B1(stage4Out[2]), .B2(stage4Out[3]), .C1(s5_n7), 
        .C2(s5_n8), .A(s5_mul2_1_0_n69), .ZN(s5_mul2_1_0_n73) );
  OAI22_X1 s5_mul2_1_0_U21 ( .A1(stage4Out[2]), .A2(stage4Out[3]), .B1(s5_n8), 
        .B2(s5_n7), .ZN(s5_mul2_1_0_n69) );
  XNOR2_X1 s5_mul2_1_0_U20 ( .A(s5_mul2_1_0_n68), .B(s5_mul2_1_0_n67), .ZN(
        s5_concat[29]) );
  NAND2_X1 s5_mul2_1_0_U19 ( .A1(stage4Out[1]), .A2(s5_n6), .ZN(
        s5_mul2_1_0_n67) );
  XOR2_X1 s5_mul2_1_0_U18 ( .A(s5_mul2_1_0_n74), .B(s5_mul2_1_0_n66), .Z(
        s5_mul2_1_0_n68) );
  OAI22_X1 s5_mul2_1_0_U17 ( .A1(s5_mul2_1_0_n65), .A2(s5_mul2_1_0_n64), .B1(
        s5_mul2_1_0_n63), .B2(s5_mul2_1_0_n62), .ZN(s5_mul2_1_0_n74) );
  NAND2_X1 s5_mul2_1_0_U16 ( .A1(s5_mul2_1_0_n61), .A2(s5_mul2_1_0_n65), .ZN(
        s5_mul2_1_0_n62) );
  XNOR2_X1 s5_mul2_1_0_U15 ( .A(s5_mul2_1_0_n60), .B(s5_mul2_1_0_n59), .ZN(
        s5_mul2_1_0_n64) );
  NAND2_X1 s5_mul2_1_0_U14 ( .A1(s5_mul2_1_0_n61), .A2(s5_mul2_1_0_n63), .ZN(
        s5_mul2_1_0_n59) );
  INV_X1 s5_mul2_1_0_U13 ( .A(s5_mul2_1_0_n58), .ZN(s5_mul2_1_0_n65) );
  XNOR2_X1 s5_mul2_1_0_U12 ( .A(s5_mul2_1_0_n57), .B(s5_mul2_1_0_n56), .ZN(
        s5_concat[28]) );
  NAND2_X1 s5_mul2_1_0_U11 ( .A1(s5_n5), .A2(stage4Out[0]), .ZN(
        s5_mul2_1_0_n56) );
  XOR2_X1 s5_mul2_1_0_U10 ( .A(s5_mul2_1_0_n66), .B(s5_mul2_1_0_n70), .Z(
        s5_mul2_1_0_n57) );
  XNOR2_X1 s5_mul2_1_0_U9 ( .A(s5_mul2_1_0_n55), .B(s5_mul2_1_0_n54), .ZN(
        s5_mul2_1_0_n70) );
  NAND2_X1 s5_mul2_1_0_U8 ( .A1(s5_mul2_1_0_n61), .A2(s5_mul2_1_0_n58), .ZN(
        s5_mul2_1_0_n54) );
  XOR2_X1 s5_mul2_1_0_U7 ( .A(stage4Out[1]), .B(stage4Out[3]), .Z(
        s5_mul2_1_0_n58) );
  XOR2_X1 s5_mul2_1_0_U6 ( .A(s5_n6), .B(s5_n8), .Z(s5_mul2_1_0_n61) );
  NOR2_X1 s5_mul2_1_0_U5 ( .A1(s5_mul2_1_0_n63), .A2(s5_mul2_1_0_n60), .ZN(
        s5_mul2_1_0_n55) );
  XNOR2_X1 s5_mul2_1_0_U4 ( .A(s5_n5), .B(s5_n7), .ZN(s5_mul2_1_0_n60) );
  XNOR2_X1 s5_mul2_1_0_U3 ( .A(stage4Out[0]), .B(stage4Out[2]), .ZN(
        s5_mul2_1_0_n63) );
  AOI221_X1 s5_mul2_1_0_U2 ( .B1(stage4Out[0]), .B2(stage4Out[1]), .C1(s5_n5), 
        .C2(s5_n6), .A(s5_mul2_1_0_n53), .ZN(s5_mul2_1_0_n66) );
  OAI22_X1 s5_mul2_1_0_U1 ( .A1(stage4Out[0]), .A2(stage4Out[1]), .B1(s5_n6), 
        .B2(s5_n5), .ZN(s5_mul2_1_0_n53) );
  XNOR2_X1 s5_mul2_0_2_U28 ( .A(s5_mul2_0_2_n76), .B(s5_mul2_0_2_n75), .ZN(
        s5_concat[23]) );
  NAND2_X1 s5_mul2_0_2_U27 ( .A1(stage4Out[27]), .A2(s5_n4), .ZN(
        s5_mul2_0_2_n75) );
  XOR2_X1 s5_mul2_0_2_U26 ( .A(s5_mul2_0_2_n74), .B(s5_mul2_0_2_n73), .Z(
        s5_mul2_0_2_n76) );
  XNOR2_X1 s5_mul2_0_2_U25 ( .A(s5_mul2_0_2_n72), .B(s5_mul2_0_2_n71), .ZN(
        s5_concat[22]) );
  NAND2_X1 s5_mul2_0_2_U24 ( .A1(s5_n3), .A2(stage4Out[26]), .ZN(
        s5_mul2_0_2_n71) );
  XOR2_X1 s5_mul2_0_2_U23 ( .A(s5_mul2_0_2_n73), .B(s5_mul2_0_2_n70), .Z(
        s5_mul2_0_2_n72) );
  AOI221_X1 s5_mul2_0_2_U22 ( .B1(stage4Out[26]), .B2(stage4Out[27]), .C1(
        s5_n3), .C2(s5_n4), .A(s5_mul2_0_2_n69), .ZN(s5_mul2_0_2_n73) );
  OAI22_X1 s5_mul2_0_2_U21 ( .A1(stage4Out[26]), .A2(stage4Out[27]), .B1(s5_n4), .B2(s5_n3), .ZN(s5_mul2_0_2_n69) );
  XNOR2_X1 s5_mul2_0_2_U20 ( .A(s5_mul2_0_2_n68), .B(s5_mul2_0_2_n67), .ZN(
        s5_concat[21]) );
  NAND2_X1 s5_mul2_0_2_U19 ( .A1(stage4Out[25]), .A2(s5_n2), .ZN(
        s5_mul2_0_2_n67) );
  XOR2_X1 s5_mul2_0_2_U18 ( .A(s5_mul2_0_2_n74), .B(s5_mul2_0_2_n66), .Z(
        s5_mul2_0_2_n68) );
  OAI22_X1 s5_mul2_0_2_U17 ( .A1(s5_mul2_0_2_n65), .A2(s5_mul2_0_2_n64), .B1(
        s5_mul2_0_2_n63), .B2(s5_mul2_0_2_n62), .ZN(s5_mul2_0_2_n74) );
  NAND2_X1 s5_mul2_0_2_U16 ( .A1(s5_mul2_0_2_n61), .A2(s5_mul2_0_2_n65), .ZN(
        s5_mul2_0_2_n62) );
  XNOR2_X1 s5_mul2_0_2_U15 ( .A(s5_mul2_0_2_n60), .B(s5_mul2_0_2_n59), .ZN(
        s5_mul2_0_2_n64) );
  NAND2_X1 s5_mul2_0_2_U14 ( .A1(s5_mul2_0_2_n61), .A2(s5_mul2_0_2_n63), .ZN(
        s5_mul2_0_2_n59) );
  INV_X1 s5_mul2_0_2_U13 ( .A(s5_mul2_0_2_n58), .ZN(s5_mul2_0_2_n65) );
  XNOR2_X1 s5_mul2_0_2_U12 ( .A(s5_mul2_0_2_n57), .B(s5_mul2_0_2_n56), .ZN(
        s5_concat[20]) );
  NAND2_X1 s5_mul2_0_2_U11 ( .A1(s5_n1), .A2(stage4Out[24]), .ZN(
        s5_mul2_0_2_n56) );
  XOR2_X1 s5_mul2_0_2_U10 ( .A(s5_mul2_0_2_n66), .B(s5_mul2_0_2_n70), .Z(
        s5_mul2_0_2_n57) );
  XNOR2_X1 s5_mul2_0_2_U9 ( .A(s5_mul2_0_2_n55), .B(s5_mul2_0_2_n54), .ZN(
        s5_mul2_0_2_n70) );
  NAND2_X1 s5_mul2_0_2_U8 ( .A1(s5_mul2_0_2_n61), .A2(s5_mul2_0_2_n58), .ZN(
        s5_mul2_0_2_n54) );
  XOR2_X1 s5_mul2_0_2_U7 ( .A(stage4Out[25]), .B(stage4Out[27]), .Z(
        s5_mul2_0_2_n58) );
  XOR2_X1 s5_mul2_0_2_U6 ( .A(s5_n2), .B(s5_n4), .Z(s5_mul2_0_2_n61) );
  NOR2_X1 s5_mul2_0_2_U5 ( .A1(s5_mul2_0_2_n63), .A2(s5_mul2_0_2_n60), .ZN(
        s5_mul2_0_2_n55) );
  XNOR2_X1 s5_mul2_0_2_U4 ( .A(s5_n1), .B(s5_n3), .ZN(s5_mul2_0_2_n60) );
  XNOR2_X1 s5_mul2_0_2_U3 ( .A(stage4Out[24]), .B(stage4Out[26]), .ZN(
        s5_mul2_0_2_n63) );
  AOI221_X1 s5_mul2_0_2_U2 ( .B1(stage4Out[24]), .B2(stage4Out[25]), .C1(s5_n1), .C2(s5_n2), .A(s5_mul2_0_2_n53), .ZN(s5_mul2_0_2_n66) );
  OAI22_X1 s5_mul2_0_2_U1 ( .A1(stage4Out[24]), .A2(stage4Out[25]), .B1(s5_n2), 
        .B2(s5_n1), .ZN(s5_mul2_0_2_n53) );
  XNOR2_X1 s5_mul2_0_1_U28 ( .A(s5_mul2_0_1_n76), .B(s5_mul2_0_1_n75), .ZN(
        s5_concat[15]) );
  NAND2_X1 s5_mul2_0_1_U27 ( .A1(stage4Out[15]), .A2(s5_n4), .ZN(
        s5_mul2_0_1_n75) );
  XOR2_X1 s5_mul2_0_1_U26 ( .A(s5_mul2_0_1_n74), .B(s5_mul2_0_1_n73), .Z(
        s5_mul2_0_1_n76) );
  XNOR2_X1 s5_mul2_0_1_U25 ( .A(s5_mul2_0_1_n72), .B(s5_mul2_0_1_n71), .ZN(
        s5_concat[14]) );
  NAND2_X1 s5_mul2_0_1_U24 ( .A1(s5_n3), .A2(stage4Out[14]), .ZN(
        s5_mul2_0_1_n71) );
  XOR2_X1 s5_mul2_0_1_U23 ( .A(s5_mul2_0_1_n73), .B(s5_mul2_0_1_n70), .Z(
        s5_mul2_0_1_n72) );
  AOI221_X1 s5_mul2_0_1_U22 ( .B1(stage4Out[14]), .B2(stage4Out[15]), .C1(
        s5_n3), .C2(s5_n4), .A(s5_mul2_0_1_n69), .ZN(s5_mul2_0_1_n73) );
  OAI22_X1 s5_mul2_0_1_U21 ( .A1(stage4Out[14]), .A2(stage4Out[15]), .B1(s5_n4), .B2(s5_n3), .ZN(s5_mul2_0_1_n69) );
  XNOR2_X1 s5_mul2_0_1_U20 ( .A(s5_mul2_0_1_n68), .B(s5_mul2_0_1_n67), .ZN(
        s5_concat[13]) );
  NAND2_X1 s5_mul2_0_1_U19 ( .A1(stage4Out[13]), .A2(s5_n2), .ZN(
        s5_mul2_0_1_n67) );
  XOR2_X1 s5_mul2_0_1_U18 ( .A(s5_mul2_0_1_n74), .B(s5_mul2_0_1_n66), .Z(
        s5_mul2_0_1_n68) );
  OAI22_X1 s5_mul2_0_1_U17 ( .A1(s5_mul2_0_1_n65), .A2(s5_mul2_0_1_n64), .B1(
        s5_mul2_0_1_n63), .B2(s5_mul2_0_1_n62), .ZN(s5_mul2_0_1_n74) );
  NAND2_X1 s5_mul2_0_1_U16 ( .A1(s5_mul2_0_1_n61), .A2(s5_mul2_0_1_n65), .ZN(
        s5_mul2_0_1_n62) );
  XNOR2_X1 s5_mul2_0_1_U15 ( .A(s5_mul2_0_1_n60), .B(s5_mul2_0_1_n59), .ZN(
        s5_mul2_0_1_n64) );
  NAND2_X1 s5_mul2_0_1_U14 ( .A1(s5_mul2_0_1_n61), .A2(s5_mul2_0_1_n63), .ZN(
        s5_mul2_0_1_n59) );
  INV_X1 s5_mul2_0_1_U13 ( .A(s5_mul2_0_1_n58), .ZN(s5_mul2_0_1_n65) );
  XNOR2_X1 s5_mul2_0_1_U12 ( .A(s5_mul2_0_1_n57), .B(s5_mul2_0_1_n56), .ZN(
        s5_concat[12]) );
  NAND2_X1 s5_mul2_0_1_U11 ( .A1(s5_n1), .A2(stage4Out[12]), .ZN(
        s5_mul2_0_1_n56) );
  XOR2_X1 s5_mul2_0_1_U10 ( .A(s5_mul2_0_1_n66), .B(s5_mul2_0_1_n70), .Z(
        s5_mul2_0_1_n57) );
  XNOR2_X1 s5_mul2_0_1_U9 ( .A(s5_mul2_0_1_n55), .B(s5_mul2_0_1_n54), .ZN(
        s5_mul2_0_1_n70) );
  NAND2_X1 s5_mul2_0_1_U8 ( .A1(s5_mul2_0_1_n61), .A2(s5_mul2_0_1_n58), .ZN(
        s5_mul2_0_1_n54) );
  XOR2_X1 s5_mul2_0_1_U7 ( .A(stage4Out[13]), .B(stage4Out[15]), .Z(
        s5_mul2_0_1_n58) );
  XOR2_X1 s5_mul2_0_1_U6 ( .A(s5_n2), .B(s5_n4), .Z(s5_mul2_0_1_n61) );
  NOR2_X1 s5_mul2_0_1_U5 ( .A1(s5_mul2_0_1_n63), .A2(s5_mul2_0_1_n60), .ZN(
        s5_mul2_0_1_n55) );
  XNOR2_X1 s5_mul2_0_1_U4 ( .A(s5_n1), .B(s5_n3), .ZN(s5_mul2_0_1_n60) );
  XNOR2_X1 s5_mul2_0_1_U3 ( .A(stage4Out[12]), .B(stage4Out[14]), .ZN(
        s5_mul2_0_1_n63) );
  AOI221_X1 s5_mul2_0_1_U2 ( .B1(stage4Out[12]), .B2(stage4Out[13]), .C1(s5_n1), .C2(s5_n2), .A(s5_mul2_0_1_n53), .ZN(s5_mul2_0_1_n66) );
  OAI22_X1 s5_mul2_0_1_U1 ( .A1(stage4Out[12]), .A2(stage4Out[13]), .B1(s5_n2), 
        .B2(s5_n1), .ZN(s5_mul2_0_1_n53) );
  XNOR2_X1 s5_mul2_0_0_U28 ( .A(s5_mul2_0_0_n76), .B(s5_mul2_0_0_n75), .ZN(
        s5_concat[7]) );
  NAND2_X1 s5_mul2_0_0_U27 ( .A1(stage4Out[3]), .A2(s5_n4), .ZN(
        s5_mul2_0_0_n75) );
  XOR2_X1 s5_mul2_0_0_U26 ( .A(s5_mul2_0_0_n74), .B(s5_mul2_0_0_n73), .Z(
        s5_mul2_0_0_n76) );
  XNOR2_X1 s5_mul2_0_0_U25 ( .A(s5_mul2_0_0_n72), .B(s5_mul2_0_0_n71), .ZN(
        s5_concat[6]) );
  NAND2_X1 s5_mul2_0_0_U24 ( .A1(s5_n3), .A2(stage4Out[2]), .ZN(
        s5_mul2_0_0_n71) );
  XOR2_X1 s5_mul2_0_0_U23 ( .A(s5_mul2_0_0_n73), .B(s5_mul2_0_0_n70), .Z(
        s5_mul2_0_0_n72) );
  AOI221_X1 s5_mul2_0_0_U22 ( .B1(stage4Out[2]), .B2(stage4Out[3]), .C1(s5_n3), 
        .C2(s5_n4), .A(s5_mul2_0_0_n69), .ZN(s5_mul2_0_0_n73) );
  OAI22_X1 s5_mul2_0_0_U21 ( .A1(stage4Out[2]), .A2(stage4Out[3]), .B1(s5_n4), 
        .B2(s5_n3), .ZN(s5_mul2_0_0_n69) );
  XNOR2_X1 s5_mul2_0_0_U20 ( .A(s5_mul2_0_0_n68), .B(s5_mul2_0_0_n67), .ZN(
        s5_concat[5]) );
  NAND2_X1 s5_mul2_0_0_U19 ( .A1(stage4Out[1]), .A2(s5_n2), .ZN(
        s5_mul2_0_0_n67) );
  XOR2_X1 s5_mul2_0_0_U18 ( .A(s5_mul2_0_0_n74), .B(s5_mul2_0_0_n66), .Z(
        s5_mul2_0_0_n68) );
  OAI22_X1 s5_mul2_0_0_U17 ( .A1(s5_mul2_0_0_n65), .A2(s5_mul2_0_0_n64), .B1(
        s5_mul2_0_0_n63), .B2(s5_mul2_0_0_n62), .ZN(s5_mul2_0_0_n74) );
  NAND2_X1 s5_mul2_0_0_U16 ( .A1(s5_mul2_0_0_n61), .A2(s5_mul2_0_0_n65), .ZN(
        s5_mul2_0_0_n62) );
  XNOR2_X1 s5_mul2_0_0_U15 ( .A(s5_mul2_0_0_n60), .B(s5_mul2_0_0_n59), .ZN(
        s5_mul2_0_0_n64) );
  NAND2_X1 s5_mul2_0_0_U14 ( .A1(s5_mul2_0_0_n61), .A2(s5_mul2_0_0_n63), .ZN(
        s5_mul2_0_0_n59) );
  INV_X1 s5_mul2_0_0_U13 ( .A(s5_mul2_0_0_n58), .ZN(s5_mul2_0_0_n65) );
  XNOR2_X1 s5_mul2_0_0_U12 ( .A(s5_mul2_0_0_n57), .B(s5_mul2_0_0_n56), .ZN(
        s5_concat[4]) );
  NAND2_X1 s5_mul2_0_0_U11 ( .A1(s5_n1), .A2(stage4Out[0]), .ZN(
        s5_mul2_0_0_n56) );
  XOR2_X1 s5_mul2_0_0_U10 ( .A(s5_mul2_0_0_n66), .B(s5_mul2_0_0_n70), .Z(
        s5_mul2_0_0_n57) );
  XNOR2_X1 s5_mul2_0_0_U9 ( .A(s5_mul2_0_0_n55), .B(s5_mul2_0_0_n54), .ZN(
        s5_mul2_0_0_n70) );
  NAND2_X1 s5_mul2_0_0_U8 ( .A1(s5_mul2_0_0_n61), .A2(s5_mul2_0_0_n58), .ZN(
        s5_mul2_0_0_n54) );
  XOR2_X1 s5_mul2_0_0_U7 ( .A(stage4Out[1]), .B(stage4Out[3]), .Z(
        s5_mul2_0_0_n58) );
  XOR2_X1 s5_mul2_0_0_U6 ( .A(s5_n2), .B(s5_n4), .Z(s5_mul2_0_0_n61) );
  NOR2_X1 s5_mul2_0_0_U5 ( .A1(s5_mul2_0_0_n63), .A2(s5_mul2_0_0_n60), .ZN(
        s5_mul2_0_0_n55) );
  XNOR2_X1 s5_mul2_0_0_U4 ( .A(s5_n1), .B(s5_n3), .ZN(s5_mul2_0_0_n60) );
  XNOR2_X1 s5_mul2_0_0_U3 ( .A(stage4Out[0]), .B(stage4Out[2]), .ZN(
        s5_mul2_0_0_n63) );
  AOI221_X1 s5_mul2_0_0_U2 ( .B1(stage4Out[0]), .B2(stage4Out[1]), .C1(s5_n1), 
        .C2(s5_n2), .A(s5_mul2_0_0_n53), .ZN(s5_mul2_0_0_n66) );
  OAI22_X1 s5_mul2_0_0_U1 ( .A1(stage4Out[0]), .A2(stage4Out[1]), .B1(s5_n2), 
        .B2(s5_n1), .ZN(s5_mul2_0_0_n53) );
  XOR2_X1 s5_compr_0_0_U8 ( .A(s5_regOut[7]), .B(s5_regOut[15]), .Z(
        s5_chain_0__1__7_) );
  XOR2_X1 s5_compr_0_0_U7 ( .A(s5_regOut[6]), .B(s5_regOut[14]), .Z(
        s5_chain_0__1__6_) );
  XOR2_X1 s5_compr_0_0_U6 ( .A(s5_regOut[5]), .B(s5_regOut[13]), .Z(
        s5_chain_0__1__5_) );
  XOR2_X1 s5_compr_0_0_U5 ( .A(s5_regOut[4]), .B(s5_regOut[12]), .Z(
        s5_chain_0__1__4_) );
  XOR2_X1 s5_compr_0_0_U4 ( .A(s5_regOut[3]), .B(s5_regOut[11]), .Z(
        s5_chain_0__1__3_) );
  XOR2_X1 s5_compr_0_0_U3 ( .A(s5_regOut[2]), .B(s5_regOut[10]), .Z(
        s5_chain_0__1__2_) );
  XOR2_X1 s5_compr_0_0_U2 ( .A(s5_regOut[1]), .B(s5_regOut[9]), .Z(
        s5_chain_0__1__1_) );
  XOR2_X1 s5_compr_0_0_U1 ( .A(s5_regOut[0]), .B(s5_regOut[8]), .Z(
        s5_chain_0__1__0_) );
  XOR2_X1 s5_compr_0_1_U8 ( .A(s5_chain_0__1__7_), .B(s5_regOut[23]), .Z(
        stage5Out[7]) );
  XOR2_X1 s5_compr_0_1_U7 ( .A(s5_chain_0__1__6_), .B(s5_regOut[22]), .Z(
        stage5Out[6]) );
  XOR2_X1 s5_compr_0_1_U6 ( .A(s5_chain_0__1__5_), .B(s5_regOut[21]), .Z(
        stage5Out[5]) );
  XOR2_X1 s5_compr_0_1_U5 ( .A(s5_chain_0__1__4_), .B(s5_regOut[20]), .Z(
        stage5Out[4]) );
  XOR2_X1 s5_compr_0_1_U4 ( .A(s5_chain_0__1__3_), .B(s5_regOut[19]), .Z(
        stage5Out[3]) );
  XOR2_X1 s5_compr_0_1_U3 ( .A(s5_chain_0__1__2_), .B(s5_regOut[18]), .Z(
        stage5Out[2]) );
  XOR2_X1 s5_compr_0_1_U2 ( .A(s5_chain_0__1__1_), .B(s5_regOut[17]), .Z(
        stage5Out[1]) );
  XOR2_X1 s5_compr_0_1_U1 ( .A(s5_chain_0__1__0_), .B(s5_regOut[16]), .Z(
        stage5Out[0]) );
  XOR2_X1 s5_compr_1_0_U8 ( .A(s5_regOut[31]), .B(s5_regOut[39]), .Z(
        s5_chain_1__1__7_) );
  XOR2_X1 s5_compr_1_0_U7 ( .A(s5_regOut[30]), .B(s5_regOut[38]), .Z(
        s5_chain_1__1__6_) );
  XOR2_X1 s5_compr_1_0_U6 ( .A(s5_regOut[29]), .B(s5_regOut[37]), .Z(
        s5_chain_1__1__5_) );
  XOR2_X1 s5_compr_1_0_U5 ( .A(s5_regOut[28]), .B(s5_regOut[36]), .Z(
        s5_chain_1__1__4_) );
  XOR2_X1 s5_compr_1_0_U4 ( .A(s5_regOut[27]), .B(s5_regOut[35]), .Z(
        s5_chain_1__1__3_) );
  XOR2_X1 s5_compr_1_0_U3 ( .A(s5_regOut[26]), .B(s5_regOut[34]), .Z(
        s5_chain_1__1__2_) );
  XOR2_X1 s5_compr_1_0_U2 ( .A(s5_regOut[25]), .B(s5_regOut[33]), .Z(
        s5_chain_1__1__1_) );
  XOR2_X1 s5_compr_1_0_U1 ( .A(s5_regOut[24]), .B(s5_regOut[32]), .Z(
        s5_chain_1__1__0_) );
  XOR2_X1 s5_compr_1_1_U8 ( .A(s5_chain_1__1__7_), .B(s5_regOut[47]), .Z(
        stage5Out[15]) );
  XOR2_X1 s5_compr_1_1_U7 ( .A(s5_chain_1__1__6_), .B(s5_regOut[46]), .Z(
        stage5Out[14]) );
  XOR2_X1 s5_compr_1_1_U6 ( .A(s5_chain_1__1__5_), .B(s5_regOut[45]), .Z(
        stage5Out[13]) );
  XOR2_X1 s5_compr_1_1_U5 ( .A(s5_chain_1__1__4_), .B(s5_regOut[44]), .Z(
        stage5Out[12]) );
  XOR2_X1 s5_compr_1_1_U4 ( .A(s5_chain_1__1__3_), .B(s5_regOut[43]), .Z(
        stage5Out[11]) );
  XOR2_X1 s5_compr_1_1_U3 ( .A(s5_chain_1__1__2_), .B(s5_regOut[42]), .Z(
        stage5Out[10]) );
  XOR2_X1 s5_compr_1_1_U2 ( .A(s5_chain_1__1__1_), .B(s5_regOut[41]), .Z(
        stage5Out[9]) );
  XOR2_X1 s5_compr_1_1_U1 ( .A(s5_chain_1__1__0_), .B(s5_regOut[40]), .Z(
        stage5Out[8]) );
  XOR2_X1 s5_compr_2_0_U8 ( .A(s5_regOut[55]), .B(s5_regOut[63]), .Z(
        s5_chain_2__1__7_) );
  XOR2_X1 s5_compr_2_0_U7 ( .A(s5_regOut[54]), .B(s5_regOut[62]), .Z(
        s5_chain_2__1__6_) );
  XOR2_X1 s5_compr_2_0_U6 ( .A(s5_regOut[53]), .B(s5_regOut[61]), .Z(
        s5_chain_2__1__5_) );
  XOR2_X1 s5_compr_2_0_U5 ( .A(s5_regOut[52]), .B(s5_regOut[60]), .Z(
        s5_chain_2__1__4_) );
  XOR2_X1 s5_compr_2_0_U4 ( .A(s5_regOut[51]), .B(s5_regOut[59]), .Z(
        s5_chain_2__1__3_) );
  XOR2_X1 s5_compr_2_0_U3 ( .A(s5_regOut[50]), .B(s5_regOut[58]), .Z(
        s5_chain_2__1__2_) );
  XOR2_X1 s5_compr_2_0_U2 ( .A(s5_regOut[49]), .B(s5_regOut[57]), .Z(
        s5_chain_2__1__1_) );
  XOR2_X1 s5_compr_2_0_U1 ( .A(s5_regOut[48]), .B(s5_regOut[56]), .Z(
        s5_chain_2__1__0_) );
  XOR2_X1 s5_compr_2_1_U8 ( .A(s5_chain_2__1__7_), .B(s5_regOut[71]), .Z(
        stage5Out[23]) );
  XOR2_X1 s5_compr_2_1_U7 ( .A(s5_chain_2__1__6_), .B(s5_regOut[70]), .Z(
        stage5Out[22]) );
  XOR2_X1 s5_compr_2_1_U6 ( .A(s5_chain_2__1__5_), .B(s5_regOut[69]), .Z(
        stage5Out[21]) );
  XOR2_X1 s5_compr_2_1_U5 ( .A(s5_chain_2__1__4_), .B(s5_regOut[68]), .Z(
        stage5Out[20]) );
  XOR2_X1 s5_compr_2_1_U4 ( .A(s5_chain_2__1__3_), .B(s5_regOut[67]), .Z(
        stage5Out[19]) );
  XOR2_X1 s5_compr_2_1_U3 ( .A(s5_chain_2__1__2_), .B(s5_regOut[66]), .Z(
        stage5Out[18]) );
  XOR2_X1 s5_compr_2_1_U2 ( .A(s5_chain_2__1__1_), .B(s5_regOut[65]), .Z(
        stage5Out[17]) );
  XOR2_X1 s5_compr_2_1_U1 ( .A(s5_chain_2__1__0_), .B(s5_regOut[64]), .Z(
        stage5Out[16]) );
  XOR2_X1 s6_2_U11 ( .A(stage5Out[19]), .B(stage5Out[23]), .Z(stage6Out[22])
         );
  XNOR2_X1 s6_2_U10 ( .A(stage6Out[20]), .B(s6_2_n9), .ZN(stage6Out[19]) );
  XOR2_X1 s6_2_U9 ( .A(stage6Out[23]), .B(stage5Out[23]), .Z(stage6Out[20]) );
  XNOR2_X1 s6_2_U8 ( .A(s6_2_n8), .B(stage6Out[21]), .ZN(stage6Out[18]) );
  XNOR2_X1 s6_2_U7 ( .A(stage6Out[23]), .B(stage5Out[18]), .ZN(s6_2_n8) );
  XOR2_X1 s6_2_U6 ( .A(stage5Out[22]), .B(stage5Out[16]), .Z(stage6Out[21]) );
  XOR2_X1 s6_2_U5 ( .A(stage5Out[19]), .B(stage5Out[21]), .Z(stage6Out[23]) );
  XNOR2_X1 s6_2_U4 ( .A(s6_2_n7), .B(stage5Out[17]), .ZN(stage6Out[17]) );
  XNOR2_X1 s6_2_U3 ( .A(stage5Out[21]), .B(stage5Out[20]), .ZN(s6_2_n7) );
  XNOR2_X1 s6_2_U2 ( .A(stage5Out[17]), .B(s6_2_n9), .ZN(stage6Out[16]) );
  XNOR2_X1 s6_2_U1 ( .A(stage5Out[22]), .B(stage5Out[20]), .ZN(s6_2_n9) );
  XOR2_X1 s6_1_U11 ( .A(stage5Out[11]), .B(stage5Out[15]), .Z(stage6Out[14])
         );
  XNOR2_X1 s6_1_U10 ( .A(stage6Out[12]), .B(s6_1_n9), .ZN(stage6Out[11]) );
  XOR2_X1 s6_1_U9 ( .A(stage6Out[15]), .B(stage5Out[15]), .Z(stage6Out[12]) );
  XNOR2_X1 s6_1_U8 ( .A(s6_1_n8), .B(stage6Out[13]), .ZN(stage6Out[10]) );
  XNOR2_X1 s6_1_U7 ( .A(stage6Out[15]), .B(stage5Out[10]), .ZN(s6_1_n8) );
  XOR2_X1 s6_1_U6 ( .A(stage5Out[14]), .B(stage5Out[8]), .Z(stage6Out[13]) );
  XOR2_X1 s6_1_U5 ( .A(stage5Out[11]), .B(stage5Out[13]), .Z(stage6Out[15]) );
  XNOR2_X1 s6_1_U4 ( .A(s6_1_n7), .B(stage5Out[9]), .ZN(stage6Out[9]) );
  XNOR2_X1 s6_1_U3 ( .A(stage5Out[13]), .B(stage5Out[12]), .ZN(s6_1_n7) );
  XNOR2_X1 s6_1_U2 ( .A(stage5Out[9]), .B(s6_1_n9), .ZN(stage6Out[8]) );
  XNOR2_X1 s6_1_U1 ( .A(stage5Out[14]), .B(stage5Out[12]), .ZN(s6_1_n9) );
  XOR2_X1 s6_0_U11 ( .A(stage5Out[3]), .B(stage5Out[7]), .Z(stage6Out[6]) );
  XNOR2_X1 s6_0_U10 ( .A(stage6Out[4]), .B(s6_0_n9), .ZN(stage6Out[3]) );
  XOR2_X1 s6_0_U9 ( .A(stage6Out[7]), .B(stage5Out[7]), .Z(stage6Out[4]) );
  XNOR2_X1 s6_0_U8 ( .A(s6_0_n8), .B(stage6Out[5]), .ZN(stage6Out[2]) );
  XNOR2_X1 s6_0_U7 ( .A(stage6Out[7]), .B(stage5Out[2]), .ZN(s6_0_n8) );
  XOR2_X1 s6_0_U6 ( .A(stage5Out[6]), .B(stage5Out[0]), .Z(stage6Out[5]) );
  XOR2_X1 s6_0_U5 ( .A(stage5Out[3]), .B(stage5Out[5]), .Z(stage6Out[7]) );
  XNOR2_X1 s6_0_U4 ( .A(s6_0_n7), .B(stage5Out[1]), .ZN(stage6Out[1]) );
  XNOR2_X1 s6_0_U3 ( .A(stage5Out[5]), .B(stage5Out[4]), .ZN(s6_0_n7) );
  XNOR2_X1 s6_0_U2 ( .A(stage5Out[1]), .B(s6_0_n9), .ZN(stage6Out[0]) );
  XNOR2_X1 s6_0_U1 ( .A(stage5Out[6]), .B(stage5Out[4]), .ZN(s6_0_n9) );
endmodule

