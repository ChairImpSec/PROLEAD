
module circuit ( Clock, Reset, InData, FreshRand, Ready, OutData );
  input [49:0] InData;
  input [24:0] FreshRand;
  output [49:0] OutData;
  input Clock, Reset;
  output Ready;
  wire   Lastround, IotaRC_0_, n2, all_mux_linear_0__MUX_theta_state_inst_n217,
         all_mux_linear_0__MUX_theta_state_inst_n216,
         all_mux_linear_0__MUX_theta_state_inst_n215,
         all_mux_linear_0__MUX_theta_state_inst_n214,
         all_mux_linear_0__MUX_theta_state_inst_n213,
         all_mux_linear_0__MUX_theta_state_inst_n212,
         all_mux_linear_0__MUX_theta_state_inst_n211,
         all_mux_linear_0__MUX_theta_state_inst_n210,
         all_mux_linear_0__MUX_theta_state_inst_n209,
         all_mux_linear_0__MUX_theta_state_inst_n208,
         all_mux_linear_0__MUX_theta_state_inst_n207,
         all_mux_linear_0__MUX_theta_state_inst_n206,
         all_mux_linear_0__MUX_theta_state_inst_n205,
         all_mux_linear_0__MUX_theta_state_inst_n204,
         all_mux_linear_0__MUX_theta_state_inst_n203,
         all_mux_linear_0__MUX_theta_state_inst_n202,
         all_mux_linear_0__MUX_theta_state_inst_n201,
         all_mux_linear_0__MUX_theta_state_inst_n200,
         all_mux_linear_0__MUX_theta_state_inst_n199,
         all_mux_linear_0__MUX_theta_state_inst_n198,
         all_mux_linear_0__MUX_theta_state_inst_n197,
         all_mux_linear_0__MUX_theta_state_inst_n196,
         all_mux_linear_0__MUX_theta_state_inst_n195,
         all_mux_linear_0__MUX_theta_state_inst_n194,
         all_mux_linear_0__MUX_theta_state_inst_n193,
         all_mux_linear_0__MUX_theta_state_inst_n192,
         all_mux_linear_0__MUX_theta_state_inst_n191,
         all_mux_linear_0__MUX_theta_state_inst_n190,
         all_mux_linear_0__MUX_theta_state_inst_n189,
         all_mux_linear_0__MUX_theta_state_inst_n188,
         all_mux_linear_0__MUX_theta_state_inst_n187,
         all_mux_linear_0__MUX_theta_state_inst_n186,
         all_mux_linear_0__MUX_theta_state_inst_n185,
         all_mux_linear_0__MUX_theta_state_inst_n184,
         all_mux_linear_0__MUX_theta_state_inst_n183,
         all_mux_linear_0__MUX_theta_state_inst_n182,
         all_mux_linear_0__MUX_theta_state_inst_n181,
         all_mux_linear_0__MUX_theta_state_inst_n180,
         all_mux_linear_0__MUX_theta_state_inst_n179,
         all_mux_linear_0__MUX_theta_state_inst_n178,
         all_mux_linear_0__MUX_theta_state_inst_n177,
         all_mux_linear_0__MUX_theta_state_inst_n176,
         all_mux_linear_0__MUX_theta_state_inst_n175,
         all_mux_linear_0__MUX_theta_state_inst_n174,
         all_mux_linear_0__MUX_theta_state_inst_n173,
         all_mux_linear_0__MUX_theta_state_inst_n172,
         all_mux_linear_0__MUX_theta_state_inst_n171,
         all_mux_linear_0__MUX_theta_state_inst_n170,
         all_mux_linear_0__MUX_theta_state_inst_n169,
         all_mux_linear_0__MUX_theta_state_inst_n168,
         all_mux_linear_0__MUX_theta_state_inst_n167,
         all_mux_linear_0__MUX_theta_state_inst_n166,
         all_mux_linear_0__MUX_theta_state_inst_n165,
         all_mux_linear_0__MUX_theta_state_inst_n164,
         all_mux_linear_0__MUX_theta_state_inst_n163,
         all_mux_linear_0__MUX_theta_state_inst_n162,
         all_mux_linear_0__MUX_theta_state_inst_n161,
         all_mux_linear_0__MUX_theta_state_inst_n160,
         all_mux_linear_0__MUX_theta_state_inst_n159,
         all_mux_linear_0__MUX_theta_state_inst_n158,
         all_mux_linear_0__MUX_theta_state_inst_n157,
         all_mux_linear_0__MUX_theta_state_inst_n156,
         all_mux_linear_0__MUX_theta_state_inst_n155,
         all_mux_linear_0__MUX_theta_state_inst_n154,
         all_mux_linear_0__MUX_theta_state_inst_n153,
         all_mux_linear_0__MUX_theta_state_inst_n152,
         all_mux_linear_0__MUX_theta_state_inst_n151,
         all_mux_linear_0__MUX_theta_state_inst_n150,
         all_mux_linear_0__MUX_theta_state_inst_n149,
         all_mux_linear_0__MUX_theta_state_inst_n148,
         all_mux_linear_0__MUX_theta_state_inst_n147,
         all_mux_linear_0__MUX_theta_state_inst_n146,
         all_mux_linear_0__MUX_theta_state_inst_n145,
         all_mux_linear_0__MUX_theta_state_inst_n144,
         all_mux_linear_0__MUX_theta_state_inst_n143,
         all_mux_linear_0__MUX_theta_state_inst_n142,
         all_mux_linear_0__MUX_theta_state_inst_n141,
         all_mux_linear_0__MUX_theta_state_inst_n140,
         all_mux_linear_0__MUX_theta_state_inst_n139,
         all_mux_linear_0__MUX_theta_state_inst_n138,
         all_mux_linear_0__MUX_theta_state_inst_n137,
         all_mux_linear_0__MUX_theta_state_inst_n136,
         all_mux_linear_0__MUX_theta_state_inst_n135,
         all_mux_linear_0__MUX_theta_state_inst_n134,
         all_mux_linear_0__MUX_theta_state_inst_n133,
         all_mux_linear_0__MUX_theta_state_inst_n132,
         all_mux_linear_0__MUX_theta_state_inst_n131,
         all_mux_linear_0__MUX_theta_state_inst_n130,
         all_mux_linear_0__MUX_theta_state_inst_n129,
         all_mux_linear_1__MUX_theta_state_inst_n335,
         all_mux_linear_1__MUX_theta_state_inst_n334,
         all_mux_linear_1__MUX_theta_state_inst_n333,
         all_mux_linear_1__MUX_theta_state_inst_n332,
         all_mux_linear_1__MUX_theta_state_inst_n331,
         all_mux_linear_1__MUX_theta_state_inst_n330,
         all_mux_linear_1__MUX_theta_state_inst_n329,
         all_mux_linear_1__MUX_theta_state_inst_n328,
         all_mux_linear_1__MUX_theta_state_inst_n327,
         all_mux_linear_1__MUX_theta_state_inst_n326,
         all_mux_linear_1__MUX_theta_state_inst_n325,
         all_mux_linear_1__MUX_theta_state_inst_n324,
         all_mux_linear_1__MUX_theta_state_inst_n323,
         all_mux_linear_1__MUX_theta_state_inst_n322,
         all_mux_linear_1__MUX_theta_state_inst_n321,
         all_mux_linear_1__MUX_theta_state_inst_n320,
         all_mux_linear_1__MUX_theta_state_inst_n319,
         all_mux_linear_1__MUX_theta_state_inst_n318,
         all_mux_linear_1__MUX_theta_state_inst_n317,
         all_mux_linear_1__MUX_theta_state_inst_n316,
         all_mux_linear_1__MUX_theta_state_inst_n315,
         all_mux_linear_1__MUX_theta_state_inst_n314,
         all_mux_linear_1__MUX_theta_state_inst_n313,
         all_mux_linear_1__MUX_theta_state_inst_n312,
         all_mux_linear_1__MUX_theta_state_inst_n311,
         all_mux_linear_1__MUX_theta_state_inst_n310,
         all_mux_linear_1__MUX_theta_state_inst_n309,
         all_mux_linear_1__MUX_theta_state_inst_n308,
         all_mux_linear_1__MUX_theta_state_inst_n307,
         all_mux_linear_1__MUX_theta_state_inst_n306,
         all_mux_linear_1__MUX_theta_state_inst_n305,
         all_mux_linear_1__MUX_theta_state_inst_n304,
         all_mux_linear_1__MUX_theta_state_inst_n303,
         all_mux_linear_1__MUX_theta_state_inst_n302,
         all_mux_linear_1__MUX_theta_state_inst_n301,
         all_mux_linear_1__MUX_theta_state_inst_n300,
         all_mux_linear_1__MUX_theta_state_inst_n299,
         all_mux_linear_1__MUX_theta_state_inst_n298,
         all_mux_linear_1__MUX_theta_state_inst_n297,
         all_mux_linear_1__MUX_theta_state_inst_n296,
         all_mux_linear_1__MUX_theta_state_inst_n295,
         all_mux_linear_1__MUX_theta_state_inst_n294,
         all_mux_linear_1__MUX_theta_state_inst_n293,
         all_mux_linear_1__MUX_theta_state_inst_n292,
         all_mux_linear_1__MUX_theta_state_inst_n291,
         all_mux_linear_1__MUX_theta_state_inst_n290,
         all_mux_linear_1__MUX_theta_state_inst_n289,
         all_mux_linear_1__MUX_theta_state_inst_n288,
         all_mux_linear_1__MUX_theta_state_inst_n287,
         all_mux_linear_1__MUX_theta_state_inst_n286,
         all_mux_linear_1__MUX_theta_state_inst_n285,
         all_mux_linear_1__MUX_theta_state_inst_n284,
         all_mux_linear_1__MUX_theta_state_inst_n283,
         all_mux_linear_1__MUX_theta_state_inst_n282,
         all_mux_linear_1__MUX_theta_state_inst_n281,
         all_mux_linear_1__MUX_theta_state_inst_n280,
         all_mux_linear_1__MUX_theta_state_inst_n279,
         all_mux_linear_1__MUX_theta_state_inst_n278,
         all_mux_linear_1__MUX_theta_state_inst_n277,
         all_mux_linear_1__MUX_theta_state_inst_n276,
         all_mux_linear_1__MUX_theta_state_inst_n275,
         all_mux_linear_1__MUX_theta_state_inst_n274,
         all_mux_linear_1__MUX_theta_state_inst_n273,
         all_mux_linear_1__MUX_theta_state_inst_n272,
         all_mux_linear_1__MUX_theta_state_inst_n271,
         all_mux_linear_1__MUX_theta_state_inst_n270,
         all_mux_linear_1__MUX_theta_state_inst_n269,
         all_mux_linear_1__MUX_theta_state_inst_n268,
         all_mux_linear_1__MUX_theta_state_inst_n267,
         all_mux_linear_1__MUX_theta_state_inst_n266,
         all_mux_linear_1__MUX_theta_state_inst_n265,
         all_mux_linear_1__MUX_theta_state_inst_n264,
         all_mux_linear_1__MUX_theta_state_inst_n263,
         all_mux_linear_1__MUX_theta_state_inst_n262,
         all_mux_linear_1__MUX_theta_state_inst_n261,
         all_mux_linear_1__MUX_theta_state_inst_n260,
         all_mux_linear_1__MUX_theta_state_inst_n259,
         all_mux_linear_1__MUX_theta_state_inst_n258,
         all_mux_linear_1__MUX_theta_state_inst_n257,
         all_mux_linear_1__MUX_theta_state_inst_n256,
         all_mux_linear_1__MUX_theta_state_inst_n255,
         all_mux_linear_1__MUX_theta_state_inst_n254,
         all_mux_linear_1__MUX_theta_state_inst_n253,
         all_mux_linear_1__MUX_theta_state_inst_n252,
         all_mux_linear_1__MUX_theta_state_inst_n251,
         all_mux_linear_1__MUX_theta_state_inst_n250,
         all_mux_linear_1__MUX_theta_state_inst_n249,
         all_mux_linear_1__MUX_theta_state_inst_n248,
         all_mux_linear_1__MUX_theta_state_inst_n247,
         all_mux_linear_1__MUX_theta_state_inst_n246,
         all_mux_linear_1__MUX_theta_state_inst_n245,
         all_mux_linear_1__MUX_theta_state_inst_n244,
         all_mux_linear_1__MUX_theta_state_inst_n243,
         all_mux_linear_1__MUX_theta_state_inst_n242,
         all_mux_linear_1__MUX_theta_state_inst_n241,
         all_mux_linear_1__MUX_theta_state_inst_n240,
         all_mux_linear_1__MUX_theta_state_inst_n239,
         all_mux_linear_1__MUX_theta_state_inst_n238,
         all_mux_linear_1__MUX_theta_state_inst_n237,
         all_mux_linear_1__MUX_theta_state_inst_n236,
         all_mux_linear_1__MUX_theta_state_inst_n235,
         all_mux_linear_1__MUX_theta_state_inst_n234,
         all_mux_linear_1__MUX_theta_state_inst_n233,
         all_mux_linear_1__MUX_theta_state_inst_n232,
         all_mux_linear_1__MUX_theta_state_inst_n231,
         all_mux_linear_1__MUX_theta_state_inst_n230,
         all_mux_linear_1__MUX_theta_state_inst_n229,
         all_mux_linear_2__MUX_theta_state_inst_n335,
         all_mux_linear_2__MUX_theta_state_inst_n334,
         all_mux_linear_2__MUX_theta_state_inst_n333,
         all_mux_linear_2__MUX_theta_state_inst_n332,
         all_mux_linear_2__MUX_theta_state_inst_n331,
         all_mux_linear_2__MUX_theta_state_inst_n330,
         all_mux_linear_2__MUX_theta_state_inst_n329,
         all_mux_linear_2__MUX_theta_state_inst_n328,
         all_mux_linear_2__MUX_theta_state_inst_n327,
         all_mux_linear_2__MUX_theta_state_inst_n326,
         all_mux_linear_2__MUX_theta_state_inst_n325,
         all_mux_linear_2__MUX_theta_state_inst_n324,
         all_mux_linear_2__MUX_theta_state_inst_n323,
         all_mux_linear_2__MUX_theta_state_inst_n322,
         all_mux_linear_2__MUX_theta_state_inst_n321,
         all_mux_linear_2__MUX_theta_state_inst_n320,
         all_mux_linear_2__MUX_theta_state_inst_n319,
         all_mux_linear_2__MUX_theta_state_inst_n318,
         all_mux_linear_2__MUX_theta_state_inst_n317,
         all_mux_linear_2__MUX_theta_state_inst_n316,
         all_mux_linear_2__MUX_theta_state_inst_n315,
         all_mux_linear_2__MUX_theta_state_inst_n314,
         all_mux_linear_2__MUX_theta_state_inst_n313,
         all_mux_linear_2__MUX_theta_state_inst_n312,
         all_mux_linear_2__MUX_theta_state_inst_n311,
         all_mux_linear_2__MUX_theta_state_inst_n310,
         all_mux_linear_2__MUX_theta_state_inst_n309,
         all_mux_linear_2__MUX_theta_state_inst_n308,
         all_mux_linear_2__MUX_theta_state_inst_n307,
         all_mux_linear_2__MUX_theta_state_inst_n306,
         all_mux_linear_2__MUX_theta_state_inst_n305,
         all_mux_linear_2__MUX_theta_state_inst_n304,
         all_mux_linear_2__MUX_theta_state_inst_n303,
         all_mux_linear_2__MUX_theta_state_inst_n302,
         all_mux_linear_2__MUX_theta_state_inst_n301,
         all_mux_linear_2__MUX_theta_state_inst_n300,
         all_mux_linear_2__MUX_theta_state_inst_n299,
         all_mux_linear_2__MUX_theta_state_inst_n298,
         all_mux_linear_2__MUX_theta_state_inst_n297,
         all_mux_linear_2__MUX_theta_state_inst_n296,
         all_mux_linear_2__MUX_theta_state_inst_n295,
         all_mux_linear_2__MUX_theta_state_inst_n294,
         all_mux_linear_2__MUX_theta_state_inst_n293,
         all_mux_linear_2__MUX_theta_state_inst_n292,
         all_mux_linear_2__MUX_theta_state_inst_n291,
         all_mux_linear_2__MUX_theta_state_inst_n290,
         all_mux_linear_2__MUX_theta_state_inst_n289,
         all_mux_linear_2__MUX_theta_state_inst_n288,
         all_mux_linear_2__MUX_theta_state_inst_n287,
         all_mux_linear_2__MUX_theta_state_inst_n286,
         all_mux_linear_2__MUX_theta_state_inst_n285,
         all_mux_linear_2__MUX_theta_state_inst_n284,
         all_mux_linear_2__MUX_theta_state_inst_n283,
         all_mux_linear_2__MUX_theta_state_inst_n282,
         all_mux_linear_2__MUX_theta_state_inst_n281,
         all_mux_linear_2__MUX_theta_state_inst_n280,
         all_mux_linear_2__MUX_theta_state_inst_n279,
         all_mux_linear_2__MUX_theta_state_inst_n278,
         all_mux_linear_2__MUX_theta_state_inst_n277,
         all_mux_linear_2__MUX_theta_state_inst_n276,
         all_mux_linear_2__MUX_theta_state_inst_n275,
         all_mux_linear_2__MUX_theta_state_inst_n274,
         all_mux_linear_2__MUX_theta_state_inst_n273,
         all_mux_linear_2__MUX_theta_state_inst_n272,
         all_mux_linear_2__MUX_theta_state_inst_n271,
         all_mux_linear_2__MUX_theta_state_inst_n270,
         all_mux_linear_2__MUX_theta_state_inst_n269,
         all_mux_linear_2__MUX_theta_state_inst_n268,
         all_mux_linear_2__MUX_theta_state_inst_n267,
         all_mux_linear_2__MUX_theta_state_inst_n266,
         all_mux_linear_2__MUX_theta_state_inst_n265,
         all_mux_linear_2__MUX_theta_state_inst_n264,
         all_mux_linear_2__MUX_theta_state_inst_n263,
         all_mux_linear_2__MUX_theta_state_inst_n262,
         all_mux_linear_2__MUX_theta_state_inst_n261,
         all_mux_linear_2__MUX_theta_state_inst_n260,
         all_mux_linear_2__MUX_theta_state_inst_n259,
         all_mux_linear_2__MUX_theta_state_inst_n258,
         all_mux_linear_2__MUX_theta_state_inst_n257,
         all_mux_linear_2__MUX_theta_state_inst_n256,
         all_mux_linear_2__MUX_theta_state_inst_n255,
         all_mux_linear_2__MUX_theta_state_inst_n254,
         all_mux_linear_2__MUX_theta_state_inst_n253,
         all_mux_linear_2__MUX_theta_state_inst_n252,
         all_mux_linear_2__MUX_theta_state_inst_n251,
         all_mux_linear_2__MUX_theta_state_inst_n250,
         all_mux_linear_2__MUX_theta_state_inst_n249,
         all_mux_linear_2__MUX_theta_state_inst_n248,
         all_mux_linear_2__MUX_theta_state_inst_n247,
         all_mux_linear_2__MUX_theta_state_inst_n246,
         all_mux_linear_2__MUX_theta_state_inst_n245,
         all_mux_linear_2__MUX_theta_state_inst_n244,
         all_mux_linear_2__MUX_theta_state_inst_n243,
         all_mux_linear_2__MUX_theta_state_inst_n242,
         all_mux_linear_2__MUX_theta_state_inst_n241,
         all_mux_linear_2__MUX_theta_state_inst_n240,
         all_mux_linear_2__MUX_theta_state_inst_n239,
         all_mux_linear_2__MUX_theta_state_inst_n238,
         all_mux_linear_2__MUX_theta_state_inst_n237,
         all_mux_linear_2__MUX_theta_state_inst_n236,
         all_mux_linear_2__MUX_theta_state_inst_n235,
         all_mux_linear_2__MUX_theta_state_inst_n234,
         all_mux_linear_2__MUX_theta_state_inst_n233,
         all_mux_linear_2__MUX_theta_state_inst_n232,
         all_mux_linear_2__MUX_theta_state_inst_n231,
         all_mux_linear_2__MUX_theta_state_inst_n230,
         all_mux_linear_2__MUX_theta_state_inst_n229,
         all_mux_linear_3__MUX_theta_state_inst_n318,
         all_mux_linear_3__MUX_theta_state_inst_n317,
         all_mux_linear_3__MUX_theta_state_inst_n316,
         all_mux_linear_3__MUX_theta_state_inst_n315,
         all_mux_linear_3__MUX_theta_state_inst_n314,
         all_mux_linear_3__MUX_theta_state_inst_n313,
         all_mux_linear_3__MUX_theta_state_inst_n312,
         all_mux_linear_3__MUX_theta_state_inst_n311,
         all_mux_linear_3__MUX_theta_state_inst_n310,
         all_mux_linear_3__MUX_theta_state_inst_n309,
         all_mux_linear_3__MUX_theta_state_inst_n308,
         all_mux_linear_3__MUX_theta_state_inst_n307,
         all_mux_linear_3__MUX_theta_state_inst_n306,
         all_mux_linear_3__MUX_theta_state_inst_n305,
         all_mux_linear_3__MUX_theta_state_inst_n304,
         all_mux_linear_3__MUX_theta_state_inst_n303,
         all_mux_linear_3__MUX_theta_state_inst_n302,
         all_mux_linear_3__MUX_theta_state_inst_n301,
         all_mux_linear_3__MUX_theta_state_inst_n300,
         all_mux_linear_3__MUX_theta_state_inst_n299,
         all_mux_linear_3__MUX_theta_state_inst_n298,
         all_mux_linear_3__MUX_theta_state_inst_n297,
         all_mux_linear_3__MUX_theta_state_inst_n296,
         all_mux_linear_3__MUX_theta_state_inst_n295,
         all_mux_linear_3__MUX_theta_state_inst_n294,
         all_mux_linear_3__MUX_theta_state_inst_n293,
         all_mux_linear_3__MUX_theta_state_inst_n292,
         all_mux_linear_3__MUX_theta_state_inst_n291,
         all_mux_linear_3__MUX_theta_state_inst_n290,
         all_mux_linear_3__MUX_theta_state_inst_n289,
         all_mux_linear_3__MUX_theta_state_inst_n288,
         all_mux_linear_3__MUX_theta_state_inst_n287,
         all_mux_linear_3__MUX_theta_state_inst_n286,
         all_mux_linear_3__MUX_theta_state_inst_n285,
         all_mux_linear_3__MUX_theta_state_inst_n284,
         all_mux_linear_3__MUX_theta_state_inst_n283,
         all_mux_linear_3__MUX_theta_state_inst_n282,
         all_mux_linear_3__MUX_theta_state_inst_n281,
         all_mux_linear_3__MUX_theta_state_inst_n280,
         all_mux_linear_3__MUX_theta_state_inst_n279,
         all_mux_linear_3__MUX_theta_state_inst_n278,
         all_mux_linear_3__MUX_theta_state_inst_n277,
         all_mux_linear_3__MUX_theta_state_inst_n276,
         all_mux_linear_3__MUX_theta_state_inst_n275,
         all_mux_linear_3__MUX_theta_state_inst_n274,
         all_mux_linear_3__MUX_theta_state_inst_n273,
         all_mux_linear_3__MUX_theta_state_inst_n272,
         all_mux_linear_3__MUX_theta_state_inst_n271,
         all_mux_linear_3__MUX_theta_state_inst_n270,
         all_mux_linear_3__MUX_theta_state_inst_n269,
         all_mux_linear_3__MUX_theta_state_inst_n268,
         all_mux_linear_3__MUX_theta_state_inst_n267,
         all_mux_linear_3__MUX_theta_state_inst_n266,
         all_mux_linear_3__MUX_theta_state_inst_n265,
         all_mux_linear_3__MUX_theta_state_inst_n264,
         all_mux_linear_3__MUX_theta_state_inst_n263,
         all_mux_linear_3__MUX_theta_state_inst_n262,
         all_mux_linear_3__MUX_theta_state_inst_n261,
         all_mux_linear_3__MUX_theta_state_inst_n260,
         all_mux_linear_3__MUX_theta_state_inst_n259,
         all_mux_linear_3__MUX_theta_state_inst_n258,
         all_mux_linear_3__MUX_theta_state_inst_n257,
         all_mux_linear_3__MUX_theta_state_inst_n256,
         all_mux_linear_3__MUX_theta_state_inst_n255,
         all_mux_linear_3__MUX_theta_state_inst_n254,
         all_mux_linear_3__MUX_theta_state_inst_n253,
         all_mux_linear_3__MUX_theta_state_inst_n252,
         all_mux_linear_3__MUX_theta_state_inst_n251,
         all_mux_linear_3__MUX_theta_state_inst_n250,
         all_mux_linear_3__MUX_theta_state_inst_n249,
         all_mux_linear_3__MUX_theta_state_inst_n248,
         all_mux_linear_3__MUX_theta_state_inst_n247,
         all_mux_linear_3__MUX_theta_state_inst_n246,
         all_mux_linear_3__MUX_theta_state_inst_n245,
         all_mux_linear_3__MUX_theta_state_inst_n244,
         all_mux_linear_3__MUX_theta_state_inst_n243,
         all_mux_linear_3__MUX_theta_state_inst_n242,
         all_mux_linear_3__MUX_theta_state_inst_n241,
         all_mux_linear_3__MUX_theta_state_inst_n240,
         all_mux_linear_3__MUX_theta_state_inst_n239,
         all_mux_linear_3__MUX_theta_state_inst_n238,
         all_mux_linear_3__MUX_theta_state_inst_n237,
         all_mux_linear_3__MUX_theta_state_inst_n236,
         all_mux_linear_3__MUX_theta_state_inst_n235,
         all_mux_linear_3__MUX_theta_state_inst_n234,
         all_mux_linear_3__MUX_theta_state_inst_n233,
         all_mux_linear_3__MUX_theta_state_inst_n232,
         all_mux_linear_3__MUX_theta_state_inst_n231,
         all_mux_linear_3__MUX_theta_state_inst_n230, CHI_ChiOut_0_,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n2,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4,
         KECCAK_CONTROL_n62, KECCAK_CONTROL_n61, KECCAK_CONTROL_n60,
         KECCAK_CONTROL_n59, KECCAK_CONTROL_n58, KECCAK_CONTROL_n57,
         KECCAK_CONTROL_n56, KECCAK_CONTROL_n55, KECCAK_CONTROL_n54,
         KECCAK_CONTROL_n53, KECCAK_CONTROL_n52, KECCAK_CONTROL_n51,
         KECCAK_CONTROL_n50, KECCAK_CONTROL_n49, KECCAK_CONTROL_n48,
         KECCAK_CONTROL_n47, KECCAK_CONTROL_n46, KECCAK_CONTROL_n45,
         KECCAK_CONTROL_n44, KECCAK_CONTROL_n43, KECCAK_CONTROL_n42,
         KECCAK_CONTROL_n41, KECCAK_CONTROL_n40, KECCAK_CONTROL_n39,
         KECCAK_CONTROL_n38, KECCAK_CONTROL_n37, KECCAK_CONTROL_n36,
         KECCAK_CONTROL_n35, KECCAK_CONTROL_n34, KECCAK_CONTROL_n32,
         KECCAK_CONTROL_n31, KECCAK_CONTROL_n27, KECCAK_CONTROL_n26,
         KECCAK_CONTROL_n6, KECCAK_CONTROL_n29, KECCAK_CONTROL_n28,
         KECCAK_CONTROL_n15, KECCAK_CONTROL_n14, KECCAK_CONTROL_n5,
         KECCAK_CONTROL_N32, KECCAK_CONTROL_RoundCountxDP_0_,
         KECCAK_CONTROL_RoundCountxDP_1_, KECCAK_CONTROL_RoundCountxDP_2_,
         KECCAK_CONTROL_RoundCountxDP_3_, KECCAK_CONTROL_RoundCountxDP_4_,
         KECCAK_CONTROL_RC_GEN_n3, KECCAK_CONTROL_RC_GEN_n2;
  wire   [99:0] SlicesFromChi;
  wire   [99:0] StateOut;
  wire   [24:0] all_mux_linear_0__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_1__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_2__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_3__MUX_theta_state_inst_StateIn;

  BUF_X1 U2 ( .A(Lastround), .Z(n2) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U116 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n217), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n216), .A(
        all_mux_linear_0__MUX_theta_state_inst_n215), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U115 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[9]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n217), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n214), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n215) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U114 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n213), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n216), .A(
        all_mux_linear_0__MUX_theta_state_inst_n212), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U113 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[8]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n213), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n214), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n212) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U112 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n211), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n216), .A(
        all_mux_linear_0__MUX_theta_state_inst_n210), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U111 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[7]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n211), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n214), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n210) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U110 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n209), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n216), .A(
        all_mux_linear_0__MUX_theta_state_inst_n208), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U109 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[6]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n209), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n214), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n208) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U108 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n207), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n216), .A(
        all_mux_linear_0__MUX_theta_state_inst_n206), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U107 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[5]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n207), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n214), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n206) );
  NOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U106 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n205), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n214) );
  NAND2_X1 all_mux_linear_0__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n205), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n216) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U104 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n204), .B(
        all_mux_linear_0__MUX_theta_state_inst_n203), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n205) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U103 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n202), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n201), .A(
        all_mux_linear_0__MUX_theta_state_inst_n200), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[4]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U102 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[4]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n199), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n202), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n200) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U101 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n198), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n201), .A(
        all_mux_linear_0__MUX_theta_state_inst_n197), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[3]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U100 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[3]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n199), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n198), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n197) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U99 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n196), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n201), .A(
        all_mux_linear_0__MUX_theta_state_inst_n195), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[2]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U98 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[2]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n199), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n196), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n195) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U97 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n194), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n193), .A(
        all_mux_linear_0__MUX_theta_state_inst_n192), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[24]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U96 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[24]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n194), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n191), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n192) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n190), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n193), .A(
        all_mux_linear_0__MUX_theta_state_inst_n189), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[23]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[23]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n190), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n191), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n189) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U93 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n188), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n193), .A(
        all_mux_linear_0__MUX_theta_state_inst_n187), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[22]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U92 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[22]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n188), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n191), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n187) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n186), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n193), .A(
        all_mux_linear_0__MUX_theta_state_inst_n185), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[21]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[21]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n186), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n191), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n185) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U89 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n184), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n193), .A(
        all_mux_linear_0__MUX_theta_state_inst_n183), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[20]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U88 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[20]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n184), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n191), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n183) );
  NOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U87 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n182), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n191) );
  NAND2_X1 all_mux_linear_0__MUX_theta_state_inst_U86 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n182), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n193) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U85 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n181), .B(
        all_mux_linear_0__MUX_theta_state_inst_n203), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n182) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n180), .B(
        all_mux_linear_0__MUX_theta_state_inst_n179), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n203) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U83 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n178), .B(
        all_mux_linear_0__MUX_theta_state_inst_n177), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n179) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U82 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n176), .B(
        all_mux_linear_0__MUX_theta_state_inst_n202), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n177) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U81 ( .A1(Reset), .A2(
        InData[4]), .B1(SlicesFromChi[4]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n202) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U80 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n198), .B(
        all_mux_linear_0__MUX_theta_state_inst_n196), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n178) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U79 ( .A1(Reset), .A2(
        InData[2]), .B1(SlicesFromChi[2]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n196) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U78 ( .A1(Reset), .A2(
        InData[3]), .B1(SlicesFromChi[3]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n198) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n176), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n201), .A(
        all_mux_linear_0__MUX_theta_state_inst_n175), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[1]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[1]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n199), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n176), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n175) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U75 ( .A1(Reset), .A2(
        InData[1]), .B1(SlicesFromChi[1]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n176) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U74 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n174), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n173), .A(
        all_mux_linear_0__MUX_theta_state_inst_n172), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[19]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U73 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[19]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n174), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n171), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n172) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U72 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n170), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n173), .A(
        all_mux_linear_0__MUX_theta_state_inst_n169), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[18]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U71 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[18]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n170), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n171), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n169) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U70 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n168), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n173), .A(
        all_mux_linear_0__MUX_theta_state_inst_n167), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[17]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U69 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[17]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n168), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n171), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n167) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U68 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n166), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n173), .A(
        all_mux_linear_0__MUX_theta_state_inst_n165), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[16]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U67 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[16]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n166), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n171), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n165) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n164), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n173), .A(
        all_mux_linear_0__MUX_theta_state_inst_n163), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[15]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[15]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n164), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n171), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n163) );
  NOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U64 ( .A1(n2), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n162), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n171) );
  NAND2_X1 all_mux_linear_0__MUX_theta_state_inst_U63 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n162), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n173) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U62 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n161), .B(
        all_mux_linear_0__MUX_theta_state_inst_n204), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n162) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U61 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n160), .B(
        all_mux_linear_0__MUX_theta_state_inst_n159), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n204) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U60 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n158), .B(
        all_mux_linear_0__MUX_theta_state_inst_n157), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n159) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n156), .B(
        all_mux_linear_0__MUX_theta_state_inst_n155), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n157) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n154), .B(
        all_mux_linear_0__MUX_theta_state_inst_n153), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n158) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U57 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n154), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n152), .A(
        all_mux_linear_0__MUX_theta_state_inst_n151), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[14]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U56 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[14]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n150), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n154), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n151) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U55 ( .A1(Reset), .A2(
        InData[14]), .B1(SlicesFromChi[14]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n154) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n153), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n152), .A(
        all_mux_linear_0__MUX_theta_state_inst_n149), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[13]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[13]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n150), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n153), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n149) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U52 ( .A1(Reset), .A2(
        InData[13]), .B1(SlicesFromChi[13]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n153) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U51 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n155), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n152), .A(
        all_mux_linear_0__MUX_theta_state_inst_n148), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[12]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U50 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[12]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n150), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n155), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n148) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U49 ( .A1(Reset), .A2(
        InData[12]), .B1(SlicesFromChi[12]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n155) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U48 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n156), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n152), .A(
        all_mux_linear_0__MUX_theta_state_inst_n147), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[11]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U47 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[11]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n150), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n156), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n147) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U46 ( .A1(Reset), .A2(
        InData[11]), .B1(SlicesFromChi[11]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n156) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U45 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n160), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n152), .A(
        all_mux_linear_0__MUX_theta_state_inst_n146), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[10]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U44 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n129), .A2(SlicesFromChi[10]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n160), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n150), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n146) );
  NOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U43 ( .A1(n2), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n145), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n150) );
  NAND2_X1 all_mux_linear_0__MUX_theta_state_inst_U42 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n145), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n152) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U41 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n144), .B(
        all_mux_linear_0__MUX_theta_state_inst_n181), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n145) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U40 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n174), .B(
        all_mux_linear_0__MUX_theta_state_inst_n143), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n181) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U39 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n142), .B(
        all_mux_linear_0__MUX_theta_state_inst_n141), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n143) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U38 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n166), .B(
        all_mux_linear_0__MUX_theta_state_inst_n164), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n141) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U37 ( .A1(Reset), .A2(
        InData[15]), .B1(SlicesFromChi[15]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n164) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U36 ( .A1(Reset), .A2(
        InData[16]), .B1(SlicesFromChi[16]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n166) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n170), .B(
        all_mux_linear_0__MUX_theta_state_inst_n168), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n142) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U34 ( .A1(Reset), .A2(
        InData[17]), .B1(SlicesFromChi[17]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n168) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U33 ( .A1(Reset), .A2(
        InData[18]), .B1(SlicesFromChi[18]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n170) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U32 ( .A1(Reset), .A2(
        InData[19]), .B1(SlicesFromChi[19]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n174) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U31 ( .A1(Reset), .A2(
        InData[10]), .B1(SlicesFromChi[10]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n160) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U30 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n180), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n201), .A(
        all_mux_linear_0__MUX_theta_state_inst_n140), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[0]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[0]), 
        .A2(all_mux_linear_0__MUX_theta_state_inst_n129), .B1(
        all_mux_linear_0__MUX_theta_state_inst_n180), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n199), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n140) );
  NOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U28 ( .A1(n2), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n139), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n199) );
  NAND2_X1 all_mux_linear_0__MUX_theta_state_inst_U27 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n139), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n201) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U26 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n161), .B(
        all_mux_linear_0__MUX_theta_state_inst_n144), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n139) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U25 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n211), .B(
        all_mux_linear_0__MUX_theta_state_inst_n138), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n144) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n137), .B(
        all_mux_linear_0__MUX_theta_state_inst_n136), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n138) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U23 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n209), .B(
        all_mux_linear_0__MUX_theta_state_inst_n207), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n136) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U22 ( .A1(Reset), .A2(
        InData[5]), .B1(SlicesFromChi[5]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n207) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U21 ( .A1(Reset), .A2(
        InData[6]), .B1(SlicesFromChi[6]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n209) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U20 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n213), .B(
        all_mux_linear_0__MUX_theta_state_inst_n217), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n137) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U19 ( .A1(Reset), .A2(
        InData[9]), .B1(SlicesFromChi[9]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n217) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U18 ( .A1(Reset), .A2(
        InData[8]), .B1(SlicesFromChi[8]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n213) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U17 ( .A1(Reset), .A2(
        InData[7]), .B1(SlicesFromChi[7]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n211) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U16 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n194), .B(
        all_mux_linear_0__MUX_theta_state_inst_n135), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n161) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U15 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n134), .B(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n135) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U14 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n186), .B(
        all_mux_linear_0__MUX_theta_state_inst_n184), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n133) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U13 ( .A1(Reset), .A2(
        InData[20]), .B1(SlicesFromChi[20]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n184) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U12 ( .A1(Reset), .A2(
        InData[21]), .B1(SlicesFromChi[21]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n186) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U11 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n190), .B(
        all_mux_linear_0__MUX_theta_state_inst_n188), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n134) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U10 ( .A1(Reset), .A2(
        InData[22]), .B1(SlicesFromChi[22]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n188) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U9 ( .A1(Reset), .A2(
        InData[23]), .B1(SlicesFromChi[23]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n190) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U8 ( .A1(Reset), .A2(
        InData[24]), .B1(SlicesFromChi[24]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n194) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U7 ( .A1(Reset), .A2(
        InData[0]), .B1(SlicesFromChi[0]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n180) );
  INV_X2 all_mux_linear_0__MUX_theta_state_inst_U6 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n130), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n129) );
  INV_X1 all_mux_linear_0__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n132) );
  INV_X1 all_mux_linear_0__MUX_theta_state_inst_U4 ( .A(Reset), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n131) );
  INV_X1 all_mux_linear_0__MUX_theta_state_inst_U3 ( .A(n2), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n130) );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[9]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[5]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[6]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[7]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[8]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[0]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[1]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[2]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[3]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[4]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[10]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[11]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[12]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[13]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[14]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[15]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[16]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[17]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[18]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[19]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[20]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[21]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[22]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[23]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[24]), .QN() );
  OAI21_X1 all_mux_linear_1__MUX_theta_state_inst_U134 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n334), .A(
        all_mux_linear_1__MUX_theta_state_inst_n333), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_1__MUX_theta_state_inst_U133 ( .A1(n2), .A2(
        SlicesFromChi[34]), .B1(all_mux_linear_1__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_1__MUX_theta_state_inst_n334), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n333) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U132 ( .A1(SlicesFromChi[34]), .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n334) );
  OAI21_X1 all_mux_linear_1__MUX_theta_state_inst_U131 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n331), .A(
        all_mux_linear_1__MUX_theta_state_inst_n330), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_1__MUX_theta_state_inst_U130 ( .A1(n2), .A2(
        SlicesFromChi[33]), .B1(all_mux_linear_1__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_1__MUX_theta_state_inst_n331), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n330) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U129 ( .A1(SlicesFromChi[33]), .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n331) );
  OAI21_X1 all_mux_linear_1__MUX_theta_state_inst_U128 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n329), .A(
        all_mux_linear_1__MUX_theta_state_inst_n328), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_1__MUX_theta_state_inst_U127 ( .A1(n2), .A2(
        SlicesFromChi[32]), .B1(all_mux_linear_1__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_1__MUX_theta_state_inst_n329), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n328) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U126 ( .A1(SlicesFromChi[32]), .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n329) );
  OAI21_X1 all_mux_linear_1__MUX_theta_state_inst_U125 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n327), .A(
        all_mux_linear_1__MUX_theta_state_inst_n326), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_1__MUX_theta_state_inst_U124 ( .A1(n2), .A2(
        SlicesFromChi[31]), .B1(all_mux_linear_1__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_1__MUX_theta_state_inst_n327), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n326) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U123 ( .A1(SlicesFromChi[31]), .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n327) );
  OAI21_X1 all_mux_linear_1__MUX_theta_state_inst_U122 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n325), .A(
        all_mux_linear_1__MUX_theta_state_inst_n324), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_1__MUX_theta_state_inst_U121 ( .A1(n2), .A2(
        SlicesFromChi[30]), .B1(all_mux_linear_1__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_1__MUX_theta_state_inst_n325), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n324) );
  AND2_X1 all_mux_linear_1__MUX_theta_state_inst_U120 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n335), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n332) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U119 ( .A1(SlicesFromChi[30]), .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n325) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U118 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n323), .B(
        all_mux_linear_1__MUX_theta_state_inst_n322), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n335) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U117 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n321), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n319), .A(
        all_mux_linear_1__MUX_theta_state_inst_n318), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[4]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U116 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n321), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n318) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U115 ( .A(SlicesFromChi[29]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n319) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U114 ( .A1(SlicesFromChi[29]), .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n321) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U113 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n317), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n316), .A(
        all_mux_linear_1__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[3]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U112 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n317), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n315) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U111 ( .A(SlicesFromChi[28]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n316) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U110 ( .A1(SlicesFromChi[28]), .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n317) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U109 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n313), .A(
        all_mux_linear_1__MUX_theta_state_inst_n312), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[2]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U108 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n314), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n312) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U107 ( .A1(SlicesFromChi[27]), .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n314) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U106 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n311), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n309), .A(
        all_mux_linear_1__MUX_theta_state_inst_n308), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[24]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n311), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n308) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U104 ( .A(SlicesFromChi[49]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n309) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U103 ( .A1(SlicesFromChi[49]), .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n311) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U102 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n307), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n306), .A(
        all_mux_linear_1__MUX_theta_state_inst_n305), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[23]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U101 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n307), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n305) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U100 ( .A(SlicesFromChi[48]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n306) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U99 ( .A1(SlicesFromChi[48]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n307) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U98 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n304), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n303), .A(
        all_mux_linear_1__MUX_theta_state_inst_n302), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[22]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U97 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n304), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n302) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U96 ( .A1(SlicesFromChi[47]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n304) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n301), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n300), .A(
        all_mux_linear_1__MUX_theta_state_inst_n299), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[21]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n301), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n299) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U93 ( .A(SlicesFromChi[46]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n300) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U92 ( .A1(SlicesFromChi[46]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n301) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n298), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n297), .A(
        all_mux_linear_1__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[20]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n298), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n296) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U89 ( .A(SlicesFromChi[45]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n297) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U88 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n294), .B(
        all_mux_linear_1__MUX_theta_state_inst_n293), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n323) );
  XOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U87 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n292), .B(
        all_mux_linear_1__MUX_theta_state_inst_n291), .Z(
        all_mux_linear_1__MUX_theta_state_inst_n293) );
  OAI211_X1 all_mux_linear_1__MUX_theta_state_inst_U86 ( .C1(SlicesFromChi[29]), .C2(all_mux_linear_1__MUX_theta_state_inst_n290), .A(
        all_mux_linear_1__MUX_theta_state_inst_n232), .B(
        all_mux_linear_1__MUX_theta_state_inst_n289), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n294) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U85 ( .A1(SlicesFromChi[29]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n289) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n313), .B(SlicesFromChi[28]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n290) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U83 ( .A(SlicesFromChi[27]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n313) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U82 ( .A1(SlicesFromChi[45]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n298) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U81 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n288), .A(
        all_mux_linear_1__MUX_theta_state_inst_n287), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[1]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U80 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n291), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n287) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U79 ( .A(SlicesFromChi[26]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n288) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U78 ( .A1(SlicesFromChi[26]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n291) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n286), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n284), .A(
        all_mux_linear_1__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[19]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n286), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n283) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U75 ( .A(SlicesFromChi[44]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n284) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U74 ( .A1(SlicesFromChi[44]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n286) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U73 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n282), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n281), .A(
        all_mux_linear_1__MUX_theta_state_inst_n280), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[18]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U72 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n282), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n280) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U71 ( .A(SlicesFromChi[43]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n281) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U70 ( .A1(SlicesFromChi[43]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n282) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U69 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n279), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n278), .A(
        all_mux_linear_1__MUX_theta_state_inst_n277), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[17]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U68 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n279), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n277) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U67 ( .A1(SlicesFromChi[42]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n279) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n276), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n275), .A(
        all_mux_linear_1__MUX_theta_state_inst_n274), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[16]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n276), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n274) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U64 ( .A(SlicesFromChi[41]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n275) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U63 ( .A1(SlicesFromChi[41]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n276) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U62 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n273), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n272), .A(
        all_mux_linear_1__MUX_theta_state_inst_n271), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[15]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U61 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n273), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n271) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U60 ( .A(SlicesFromChi[40]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n272) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n269), .B(
        all_mux_linear_1__MUX_theta_state_inst_n268), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n322) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n267), .B(
        all_mux_linear_1__MUX_theta_state_inst_n266), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n268) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U57 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n265), .B(
        all_mux_linear_1__MUX_theta_state_inst_n264), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n267) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U56 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n263), .B(
        all_mux_linear_1__MUX_theta_state_inst_n262), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n269) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U55 ( .A1(SlicesFromChi[40]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n273) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n266), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n260), .A(
        all_mux_linear_1__MUX_theta_state_inst_n259), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[14]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n266), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n259) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U52 ( .A(SlicesFromChi[39]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n260) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U51 ( .A1(SlicesFromChi[39]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n266) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U50 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n264), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n258), .A(
        all_mux_linear_1__MUX_theta_state_inst_n257), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[13]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U49 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n264), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n257) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U48 ( .A(SlicesFromChi[38]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n258) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U47 ( .A1(SlicesFromChi[38]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n264) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U46 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n256), .A(
        all_mux_linear_1__MUX_theta_state_inst_n255), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[12]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U45 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n265), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n255) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U44 ( .A(SlicesFromChi[37]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n256) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U43 ( .A1(SlicesFromChi[37]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n265) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U42 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n262), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n254), .A(
        all_mux_linear_1__MUX_theta_state_inst_n253), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[11]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U41 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n262), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n253) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U40 ( .A(SlicesFromChi[36]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n254) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U39 ( .A1(SlicesFromChi[36]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n262) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U38 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n263), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n252), .A(
        all_mux_linear_1__MUX_theta_state_inst_n251), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[10]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U37 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n263), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n251) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U36 ( .A(SlicesFromChi[35]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n252) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n249), .B(
        all_mux_linear_1__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n295) );
  OAI211_X1 all_mux_linear_1__MUX_theta_state_inst_U34 ( .C1(SlicesFromChi[40]), .C2(all_mux_linear_1__MUX_theta_state_inst_n247), .A(
        all_mux_linear_1__MUX_theta_state_inst_n232), .B(
        all_mux_linear_1__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n248) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U33 ( .A1(SlicesFromChi[40]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n246) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U32 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n278), .B(SlicesFromChi[43]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n247) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U31 ( .A(SlicesFromChi[42]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n278) );
  OAI211_X1 all_mux_linear_1__MUX_theta_state_inst_U30 ( .C1(SlicesFromChi[41]), .C2(SlicesFromChi[44]), .A(all_mux_linear_1__MUX_theta_state_inst_n231), .B(
        all_mux_linear_1__MUX_theta_state_inst_n245), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n249) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[44]), 
        .A2(SlicesFromChi[41]), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n245) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U28 ( .A1(SlicesFromChi[35]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n263) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U27 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n292), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n244), .A(
        all_mux_linear_1__MUX_theta_state_inst_n243), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[0]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U26 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n292), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n243) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U25 ( .A(SlicesFromChi[25]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n244) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n242), .B(
        all_mux_linear_1__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n250) );
  AOI211_X1 all_mux_linear_1__MUX_theta_state_inst_U23 ( .C1(SlicesFromChi[31]), .C2(SlicesFromChi[32]), .A(Reset), .B(
        all_mux_linear_1__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n241) );
  NOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U22 ( .A1(SlicesFromChi[31]), 
        .A2(SlicesFromChi[32]), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n240) );
  OAI211_X1 all_mux_linear_1__MUX_theta_state_inst_U21 ( .C1(SlicesFromChi[30]), .C2(all_mux_linear_1__MUX_theta_state_inst_n239), .A(
        all_mux_linear_1__MUX_theta_state_inst_n231), .B(
        all_mux_linear_1__MUX_theta_state_inst_n238), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n242) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U20 ( .A1(SlicesFromChi[30]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n239), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n238) );
  XOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U19 ( .A(SlicesFromChi[34]), 
        .B(SlicesFromChi[33]), .Z(all_mux_linear_1__MUX_theta_state_inst_n239)
         );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U18 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n237), .B(
        all_mux_linear_1__MUX_theta_state_inst_n236), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n270) );
  AOI211_X1 all_mux_linear_1__MUX_theta_state_inst_U17 ( .C1(SlicesFromChi[46]), .C2(SlicesFromChi[49]), .A(Reset), .B(
        all_mux_linear_1__MUX_theta_state_inst_n235), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n236) );
  NOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U16 ( .A1(SlicesFromChi[46]), 
        .A2(SlicesFromChi[49]), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n235) );
  OAI211_X1 all_mux_linear_1__MUX_theta_state_inst_U15 ( .C1(SlicesFromChi[45]), .C2(all_mux_linear_1__MUX_theta_state_inst_n234), .A(
        all_mux_linear_1__MUX_theta_state_inst_n231), .B(
        all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n237) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U14 ( .A1(SlicesFromChi[45]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n233) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U13 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n303), .B(SlicesFromChi[48]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n234) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U12 ( .A(SlicesFromChi[47]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n303) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U11 ( .A1(SlicesFromChi[25]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n292) );
  XOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U10 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n270), .B(
        all_mux_linear_1__MUX_theta_state_inst_n250), .Z(
        all_mux_linear_1__MUX_theta_state_inst_n320) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U9 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n270), .B(
        all_mux_linear_1__MUX_theta_state_inst_n322), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n285) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U8 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n323), .B(
        all_mux_linear_1__MUX_theta_state_inst_n295), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n310) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U7 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n250), .B(
        all_mux_linear_1__MUX_theta_state_inst_n295), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n261) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U6 ( .A(Reset), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n231) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U4 ( .A(n2), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n230) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U3 ( .A(n2), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n229) );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[25]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[26]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[27]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[28]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[29]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[30]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[31]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[32]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[33]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[34]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[35]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[36]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[37]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[38]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[39]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[40]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[41]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[42]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[43]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[44]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[45]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[46]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[47]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[48]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[49]), .QN() );
  OAI21_X1 all_mux_linear_2__MUX_theta_state_inst_U134 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n334), .A(
        all_mux_linear_2__MUX_theta_state_inst_n333), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_2__MUX_theta_state_inst_U133 ( .A1(n2), .A2(
        SlicesFromChi[59]), .B1(all_mux_linear_2__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_2__MUX_theta_state_inst_n334), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n333) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U132 ( .A1(SlicesFromChi[59]), .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n334) );
  OAI21_X1 all_mux_linear_2__MUX_theta_state_inst_U131 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n331), .A(
        all_mux_linear_2__MUX_theta_state_inst_n330), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_2__MUX_theta_state_inst_U130 ( .A1(n2), .A2(
        SlicesFromChi[58]), .B1(all_mux_linear_2__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_2__MUX_theta_state_inst_n331), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n330) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U129 ( .A1(SlicesFromChi[58]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n331) );
  OAI21_X1 all_mux_linear_2__MUX_theta_state_inst_U128 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n329), .A(
        all_mux_linear_2__MUX_theta_state_inst_n328), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_2__MUX_theta_state_inst_U127 ( .A1(n2), .A2(
        SlicesFromChi[57]), .B1(all_mux_linear_2__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_2__MUX_theta_state_inst_n329), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n328) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U126 ( .A1(SlicesFromChi[57]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n329) );
  OAI21_X1 all_mux_linear_2__MUX_theta_state_inst_U125 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n327), .A(
        all_mux_linear_2__MUX_theta_state_inst_n326), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_2__MUX_theta_state_inst_U124 ( .A1(n2), .A2(
        SlicesFromChi[56]), .B1(all_mux_linear_2__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_2__MUX_theta_state_inst_n327), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n326) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U123 ( .A1(SlicesFromChi[56]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n327) );
  OAI21_X1 all_mux_linear_2__MUX_theta_state_inst_U122 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n325), .A(
        all_mux_linear_2__MUX_theta_state_inst_n324), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_2__MUX_theta_state_inst_U121 ( .A1(n2), .A2(
        SlicesFromChi[55]), .B1(all_mux_linear_2__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_2__MUX_theta_state_inst_n325), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n324) );
  AND2_X1 all_mux_linear_2__MUX_theta_state_inst_U120 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n335), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n332) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U119 ( .A1(SlicesFromChi[55]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n325) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U118 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n323), .B(
        all_mux_linear_2__MUX_theta_state_inst_n322), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n335) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U117 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n321), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n319), .A(
        all_mux_linear_2__MUX_theta_state_inst_n318), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[4]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U116 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n321), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n318) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U115 ( .A(SlicesFromChi[54]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n319) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U114 ( .A1(SlicesFromChi[54]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n321) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U113 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n317), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n316), .A(
        all_mux_linear_2__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[3]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U112 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n317), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n315) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U111 ( .A(SlicesFromChi[53]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n316) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U110 ( .A1(SlicesFromChi[53]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n317) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U109 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n313), .A(
        all_mux_linear_2__MUX_theta_state_inst_n312), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[2]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U108 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n314), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n312) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U107 ( .A1(SlicesFromChi[52]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n314) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U106 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n311), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n309), .A(
        all_mux_linear_2__MUX_theta_state_inst_n308), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[24]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n311), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n308) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U104 ( .A(SlicesFromChi[74]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n309) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U103 ( .A1(SlicesFromChi[74]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n311) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U102 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n307), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n306), .A(
        all_mux_linear_2__MUX_theta_state_inst_n305), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[23]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U101 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n307), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n305) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U100 ( .A(SlicesFromChi[73]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n306) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U99 ( .A1(SlicesFromChi[73]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n307) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U98 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n304), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n303), .A(
        all_mux_linear_2__MUX_theta_state_inst_n302), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[22]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U97 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n304), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n302) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U96 ( .A1(SlicesFromChi[72]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n304) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n301), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n300), .A(
        all_mux_linear_2__MUX_theta_state_inst_n299), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[21]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n301), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n299) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U93 ( .A(SlicesFromChi[71]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n300) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U92 ( .A1(SlicesFromChi[71]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n301) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n298), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n297), .A(
        all_mux_linear_2__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[20]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n298), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n296) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U89 ( .A(SlicesFromChi[70]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n297) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U88 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n294), .B(
        all_mux_linear_2__MUX_theta_state_inst_n293), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n323) );
  XOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U87 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n292), .B(
        all_mux_linear_2__MUX_theta_state_inst_n291), .Z(
        all_mux_linear_2__MUX_theta_state_inst_n293) );
  OAI211_X1 all_mux_linear_2__MUX_theta_state_inst_U86 ( .C1(SlicesFromChi[54]), .C2(all_mux_linear_2__MUX_theta_state_inst_n290), .A(
        all_mux_linear_2__MUX_theta_state_inst_n232), .B(
        all_mux_linear_2__MUX_theta_state_inst_n289), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n294) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U85 ( .A1(SlicesFromChi[54]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n289) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n313), .B(SlicesFromChi[53]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n290) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U83 ( .A(SlicesFromChi[52]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n313) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U82 ( .A1(SlicesFromChi[70]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n298) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U81 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n288), .A(
        all_mux_linear_2__MUX_theta_state_inst_n287), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[1]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U80 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n291), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n287) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U79 ( .A(SlicesFromChi[51]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n288) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U78 ( .A1(SlicesFromChi[51]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n291) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n286), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n284), .A(
        all_mux_linear_2__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[19]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n286), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n283) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U75 ( .A(SlicesFromChi[69]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n284) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U74 ( .A1(SlicesFromChi[69]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n286) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U73 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n282), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n281), .A(
        all_mux_linear_2__MUX_theta_state_inst_n280), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[18]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U72 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n282), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n280) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U71 ( .A(SlicesFromChi[68]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n281) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U70 ( .A1(SlicesFromChi[68]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n282) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U69 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n279), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n278), .A(
        all_mux_linear_2__MUX_theta_state_inst_n277), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[17]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U68 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n279), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n277) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U67 ( .A1(SlicesFromChi[67]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n279) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n276), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n275), .A(
        all_mux_linear_2__MUX_theta_state_inst_n274), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[16]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n276), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n274) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U64 ( .A(SlicesFromChi[66]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n275) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U63 ( .A1(SlicesFromChi[66]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n276) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U62 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n273), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n272), .A(
        all_mux_linear_2__MUX_theta_state_inst_n271), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[15]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U61 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n273), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n271) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U60 ( .A(SlicesFromChi[65]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n272) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n269), .B(
        all_mux_linear_2__MUX_theta_state_inst_n268), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n322) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n267), .B(
        all_mux_linear_2__MUX_theta_state_inst_n266), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n268) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U57 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n265), .B(
        all_mux_linear_2__MUX_theta_state_inst_n264), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n267) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U56 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n263), .B(
        all_mux_linear_2__MUX_theta_state_inst_n262), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n269) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U55 ( .A1(SlicesFromChi[65]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n273) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n266), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n260), .A(
        all_mux_linear_2__MUX_theta_state_inst_n259), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[14]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n266), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n259) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U52 ( .A(SlicesFromChi[64]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n260) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U51 ( .A1(SlicesFromChi[64]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n266) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U50 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n264), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n258), .A(
        all_mux_linear_2__MUX_theta_state_inst_n257), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[13]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U49 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n264), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n257) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U48 ( .A(SlicesFromChi[63]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n258) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U47 ( .A1(SlicesFromChi[63]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n264) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U46 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n256), .A(
        all_mux_linear_2__MUX_theta_state_inst_n255), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[12]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U45 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n265), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n255) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U44 ( .A(SlicesFromChi[62]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n256) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U43 ( .A1(SlicesFromChi[62]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n265) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U42 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n262), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n254), .A(
        all_mux_linear_2__MUX_theta_state_inst_n253), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[11]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U41 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n262), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n253) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U40 ( .A(SlicesFromChi[61]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n254) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U39 ( .A1(SlicesFromChi[61]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n262) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U38 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n263), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n252), .A(
        all_mux_linear_2__MUX_theta_state_inst_n251), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[10]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U37 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n263), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n251) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U36 ( .A(SlicesFromChi[60]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n252) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n249), .B(
        all_mux_linear_2__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n295) );
  OAI211_X1 all_mux_linear_2__MUX_theta_state_inst_U34 ( .C1(SlicesFromChi[65]), .C2(all_mux_linear_2__MUX_theta_state_inst_n247), .A(
        all_mux_linear_2__MUX_theta_state_inst_n232), .B(
        all_mux_linear_2__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n248) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U33 ( .A1(SlicesFromChi[65]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n246) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U32 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n278), .B(SlicesFromChi[68]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n247) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U31 ( .A(SlicesFromChi[67]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n278) );
  OAI211_X1 all_mux_linear_2__MUX_theta_state_inst_U30 ( .C1(SlicesFromChi[66]), .C2(SlicesFromChi[69]), .A(all_mux_linear_2__MUX_theta_state_inst_n231), .B(
        all_mux_linear_2__MUX_theta_state_inst_n245), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n249) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[69]), 
        .A2(SlicesFromChi[66]), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n245) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U28 ( .A1(SlicesFromChi[60]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n263) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U27 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n292), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n244), .A(
        all_mux_linear_2__MUX_theta_state_inst_n243), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[0]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U26 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n292), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n243) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U25 ( .A(SlicesFromChi[50]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n244) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n242), .B(
        all_mux_linear_2__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n250) );
  AOI211_X1 all_mux_linear_2__MUX_theta_state_inst_U23 ( .C1(SlicesFromChi[56]), .C2(SlicesFromChi[57]), .A(Reset), .B(
        all_mux_linear_2__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n241) );
  NOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U22 ( .A1(SlicesFromChi[56]), 
        .A2(SlicesFromChi[57]), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n240) );
  OAI211_X1 all_mux_linear_2__MUX_theta_state_inst_U21 ( .C1(SlicesFromChi[55]), .C2(all_mux_linear_2__MUX_theta_state_inst_n239), .A(
        all_mux_linear_2__MUX_theta_state_inst_n231), .B(
        all_mux_linear_2__MUX_theta_state_inst_n238), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n242) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U20 ( .A1(SlicesFromChi[55]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n239), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n238) );
  XOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U19 ( .A(SlicesFromChi[59]), 
        .B(SlicesFromChi[58]), .Z(all_mux_linear_2__MUX_theta_state_inst_n239)
         );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U18 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n237), .B(
        all_mux_linear_2__MUX_theta_state_inst_n236), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n270) );
  AOI211_X1 all_mux_linear_2__MUX_theta_state_inst_U17 ( .C1(SlicesFromChi[71]), .C2(SlicesFromChi[74]), .A(Reset), .B(
        all_mux_linear_2__MUX_theta_state_inst_n235), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n236) );
  NOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U16 ( .A1(SlicesFromChi[71]), 
        .A2(SlicesFromChi[74]), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n235) );
  OAI211_X1 all_mux_linear_2__MUX_theta_state_inst_U15 ( .C1(SlicesFromChi[70]), .C2(all_mux_linear_2__MUX_theta_state_inst_n234), .A(
        all_mux_linear_2__MUX_theta_state_inst_n231), .B(
        all_mux_linear_2__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n237) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U14 ( .A1(SlicesFromChi[70]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n233) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U13 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n303), .B(SlicesFromChi[73]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n234) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U12 ( .A(SlicesFromChi[72]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n303) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U11 ( .A1(SlicesFromChi[50]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n292) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U10 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n250), .B(
        all_mux_linear_2__MUX_theta_state_inst_n295), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n261) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U9 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n323), .B(
        all_mux_linear_2__MUX_theta_state_inst_n295), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n310) );
  XOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U8 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n270), .B(
        all_mux_linear_2__MUX_theta_state_inst_n250), .Z(
        all_mux_linear_2__MUX_theta_state_inst_n320) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U7 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n270), .B(
        all_mux_linear_2__MUX_theta_state_inst_n322), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n285) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U6 ( .A(Reset), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n231) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U4 ( .A(n2), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n230) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U3 ( .A(n2), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n229) );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[50]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[51]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[52]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[53]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[54]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[55]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[56]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[57]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[58]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[59]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[60]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[61]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[62]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[63]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[64]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[65]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[66]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[67]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[68]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[69]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[70]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[71]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[72]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[73]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[74]), .QN() );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U116 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n318), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n317), .A(
        all_mux_linear_3__MUX_theta_state_inst_n316), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U115 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[84]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n318), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n316) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U114 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n317), .A(
        all_mux_linear_3__MUX_theta_state_inst_n313), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U113 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[83]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n313) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U112 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n312), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n317), .A(
        all_mux_linear_3__MUX_theta_state_inst_n311), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U111 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[82]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n312), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n311) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U110 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n310), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n317), .A(
        all_mux_linear_3__MUX_theta_state_inst_n309), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U109 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[81]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n310), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n309) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U108 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n308), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n317), .A(
        all_mux_linear_3__MUX_theta_state_inst_n307), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U107 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[80]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n308), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n307) );
  NOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U106 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n306), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n315) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n306), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n317) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U104 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n305), .B(
        all_mux_linear_3__MUX_theta_state_inst_n304), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n306) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U103 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n303), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n302), .A(
        all_mux_linear_3__MUX_theta_state_inst_n301), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[4]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U102 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[79]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n303), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n301) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U101 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n299), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n302), .A(
        all_mux_linear_3__MUX_theta_state_inst_n298), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[3]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U100 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[78]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n299), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n298) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U99 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n297), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n302), .A(
        all_mux_linear_3__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[2]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U98 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[77]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n297), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n296) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U97 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n295), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n294), .A(
        all_mux_linear_3__MUX_theta_state_inst_n293), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[24]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U96 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[99]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n295), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n293) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n294), .A(
        all_mux_linear_3__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[23]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[98]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n290) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U93 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n289), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n294), .A(
        all_mux_linear_3__MUX_theta_state_inst_n288), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[22]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U92 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[97]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n289), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n288) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n287), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n294), .A(
        all_mux_linear_3__MUX_theta_state_inst_n286), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[21]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[96]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n287), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n286) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U89 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n285), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n294), .A(
        all_mux_linear_3__MUX_theta_state_inst_n284), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[20]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U88 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[95]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n285), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n284) );
  NOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U87 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n292) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U86 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n294) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U85 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n282), .B(
        all_mux_linear_3__MUX_theta_state_inst_n304), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n283) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n281), .B(
        all_mux_linear_3__MUX_theta_state_inst_n280), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n304) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U83 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n279), .B(
        all_mux_linear_3__MUX_theta_state_inst_n278), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n280) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U82 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n277), .B(
        all_mux_linear_3__MUX_theta_state_inst_n303), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n278) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U81 ( .A1(Reset), .A2(
        InData[29]), .B1(SlicesFromChi[79]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n303) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U80 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n299), .B(
        all_mux_linear_3__MUX_theta_state_inst_n297), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n279) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U79 ( .A1(Reset), .A2(
        InData[27]), .B1(SlicesFromChi[77]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n297) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U78 ( .A1(Reset), .A2(
        InData[28]), .B1(SlicesFromChi[78]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n299) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n277), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n302), .A(
        all_mux_linear_3__MUX_theta_state_inst_n276), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[1]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[76]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n277), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n276) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U75 ( .A1(Reset), .A2(
        InData[26]), .B1(SlicesFromChi[76]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n277) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U74 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n275), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n274), .A(
        all_mux_linear_3__MUX_theta_state_inst_n273), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[19]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U73 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[94]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n275), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n273) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U72 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n271), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n274), .A(
        all_mux_linear_3__MUX_theta_state_inst_n270), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[18]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U71 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[93]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n271), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n270) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U70 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n269), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n274), .A(
        all_mux_linear_3__MUX_theta_state_inst_n268), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[17]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U69 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[92]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n269), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n268) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U68 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n267), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n274), .A(
        all_mux_linear_3__MUX_theta_state_inst_n266), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[16]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U67 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[91]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n267), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n266) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n274), .A(
        all_mux_linear_3__MUX_theta_state_inst_n264), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[15]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[90]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n264) );
  NOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U64 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n263), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n272) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U63 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n263), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n274) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U62 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n262), .B(
        all_mux_linear_3__MUX_theta_state_inst_n305), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n263) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U61 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n261), .B(
        all_mux_linear_3__MUX_theta_state_inst_n260), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n305) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U60 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n259), .B(
        all_mux_linear_3__MUX_theta_state_inst_n258), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n260) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n257), .B(
        all_mux_linear_3__MUX_theta_state_inst_n256), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n258) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n255), .B(
        all_mux_linear_3__MUX_theta_state_inst_n254), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n259) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U57 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n255), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n253), .A(
        all_mux_linear_3__MUX_theta_state_inst_n252), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[14]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U56 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[89]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n255), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n252) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U55 ( .A1(Reset), .A2(
        InData[39]), .B1(SlicesFromChi[89]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n255) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n254), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n253), .A(
        all_mux_linear_3__MUX_theta_state_inst_n250), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[13]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[88]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n254), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n250) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U52 ( .A1(Reset), .A2(
        InData[38]), .B1(SlicesFromChi[88]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n254) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U51 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n256), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n253), .A(
        all_mux_linear_3__MUX_theta_state_inst_n249), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[12]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U50 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[87]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n256), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n249) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U49 ( .A1(Reset), .A2(
        InData[37]), .B1(SlicesFromChi[87]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n256) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U48 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n257), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n253), .A(
        all_mux_linear_3__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[11]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U47 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[86]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n257), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n248) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U46 ( .A1(Reset), .A2(
        InData[36]), .B1(SlicesFromChi[86]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n257) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U45 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n261), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n253), .A(
        all_mux_linear_3__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[10]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U44 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(SlicesFromChi[85]), 
        .B1(all_mux_linear_3__MUX_theta_state_inst_n261), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n251), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n247) );
  NOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U43 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n251) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U42 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n253) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U41 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n245), .B(
        all_mux_linear_3__MUX_theta_state_inst_n282), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n246) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U40 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n275), .B(
        all_mux_linear_3__MUX_theta_state_inst_n244), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n282) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U39 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n243), .B(
        all_mux_linear_3__MUX_theta_state_inst_n242), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n244) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U38 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n267), .B(
        all_mux_linear_3__MUX_theta_state_inst_n265), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n242) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U37 ( .A1(Reset), .A2(
        InData[40]), .B1(SlicesFromChi[90]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n265) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U36 ( .A1(Reset), .A2(
        InData[41]), .B1(SlicesFromChi[91]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n267) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n271), .B(
        all_mux_linear_3__MUX_theta_state_inst_n269), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n243) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U34 ( .A1(Reset), .A2(
        InData[42]), .B1(SlicesFromChi[92]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n269) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U33 ( .A1(Reset), .A2(
        InData[43]), .B1(SlicesFromChi[93]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n271) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U32 ( .A1(Reset), .A2(
        InData[44]), .B1(SlicesFromChi[94]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n275) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U31 ( .A1(Reset), .A2(
        InData[35]), .B1(SlicesFromChi[85]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n261) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U30 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n281), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n302), .A(
        all_mux_linear_3__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[0]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[75]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n230), .B1(
        all_mux_linear_3__MUX_theta_state_inst_n281), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n300), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n241) );
  NOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U28 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n300) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U27 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n302) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U26 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n262), .B(
        all_mux_linear_3__MUX_theta_state_inst_n245), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n240) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U25 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n312), .B(
        all_mux_linear_3__MUX_theta_state_inst_n239), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n245) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n238), .B(
        all_mux_linear_3__MUX_theta_state_inst_n237), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n239) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U23 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n310), .B(
        all_mux_linear_3__MUX_theta_state_inst_n308), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n237) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U22 ( .A1(Reset), .A2(
        InData[30]), .B1(SlicesFromChi[80]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n308) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U21 ( .A1(Reset), .A2(
        InData[31]), .B1(SlicesFromChi[81]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n310) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U20 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n314), .B(
        all_mux_linear_3__MUX_theta_state_inst_n318), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n238) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U19 ( .A1(Reset), .A2(
        InData[34]), .B1(SlicesFromChi[84]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n318) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U18 ( .A1(Reset), .A2(
        InData[33]), .B1(SlicesFromChi[83]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n314) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U17 ( .A1(Reset), .A2(
        InData[32]), .B1(SlicesFromChi[82]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n312) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U16 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n295), .B(
        all_mux_linear_3__MUX_theta_state_inst_n236), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n262) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U15 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n235), .B(
        all_mux_linear_3__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n236) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U14 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n287), .B(
        all_mux_linear_3__MUX_theta_state_inst_n285), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n234) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U13 ( .A1(Reset), .A2(
        InData[45]), .B1(SlicesFromChi[95]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n285) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U12 ( .A1(Reset), .A2(
        InData[46]), .B1(SlicesFromChi[96]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n287) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U11 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n291), .B(
        all_mux_linear_3__MUX_theta_state_inst_n289), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n235) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U10 ( .A1(Reset), .A2(
        InData[47]), .B1(SlicesFromChi[97]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n289) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U9 ( .A1(Reset), .A2(
        InData[48]), .B1(SlicesFromChi[98]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n291) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U8 ( .A1(Reset), .A2(
        InData[49]), .B1(SlicesFromChi[99]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n295) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U7 ( .A1(Reset), .A2(
        InData[25]), .B1(SlicesFromChi[75]), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n281) );
  INV_X2 all_mux_linear_3__MUX_theta_state_inst_U6 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n230) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n233) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U4 ( .A(Reset), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U3 ( .A(n2), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n231) );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[75]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[76]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[77]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[78]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[79]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[80]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[81]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[82]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[83]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[84]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[85]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[86]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[87]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[88]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[89]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[90]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[91]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[92]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[93]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[94]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[95]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[96]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[97]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[98]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[99]), .QN() );
  XOR2_X1 COMPRESSION_BITS_0__BIT_SHARES_0__Copression_U1 ( .A(StateOut[0]), 
        .B(StateOut[25]), .Z(OutData[0]) );
  XOR2_X1 COMPRESSION_BITS_0__BIT_SHARES_1__Copression_U1 ( .A(StateOut[50]), 
        .B(StateOut[75]), .Z(OutData[25]) );
  XOR2_X1 COMPRESSION_BITS_1__BIT_SHARES_0__Copression_U1 ( .A(StateOut[1]), 
        .B(StateOut[26]), .Z(OutData[1]) );
  XOR2_X1 COMPRESSION_BITS_1__BIT_SHARES_1__Copression_U1 ( .A(StateOut[51]), 
        .B(StateOut[76]), .Z(OutData[26]) );
  XOR2_X1 COMPRESSION_BITS_2__BIT_SHARES_0__Copression_U1 ( .A(StateOut[2]), 
        .B(StateOut[27]), .Z(OutData[2]) );
  XOR2_X1 COMPRESSION_BITS_2__BIT_SHARES_1__Copression_U1 ( .A(StateOut[52]), 
        .B(StateOut[77]), .Z(OutData[27]) );
  XOR2_X1 COMPRESSION_BITS_3__BIT_SHARES_0__Copression_U1 ( .A(StateOut[3]), 
        .B(StateOut[28]), .Z(OutData[3]) );
  XOR2_X1 COMPRESSION_BITS_3__BIT_SHARES_1__Copression_U1 ( .A(StateOut[53]), 
        .B(StateOut[78]), .Z(OutData[28]) );
  XOR2_X1 COMPRESSION_BITS_4__BIT_SHARES_0__Copression_U1 ( .A(StateOut[4]), 
        .B(StateOut[29]), .Z(OutData[4]) );
  XOR2_X1 COMPRESSION_BITS_4__BIT_SHARES_1__Copression_U1 ( .A(StateOut[54]), 
        .B(StateOut[79]), .Z(OutData[29]) );
  XOR2_X1 COMPRESSION_BITS_5__BIT_SHARES_0__Copression_U1 ( .A(StateOut[5]), 
        .B(StateOut[30]), .Z(OutData[5]) );
  XOR2_X1 COMPRESSION_BITS_5__BIT_SHARES_1__Copression_U1 ( .A(StateOut[55]), 
        .B(StateOut[80]), .Z(OutData[30]) );
  XOR2_X1 COMPRESSION_BITS_6__BIT_SHARES_0__Copression_U1 ( .A(StateOut[6]), 
        .B(StateOut[31]), .Z(OutData[6]) );
  XOR2_X1 COMPRESSION_BITS_6__BIT_SHARES_1__Copression_U1 ( .A(StateOut[56]), 
        .B(StateOut[81]), .Z(OutData[31]) );
  XOR2_X1 COMPRESSION_BITS_7__BIT_SHARES_0__Copression_U1 ( .A(StateOut[7]), 
        .B(StateOut[32]), .Z(OutData[7]) );
  XOR2_X1 COMPRESSION_BITS_7__BIT_SHARES_1__Copression_U1 ( .A(StateOut[57]), 
        .B(StateOut[82]), .Z(OutData[32]) );
  XOR2_X1 COMPRESSION_BITS_8__BIT_SHARES_0__Copression_U1 ( .A(StateOut[8]), 
        .B(StateOut[33]), .Z(OutData[8]) );
  XOR2_X1 COMPRESSION_BITS_8__BIT_SHARES_1__Copression_U1 ( .A(StateOut[58]), 
        .B(StateOut[83]), .Z(OutData[33]) );
  XOR2_X1 COMPRESSION_BITS_9__BIT_SHARES_0__Copression_U1 ( .A(StateOut[9]), 
        .B(StateOut[34]), .Z(OutData[9]) );
  XOR2_X1 COMPRESSION_BITS_9__BIT_SHARES_1__Copression_U1 ( .A(StateOut[59]), 
        .B(StateOut[84]), .Z(OutData[34]) );
  XOR2_X1 COMPRESSION_BITS_10__BIT_SHARES_0__Copression_U1 ( .A(StateOut[10]), 
        .B(StateOut[35]), .Z(OutData[10]) );
  XOR2_X1 COMPRESSION_BITS_10__BIT_SHARES_1__Copression_U1 ( .A(StateOut[60]), 
        .B(StateOut[85]), .Z(OutData[35]) );
  XOR2_X1 COMPRESSION_BITS_11__BIT_SHARES_0__Copression_U1 ( .A(StateOut[11]), 
        .B(StateOut[36]), .Z(OutData[11]) );
  XOR2_X1 COMPRESSION_BITS_11__BIT_SHARES_1__Copression_U1 ( .A(StateOut[61]), 
        .B(StateOut[86]), .Z(OutData[36]) );
  XOR2_X1 COMPRESSION_BITS_12__BIT_SHARES_0__Copression_U1 ( .A(StateOut[12]), 
        .B(StateOut[37]), .Z(OutData[12]) );
  XOR2_X1 COMPRESSION_BITS_12__BIT_SHARES_1__Copression_U1 ( .A(StateOut[62]), 
        .B(StateOut[87]), .Z(OutData[37]) );
  XOR2_X1 COMPRESSION_BITS_13__BIT_SHARES_0__Copression_U1 ( .A(StateOut[13]), 
        .B(StateOut[38]), .Z(OutData[13]) );
  XOR2_X1 COMPRESSION_BITS_13__BIT_SHARES_1__Copression_U1 ( .A(StateOut[63]), 
        .B(StateOut[88]), .Z(OutData[38]) );
  XOR2_X1 COMPRESSION_BITS_14__BIT_SHARES_0__Copression_U1 ( .A(StateOut[14]), 
        .B(StateOut[39]), .Z(OutData[14]) );
  XOR2_X1 COMPRESSION_BITS_14__BIT_SHARES_1__Copression_U1 ( .A(StateOut[64]), 
        .B(StateOut[89]), .Z(OutData[39]) );
  XOR2_X1 COMPRESSION_BITS_15__BIT_SHARES_0__Copression_U1 ( .A(StateOut[15]), 
        .B(StateOut[65]), .Z(OutData[15]) );
  XOR2_X1 COMPRESSION_BITS_15__BIT_SHARES_1__Copression_U1 ( .A(StateOut[40]), 
        .B(StateOut[90]), .Z(OutData[40]) );
  XOR2_X1 COMPRESSION_BITS_16__BIT_SHARES_0__Copression_U1 ( .A(StateOut[16]), 
        .B(StateOut[66]), .Z(OutData[16]) );
  XOR2_X1 COMPRESSION_BITS_16__BIT_SHARES_1__Copression_U1 ( .A(StateOut[41]), 
        .B(StateOut[91]), .Z(OutData[41]) );
  XOR2_X1 COMPRESSION_BITS_17__BIT_SHARES_0__Copression_U1 ( .A(StateOut[17]), 
        .B(StateOut[67]), .Z(OutData[17]) );
  XOR2_X1 COMPRESSION_BITS_17__BIT_SHARES_1__Copression_U1 ( .A(StateOut[42]), 
        .B(StateOut[92]), .Z(OutData[42]) );
  XOR2_X1 COMPRESSION_BITS_18__BIT_SHARES_0__Copression_U1 ( .A(StateOut[18]), 
        .B(StateOut[68]), .Z(OutData[18]) );
  XOR2_X1 COMPRESSION_BITS_18__BIT_SHARES_1__Copression_U1 ( .A(StateOut[43]), 
        .B(StateOut[93]), .Z(OutData[43]) );
  XOR2_X1 COMPRESSION_BITS_19__BIT_SHARES_0__Copression_U1 ( .A(StateOut[19]), 
        .B(StateOut[69]), .Z(OutData[19]) );
  XOR2_X1 COMPRESSION_BITS_19__BIT_SHARES_1__Copression_U1 ( .A(StateOut[44]), 
        .B(StateOut[94]), .Z(OutData[44]) );
  XOR2_X1 COMPRESSION_BITS_20__BIT_SHARES_0__Copression_U1 ( .A(StateOut[20]), 
        .B(StateOut[45]), .Z(OutData[20]) );
  XOR2_X1 COMPRESSION_BITS_20__BIT_SHARES_1__Copression_U1 ( .A(StateOut[70]), 
        .B(StateOut[95]), .Z(OutData[45]) );
  XOR2_X1 COMPRESSION_BITS_21__BIT_SHARES_0__Copression_U1 ( .A(StateOut[21]), 
        .B(StateOut[46]), .Z(OutData[21]) );
  XOR2_X1 COMPRESSION_BITS_21__BIT_SHARES_1__Copression_U1 ( .A(StateOut[71]), 
        .B(StateOut[96]), .Z(OutData[46]) );
  XOR2_X1 COMPRESSION_BITS_22__BIT_SHARES_0__Copression_U1 ( .A(StateOut[22]), 
        .B(StateOut[47]), .Z(OutData[22]) );
  XOR2_X1 COMPRESSION_BITS_22__BIT_SHARES_1__Copression_U1 ( .A(StateOut[72]), 
        .B(StateOut[97]), .Z(OutData[47]) );
  XOR2_X1 COMPRESSION_BITS_23__BIT_SHARES_0__Copression_U1 ( .A(StateOut[23]), 
        .B(StateOut[48]), .Z(OutData[23]) );
  XOR2_X1 COMPRESSION_BITS_23__BIT_SHARES_1__Copression_U1 ( .A(StateOut[73]), 
        .B(StateOut[98]), .Z(OutData[48]) );
  XOR2_X1 COMPRESSION_BITS_24__BIT_SHARES_0__Copression_U1 ( .A(StateOut[24]), 
        .B(StateOut[49]), .Z(OutData[24]) );
  XOR2_X1 COMPRESSION_BITS_24__BIT_SHARES_1__Copression_U1 ( .A(StateOut[74]), 
        .B(StateOut[99]), .Z(OutData[49]) );
  XOR2_X1 CHI_U1 ( .A(CHI_ChiOut_0_), .B(IotaRC_0_), .Z(SlicesFromChi[0]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(OutData[0]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n3), .ZN(CHI_ChiOut_0_) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[12]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n2), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n3) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(OutData[6]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n2) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A(OutData[6]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[5]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A1(OutData[18]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(OutData[12]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U3 ( 
        .A(OutData[12]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7), .ZN(SlicesFromChi[10]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A1(OutData[24]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A(OutData[18]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A(OutData[18]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[15]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A1(OutData[0]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(OutData[24]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U3 ( 
        .A(OutData[24]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7), .ZN(SlicesFromChi[20]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U2 ( 
        .A1(OutData[6]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A(OutData[0]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U3 ( 
        .A(FreshRand[0]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5), .ZN(SlicesFromChi[25]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A1(OutData[37]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A(OutData[6]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[1]), .ZN(SlicesFromChi[30]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[37]), .A2(OutData[18]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7), .ZN(SlicesFromChi[35]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U3 ( 
        .A1(OutData[49]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(OutData[18]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A(FreshRand[2]), .B(OutData[37]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[25]), .A2(OutData[49]), .ZN(SlicesFromChi[40]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[45]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[25]), .A2(OutData[6]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(FreshRand[4]), .B(OutData[49]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[50]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[31]), .A2(OutData[12]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[0]), .B(OutData[25]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[55]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[43]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[12]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[1]), .B(OutData[31]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[2]), .ZN(SlicesFromChi[60]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[43]), .A2(OutData[24]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[65]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[25]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[24]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[3]), .B(OutData[43]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[31]), .A2(OutData[25]), .ZN(SlicesFromChi[70]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[37]), .A2(OutData[31]), .ZN(SlicesFromChi[75]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[43]), .A2(OutData[37]), .ZN(SlicesFromChi[80]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[49]), .A2(OutData[43]), .ZN(SlicesFromChi[85]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[3]), .ZN(SlicesFromChi[90]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[49]), .A2(OutData[0]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(FreshRand[4]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[95]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[31]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(OutData[0]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(OutData[15]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7), .ZN(SlicesFromChi[1]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[2]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(OutData[21]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A(OutData[21]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[6]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A1(OutData[8]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(OutData[2]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U3 ( 
        .A(OutData[2]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7), .ZN(SlicesFromChi[11]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A1(OutData[14]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A(OutData[8]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A(OutData[8]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[16]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A1(OutData[15]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(OutData[14]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U3 ( 
        .A(OutData[14]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7), .ZN(SlicesFromChi[21]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U2 ( 
        .A1(OutData[21]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A(OutData[15]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U3 ( 
        .A(FreshRand[5]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5), .ZN(SlicesFromChi[26]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A1(OutData[27]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A(OutData[21]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[6]), .ZN(SlicesFromChi[31]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[27]), .A2(OutData[8]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7), .ZN(SlicesFromChi[36]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U3 ( 
        .A1(OutData[39]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(OutData[8]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A(FreshRand[7]), .B(OutData[27]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[40]), .A2(OutData[39]), .ZN(SlicesFromChi[41]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[46]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[40]), .A2(OutData[21]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(FreshRand[9]), .B(OutData[39]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[51]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[46]), .A2(OutData[2]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[5]), .B(OutData[40]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[56]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[33]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[2]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[6]), .B(OutData[46]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[7]), .ZN(SlicesFromChi[61]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[33]), .A2(OutData[14]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[66]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[40]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[14]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[8]), .B(OutData[33]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[46]), .A2(OutData[40]), .ZN(SlicesFromChi[71]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[27]), .A2(OutData[46]), .ZN(SlicesFromChi[76]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[33]), .A2(OutData[27]), .ZN(SlicesFromChi[81]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[39]), .A2(OutData[33]), .ZN(SlicesFromChi[86]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[8]), .ZN(SlicesFromChi[91]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[39]), .A2(OutData[15]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(FreshRand[9]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[96]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[46]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(OutData[15]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(OutData[5]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7), .ZN(SlicesFromChi[2]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[17]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(OutData[11]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A(OutData[11]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[7]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A1(OutData[23]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(OutData[17]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U3 ( 
        .A(OutData[17]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7), .ZN(SlicesFromChi[12]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A1(OutData[4]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A(OutData[23]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A(OutData[23]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[17]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A1(OutData[5]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(OutData[4]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U3 ( 
        .A(OutData[4]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7), .ZN(SlicesFromChi[22]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U2 ( 
        .A1(OutData[11]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A(OutData[5]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U3 ( 
        .A(FreshRand[10]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5), .ZN(SlicesFromChi[27]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A1(OutData[42]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A(OutData[11]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[11]), .ZN(SlicesFromChi[32]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[42]), .A2(OutData[23]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7), .ZN(SlicesFromChi[37]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U3 ( 
        .A1(OutData[29]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(OutData[23]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A(FreshRand[12]), .B(OutData[42]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[30]), .A2(OutData[29]), .ZN(SlicesFromChi[42]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[47]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[30]), .A2(OutData[11]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(FreshRand[14]), .B(OutData[29]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[52]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[36]), .A2(OutData[17]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[10]), .B(OutData[30]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[57]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[48]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[17]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[11]), .B(OutData[36]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[12]), .ZN(SlicesFromChi[62]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[48]), .A2(OutData[4]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[67]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[30]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[4]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[13]), .B(OutData[48]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[36]), .A2(OutData[30]), .ZN(SlicesFromChi[72]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[42]), .A2(OutData[36]), .ZN(SlicesFromChi[77]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[48]), .A2(OutData[42]), .ZN(SlicesFromChi[82]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[29]), .A2(OutData[48]), .ZN(SlicesFromChi[87]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[13]), .ZN(SlicesFromChi[92]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[29]), .A2(OutData[5]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(FreshRand[14]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[97]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[36]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(OutData[5]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(OutData[20]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7), .ZN(SlicesFromChi[3]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[7]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(OutData[1]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A(OutData[1]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[8]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A1(OutData[13]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(OutData[7]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U3 ( 
        .A(OutData[7]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7), .ZN(SlicesFromChi[13]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A1(OutData[19]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A(OutData[13]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A(OutData[13]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[18]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A1(OutData[20]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(OutData[19]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U3 ( 
        .A(OutData[19]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7), .ZN(SlicesFromChi[23]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U2 ( 
        .A1(OutData[1]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A(OutData[20]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U3 ( 
        .A(FreshRand[15]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5), .ZN(SlicesFromChi[28]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A1(OutData[32]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A(OutData[1]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[16]), .ZN(SlicesFromChi[33]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[32]), .A2(OutData[13]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7), .ZN(SlicesFromChi[38]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U3 ( 
        .A1(OutData[44]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(OutData[13]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A(FreshRand[17]), .B(OutData[32]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[45]), .A2(OutData[44]), .ZN(SlicesFromChi[43]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[48]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[45]), .A2(OutData[1]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(FreshRand[19]), .B(OutData[44]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[53]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[26]), .A2(OutData[7]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[15]), .B(OutData[45]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[58]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[38]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[7]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[16]), .B(OutData[26]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[17]), .ZN(SlicesFromChi[63]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[38]), .A2(OutData[19]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[68]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[45]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[19]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[18]), .B(OutData[38]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[26]), .A2(OutData[45]), .ZN(SlicesFromChi[73]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[32]), .A2(OutData[26]), .ZN(SlicesFromChi[78]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[38]), .A2(OutData[32]), .ZN(SlicesFromChi[83]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[44]), .A2(OutData[38]), .ZN(SlicesFromChi[88]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[18]), .ZN(SlicesFromChi[93]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[44]), .A2(OutData[20]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(FreshRand[19]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[98]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[26]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(OutData[20]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(OutData[10]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7), .ZN(SlicesFromChi[4]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[22]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(OutData[16]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A(OutData[16]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[9]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A1(OutData[3]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(OutData[22]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U3 ( 
        .A(OutData[22]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7), .ZN(SlicesFromChi[14]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A1(OutData[9]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A(OutData[3]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A(OutData[3]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[19]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A1(OutData[10]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(OutData[9]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U3 ( 
        .A(OutData[9]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7), .ZN(SlicesFromChi[24]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U2 ( 
        .A1(OutData[16]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A(OutData[10]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U3 ( 
        .A(FreshRand[20]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5), .ZN(SlicesFromChi[29]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A1(OutData[47]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A(OutData[16]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[21]), .ZN(SlicesFromChi[34]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[47]), .A2(OutData[3]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7), .ZN(SlicesFromChi[39]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U3 ( 
        .A1(OutData[34]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(OutData[3]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A(FreshRand[22]), .B(OutData[47]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[35]), .A2(OutData[34]), .ZN(SlicesFromChi[44]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[49]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[35]), .A2(OutData[16]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(FreshRand[24]), .B(OutData[34]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[54]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[41]), .A2(OutData[22]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[20]), .B(OutData[35]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[59]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[28]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[22]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[21]), .B(OutData[41]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[22]), .ZN(SlicesFromChi[64]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[28]), .A2(OutData[9]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[69]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[35]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[9]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[23]), .B(OutData[28]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[41]), .A2(OutData[35]), .ZN(SlicesFromChi[74]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[47]), .A2(OutData[41]), .ZN(SlicesFromChi[79]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[28]), .A2(OutData[47]), .ZN(SlicesFromChi[84]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[34]), .A2(OutData[28]), .ZN(SlicesFromChi[89]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[23]), .ZN(SlicesFromChi[94]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[34]), .A2(OutData[10]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(FreshRand[24]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[99]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[41]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(OutData[10]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n4) );
  OAI221_X1 KECCAK_CONTROL_U33 ( .B1(KECCAK_CONTROL_n6), .B2(
        KECCAK_CONTROL_n62), .C1(KECCAK_CONTROL_n6), .C2(KECCAK_CONTROL_n61), 
        .A(KECCAK_CONTROL_n60), .ZN(KECCAK_CONTROL_n34) );
  NAND3_X1 KECCAK_CONTROL_U32 ( .A1(KECCAK_CONTROL_n59), .A2(
        KECCAK_CONTROL_n58), .A3(KECCAK_CONTROL_n6), .ZN(KECCAK_CONTROL_n60)
         );
  OAI22_X1 KECCAK_CONTROL_U31 ( .A1(KECCAK_CONTROL_n27), .A2(
        KECCAK_CONTROL_n62), .B1(KECCAK_CONTROL_n57), .B2(KECCAK_CONTROL_n61), 
        .ZN(KECCAK_CONTROL_n35) );
  NAND2_X1 KECCAK_CONTROL_U30 ( .A1(KECCAK_CONTROL_n59), .A2(
        KECCAK_CONTROL_n27), .ZN(KECCAK_CONTROL_n61) );
  OR2_X1 KECCAK_CONTROL_U29 ( .A1(KECCAK_CONTROL_n40), .A2(KECCAK_CONTROL_n31), 
        .ZN(KECCAK_CONTROL_n57) );
  AOI21_X1 KECCAK_CONTROL_U28 ( .B1(KECCAK_CONTROL_n59), .B2(
        KECCAK_CONTROL_n31), .A(KECCAK_CONTROL_n56), .ZN(KECCAK_CONTROL_n62)
         );
  OAI22_X1 KECCAK_CONTROL_U27 ( .A1(KECCAK_CONTROL_n31), .A2(
        KECCAK_CONTROL_n55), .B1(KECCAK_CONTROL_n54), .B2(KECCAK_CONTROL_n40), 
        .ZN(KECCAK_CONTROL_n36) );
  NAND2_X1 KECCAK_CONTROL_U26 ( .A1(KECCAK_CONTROL_n59), .A2(
        KECCAK_CONTROL_n31), .ZN(KECCAK_CONTROL_n54) );
  INV_X1 KECCAK_CONTROL_U25 ( .A(KECCAK_CONTROL_n53), .ZN(KECCAK_CONTROL_n59)
         );
  INV_X1 KECCAK_CONTROL_U24 ( .A(KECCAK_CONTROL_n56), .ZN(KECCAK_CONTROL_n55)
         );
  OAI21_X1 KECCAK_CONTROL_U23 ( .B1(Reset), .B2(
        KECCAK_CONTROL_RoundCountxDP_0_), .A(KECCAK_CONTROL_n52), .ZN(
        KECCAK_CONTROL_n56) );
  AOI22_X1 KECCAK_CONTROL_U22 ( .A1(KECCAK_CONTROL_RoundCountxDP_0_), .A2(
        KECCAK_CONTROL_n52), .B1(KECCAK_CONTROL_n53), .B2(KECCAK_CONTROL_n40), 
        .ZN(KECCAK_CONTROL_n37) );
  OAI22_X1 KECCAK_CONTROL_U21 ( .A1(KECCAK_CONTROL_n32), .A2(
        KECCAK_CONTROL_n52), .B1(KECCAK_CONTROL_n51), .B2(KECCAK_CONTROL_n53), 
        .ZN(KECCAK_CONTROL_n38) );
  NAND2_X1 KECCAK_CONTROL_U20 ( .A1(KECCAK_CONTROL_n42), .A2(
        KECCAK_CONTROL_n52), .ZN(KECCAK_CONTROL_n53) );
  NAND3_X1 KECCAK_CONTROL_U19 ( .A1(KECCAK_CONTROL_n42), .A2(
        KECCAK_CONTROL_n50), .A3(KECCAK_CONTROL_n49), .ZN(KECCAK_CONTROL_n52)
         );
  AOI21_X1 KECCAK_CONTROL_U18 ( .B1(KECCAK_CONTROL_n39), .B2(
        KECCAK_CONTROL_n50), .A(Reset), .ZN(KECCAK_CONTROL_n48) );
  AOI21_X1 KECCAK_CONTROL_U17 ( .B1(KECCAK_CONTROL_n14), .B2(
        KECCAK_CONTROL_n47), .A(Reset), .ZN(KECCAK_CONTROL_n29) );
  INV_X1 KECCAK_CONTROL_U16 ( .A(KECCAK_CONTROL_n46), .ZN(KECCAK_CONTROL_n47)
         );
  AOI221_X1 KECCAK_CONTROL_U15 ( .B1(KECCAK_CONTROL_n26), .B2(
        KECCAK_CONTROL_n50), .C1(KECCAK_CONTROL_n46), .C2(KECCAK_CONTROL_n50), 
        .A(Reset), .ZN(KECCAK_CONTROL_n28) );
  NOR2_X1 KECCAK_CONTROL_U14 ( .A1(KECCAK_CONTROL_n5), .A2(KECCAK_CONTROL_n49), 
        .ZN(KECCAK_CONTROL_n46) );
  NAND3_X1 KECCAK_CONTROL_U13 ( .A1(KECCAK_CONTROL_n41), .A2(
        KECCAK_CONTROL_n15), .A3(KECCAK_CONTROL_n14), .ZN(KECCAK_CONTROL_n49)
         );
  NAND3_X1 KECCAK_CONTROL_U12 ( .A1(KECCAK_CONTROL_n39), .A2(
        KECCAK_CONTROL_n14), .A3(KECCAK_CONTROL_n26), .ZN(KECCAK_CONTROL_n50)
         );
  NOR3_X1 KECCAK_CONTROL_U11 ( .A1(KECCAK_CONTROL_n14), .A2(KECCAK_CONTROL_n39), .A3(KECCAK_CONTROL_n41), .ZN(Ready) );
  AOI21_X1 KECCAK_CONTROL_U10 ( .B1(KECCAK_CONTROL_n51), .B2(
        KECCAK_CONTROL_n45), .A(Reset), .ZN(KECCAK_CONTROL_N32) );
  INV_X1 KECCAK_CONTROL_U9 ( .A(KECCAK_CONTROL_n44), .ZN(KECCAK_CONTROL_n45)
         );
  AOI211_X1 KECCAK_CONTROL_U8 ( .C1(KECCAK_CONTROL_n27), .C2(
        KECCAK_CONTROL_n31), .A(KECCAK_CONTROL_n58), .B(KECCAK_CONTROL_n6), 
        .ZN(KECCAK_CONTROL_n44) );
  XNOR2_X1 KECCAK_CONTROL_U7 ( .A(KECCAK_CONTROL_n43), .B(KECCAK_CONTROL_n32), 
        .ZN(KECCAK_CONTROL_n51) );
  NAND2_X1 KECCAK_CONTROL_U6 ( .A1(KECCAK_CONTROL_RoundCountxDP_3_), .A2(
        KECCAK_CONTROL_n58), .ZN(KECCAK_CONTROL_n43) );
  NOR3_X1 KECCAK_CONTROL_U5 ( .A1(KECCAK_CONTROL_n31), .A2(KECCAK_CONTROL_n27), 
        .A3(KECCAK_CONTROL_n40), .ZN(KECCAK_CONTROL_n58) );
  NOR2_X1 KECCAK_CONTROL_U4 ( .A1(Reset), .A2(KECCAK_CONTROL_n5), .ZN(
        Lastround) );
  INV_X1 KECCAK_CONTROL_U3 ( .A(Reset), .ZN(KECCAK_CONTROL_n42) );
  DFF_X1 KECCAK_CONTROL_CtrlStatexDP_reg_0_ ( .D(KECCAK_CONTROL_n48), .CK(
        Clock), .Q(KECCAK_CONTROL_n15), .QN(KECCAK_CONTROL_n39) );
  DFF_X1 KECCAK_CONTROL_RoundCountxDP_reg_0_ ( .D(KECCAK_CONTROL_n37), .CK(
        Clock), .Q(KECCAK_CONTROL_RoundCountxDP_0_), .QN(KECCAK_CONTROL_n40)
         );
  DFF_X1 KECCAK_CONTROL_RoundCountxDP_reg_1_ ( .D(KECCAK_CONTROL_n36), .CK(
        Clock), .Q(KECCAK_CONTROL_RoundCountxDP_1_), .QN(KECCAK_CONTROL_n31)
         );
  DFF_X1 KECCAK_CONTROL_RoundCountxDP_reg_2_ ( .D(KECCAK_CONTROL_n35), .CK(
        Clock), .Q(KECCAK_CONTROL_RoundCountxDP_2_), .QN(KECCAK_CONTROL_n27)
         );
  DFF_X1 KECCAK_CONTROL_RoundCountxDP_reg_3_ ( .D(KECCAK_CONTROL_n34), .CK(
        Clock), .Q(KECCAK_CONTROL_RoundCountxDP_3_), .QN(KECCAK_CONTROL_n6) );
  DFF_X1 KECCAK_CONTROL_RoundCountxDP_reg_4_ ( .D(KECCAK_CONTROL_n38), .CK(
        Clock), .Q(KECCAK_CONTROL_RoundCountxDP_4_), .QN(KECCAK_CONTROL_n32)
         );
  DFF_X1 KECCAK_CONTROL_CtrlStatexDP_reg_1_ ( .D(KECCAK_CONTROL_n28), .CK(
        Clock), .Q(KECCAK_CONTROL_n41), .QN(KECCAK_CONTROL_n26) );
  DFF_X1 KECCAK_CONTROL_CtrlStatexDP_reg_2_ ( .D(KECCAK_CONTROL_n29), .CK(
        Clock), .Q(), .QN(KECCAK_CONTROL_n14) );
  DFF_X1 KECCAK_CONTROL_RoundCountLastxDP_reg ( .D(KECCAK_CONTROL_N32), .CK(
        Clock), .Q(), .QN(KECCAK_CONTROL_n5) );
  AOI221_X1 KECCAK_CONTROL_RC_GEN_U4 ( .B1(KECCAK_CONTROL_RoundCountxDP_0_), 
        .B2(KECCAK_CONTROL_RC_GEN_n3), .C1(KECCAK_CONTROL_RC_GEN_n2), .C2(
        KECCAK_CONTROL_RC_GEN_n3), .A(KECCAK_CONTROL_RoundCountxDP_4_), .ZN(
        IotaRC_0_) );
  XOR2_X1 KECCAK_CONTROL_RC_GEN_U3 ( .A(KECCAK_CONTROL_RoundCountxDP_1_), .B(
        KECCAK_CONTROL_RoundCountxDP_3_), .Z(KECCAK_CONTROL_RC_GEN_n2) );
  INV_X1 KECCAK_CONTROL_RC_GEN_U2 ( .A(KECCAK_CONTROL_RoundCountxDP_2_), .ZN(
        KECCAK_CONTROL_RC_GEN_n3) );
endmodule

