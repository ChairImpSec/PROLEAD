
module circuit ( Clock, Reset, InData, FreshRand, Ready, OutData );
  input [74:0] InData;
  input [74:0] FreshRand;
  output [74:0] OutData;
  input Clock, Reset;
  output Ready;
  wire   Lastround, IotaRC_0_, n2, n3, n4,
         all_mux_linear_0__MUX_theta_state_inst_n218,
         all_mux_linear_0__MUX_theta_state_inst_n217,
         all_mux_linear_0__MUX_theta_state_inst_n216,
         all_mux_linear_0__MUX_theta_state_inst_n215,
         all_mux_linear_0__MUX_theta_state_inst_n214,
         all_mux_linear_0__MUX_theta_state_inst_n213,
         all_mux_linear_0__MUX_theta_state_inst_n212,
         all_mux_linear_0__MUX_theta_state_inst_n211,
         all_mux_linear_0__MUX_theta_state_inst_n210,
         all_mux_linear_0__MUX_theta_state_inst_n209,
         all_mux_linear_0__MUX_theta_state_inst_n208,
         all_mux_linear_0__MUX_theta_state_inst_n207,
         all_mux_linear_0__MUX_theta_state_inst_n206,
         all_mux_linear_0__MUX_theta_state_inst_n205,
         all_mux_linear_0__MUX_theta_state_inst_n204,
         all_mux_linear_0__MUX_theta_state_inst_n203,
         all_mux_linear_0__MUX_theta_state_inst_n202,
         all_mux_linear_0__MUX_theta_state_inst_n201,
         all_mux_linear_0__MUX_theta_state_inst_n200,
         all_mux_linear_0__MUX_theta_state_inst_n199,
         all_mux_linear_0__MUX_theta_state_inst_n198,
         all_mux_linear_0__MUX_theta_state_inst_n197,
         all_mux_linear_0__MUX_theta_state_inst_n196,
         all_mux_linear_0__MUX_theta_state_inst_n195,
         all_mux_linear_0__MUX_theta_state_inst_n194,
         all_mux_linear_0__MUX_theta_state_inst_n193,
         all_mux_linear_0__MUX_theta_state_inst_n192,
         all_mux_linear_0__MUX_theta_state_inst_n191,
         all_mux_linear_0__MUX_theta_state_inst_n190,
         all_mux_linear_0__MUX_theta_state_inst_n189,
         all_mux_linear_0__MUX_theta_state_inst_n188,
         all_mux_linear_0__MUX_theta_state_inst_n187,
         all_mux_linear_0__MUX_theta_state_inst_n186,
         all_mux_linear_0__MUX_theta_state_inst_n185,
         all_mux_linear_0__MUX_theta_state_inst_n184,
         all_mux_linear_0__MUX_theta_state_inst_n183,
         all_mux_linear_0__MUX_theta_state_inst_n182,
         all_mux_linear_0__MUX_theta_state_inst_n181,
         all_mux_linear_0__MUX_theta_state_inst_n180,
         all_mux_linear_0__MUX_theta_state_inst_n179,
         all_mux_linear_0__MUX_theta_state_inst_n178,
         all_mux_linear_0__MUX_theta_state_inst_n177,
         all_mux_linear_0__MUX_theta_state_inst_n176,
         all_mux_linear_0__MUX_theta_state_inst_n175,
         all_mux_linear_0__MUX_theta_state_inst_n174,
         all_mux_linear_0__MUX_theta_state_inst_n173,
         all_mux_linear_0__MUX_theta_state_inst_n172,
         all_mux_linear_0__MUX_theta_state_inst_n171,
         all_mux_linear_0__MUX_theta_state_inst_n170,
         all_mux_linear_0__MUX_theta_state_inst_n169,
         all_mux_linear_0__MUX_theta_state_inst_n168,
         all_mux_linear_0__MUX_theta_state_inst_n167,
         all_mux_linear_0__MUX_theta_state_inst_n166,
         all_mux_linear_0__MUX_theta_state_inst_n165,
         all_mux_linear_0__MUX_theta_state_inst_n164,
         all_mux_linear_0__MUX_theta_state_inst_n163,
         all_mux_linear_0__MUX_theta_state_inst_n162,
         all_mux_linear_0__MUX_theta_state_inst_n161,
         all_mux_linear_0__MUX_theta_state_inst_n160,
         all_mux_linear_0__MUX_theta_state_inst_n159,
         all_mux_linear_0__MUX_theta_state_inst_n158,
         all_mux_linear_0__MUX_theta_state_inst_n157,
         all_mux_linear_0__MUX_theta_state_inst_n156,
         all_mux_linear_0__MUX_theta_state_inst_n155,
         all_mux_linear_0__MUX_theta_state_inst_n154,
         all_mux_linear_0__MUX_theta_state_inst_n153,
         all_mux_linear_0__MUX_theta_state_inst_n152,
         all_mux_linear_0__MUX_theta_state_inst_n151,
         all_mux_linear_0__MUX_theta_state_inst_n150,
         all_mux_linear_0__MUX_theta_state_inst_n149,
         all_mux_linear_0__MUX_theta_state_inst_n148,
         all_mux_linear_0__MUX_theta_state_inst_n147,
         all_mux_linear_0__MUX_theta_state_inst_n146,
         all_mux_linear_0__MUX_theta_state_inst_n145,
         all_mux_linear_0__MUX_theta_state_inst_n144,
         all_mux_linear_0__MUX_theta_state_inst_n143,
         all_mux_linear_0__MUX_theta_state_inst_n142,
         all_mux_linear_0__MUX_theta_state_inst_n141,
         all_mux_linear_0__MUX_theta_state_inst_n140,
         all_mux_linear_0__MUX_theta_state_inst_n139,
         all_mux_linear_0__MUX_theta_state_inst_n138,
         all_mux_linear_0__MUX_theta_state_inst_n137,
         all_mux_linear_0__MUX_theta_state_inst_n136,
         all_mux_linear_0__MUX_theta_state_inst_n135,
         all_mux_linear_0__MUX_theta_state_inst_n134,
         all_mux_linear_0__MUX_theta_state_inst_n133,
         all_mux_linear_0__MUX_theta_state_inst_n132,
         all_mux_linear_0__MUX_theta_state_inst_n131,
         all_mux_linear_0__MUX_theta_state_inst_n130,
         all_mux_linear_1__MUX_theta_state_inst_n336,
         all_mux_linear_1__MUX_theta_state_inst_n335,
         all_mux_linear_1__MUX_theta_state_inst_n334,
         all_mux_linear_1__MUX_theta_state_inst_n333,
         all_mux_linear_1__MUX_theta_state_inst_n332,
         all_mux_linear_1__MUX_theta_state_inst_n331,
         all_mux_linear_1__MUX_theta_state_inst_n330,
         all_mux_linear_1__MUX_theta_state_inst_n329,
         all_mux_linear_1__MUX_theta_state_inst_n328,
         all_mux_linear_1__MUX_theta_state_inst_n327,
         all_mux_linear_1__MUX_theta_state_inst_n326,
         all_mux_linear_1__MUX_theta_state_inst_n325,
         all_mux_linear_1__MUX_theta_state_inst_n324,
         all_mux_linear_1__MUX_theta_state_inst_n323,
         all_mux_linear_1__MUX_theta_state_inst_n322,
         all_mux_linear_1__MUX_theta_state_inst_n321,
         all_mux_linear_1__MUX_theta_state_inst_n320,
         all_mux_linear_1__MUX_theta_state_inst_n319,
         all_mux_linear_1__MUX_theta_state_inst_n318,
         all_mux_linear_1__MUX_theta_state_inst_n317,
         all_mux_linear_1__MUX_theta_state_inst_n316,
         all_mux_linear_1__MUX_theta_state_inst_n315,
         all_mux_linear_1__MUX_theta_state_inst_n314,
         all_mux_linear_1__MUX_theta_state_inst_n313,
         all_mux_linear_1__MUX_theta_state_inst_n312,
         all_mux_linear_1__MUX_theta_state_inst_n311,
         all_mux_linear_1__MUX_theta_state_inst_n310,
         all_mux_linear_1__MUX_theta_state_inst_n309,
         all_mux_linear_1__MUX_theta_state_inst_n308,
         all_mux_linear_1__MUX_theta_state_inst_n307,
         all_mux_linear_1__MUX_theta_state_inst_n306,
         all_mux_linear_1__MUX_theta_state_inst_n305,
         all_mux_linear_1__MUX_theta_state_inst_n304,
         all_mux_linear_1__MUX_theta_state_inst_n303,
         all_mux_linear_1__MUX_theta_state_inst_n302,
         all_mux_linear_1__MUX_theta_state_inst_n301,
         all_mux_linear_1__MUX_theta_state_inst_n300,
         all_mux_linear_1__MUX_theta_state_inst_n299,
         all_mux_linear_1__MUX_theta_state_inst_n298,
         all_mux_linear_1__MUX_theta_state_inst_n297,
         all_mux_linear_1__MUX_theta_state_inst_n296,
         all_mux_linear_1__MUX_theta_state_inst_n295,
         all_mux_linear_1__MUX_theta_state_inst_n294,
         all_mux_linear_1__MUX_theta_state_inst_n293,
         all_mux_linear_1__MUX_theta_state_inst_n292,
         all_mux_linear_1__MUX_theta_state_inst_n291,
         all_mux_linear_1__MUX_theta_state_inst_n290,
         all_mux_linear_1__MUX_theta_state_inst_n289,
         all_mux_linear_1__MUX_theta_state_inst_n288,
         all_mux_linear_1__MUX_theta_state_inst_n287,
         all_mux_linear_1__MUX_theta_state_inst_n286,
         all_mux_linear_1__MUX_theta_state_inst_n285,
         all_mux_linear_1__MUX_theta_state_inst_n284,
         all_mux_linear_1__MUX_theta_state_inst_n283,
         all_mux_linear_1__MUX_theta_state_inst_n282,
         all_mux_linear_1__MUX_theta_state_inst_n281,
         all_mux_linear_1__MUX_theta_state_inst_n280,
         all_mux_linear_1__MUX_theta_state_inst_n279,
         all_mux_linear_1__MUX_theta_state_inst_n278,
         all_mux_linear_1__MUX_theta_state_inst_n277,
         all_mux_linear_1__MUX_theta_state_inst_n276,
         all_mux_linear_1__MUX_theta_state_inst_n275,
         all_mux_linear_1__MUX_theta_state_inst_n274,
         all_mux_linear_1__MUX_theta_state_inst_n273,
         all_mux_linear_1__MUX_theta_state_inst_n272,
         all_mux_linear_1__MUX_theta_state_inst_n271,
         all_mux_linear_1__MUX_theta_state_inst_n270,
         all_mux_linear_1__MUX_theta_state_inst_n269,
         all_mux_linear_1__MUX_theta_state_inst_n268,
         all_mux_linear_1__MUX_theta_state_inst_n267,
         all_mux_linear_1__MUX_theta_state_inst_n266,
         all_mux_linear_1__MUX_theta_state_inst_n265,
         all_mux_linear_1__MUX_theta_state_inst_n264,
         all_mux_linear_1__MUX_theta_state_inst_n263,
         all_mux_linear_1__MUX_theta_state_inst_n262,
         all_mux_linear_1__MUX_theta_state_inst_n261,
         all_mux_linear_1__MUX_theta_state_inst_n260,
         all_mux_linear_1__MUX_theta_state_inst_n259,
         all_mux_linear_1__MUX_theta_state_inst_n258,
         all_mux_linear_1__MUX_theta_state_inst_n257,
         all_mux_linear_1__MUX_theta_state_inst_n256,
         all_mux_linear_1__MUX_theta_state_inst_n255,
         all_mux_linear_1__MUX_theta_state_inst_n254,
         all_mux_linear_1__MUX_theta_state_inst_n253,
         all_mux_linear_1__MUX_theta_state_inst_n252,
         all_mux_linear_1__MUX_theta_state_inst_n251,
         all_mux_linear_1__MUX_theta_state_inst_n250,
         all_mux_linear_1__MUX_theta_state_inst_n249,
         all_mux_linear_1__MUX_theta_state_inst_n248,
         all_mux_linear_1__MUX_theta_state_inst_n247,
         all_mux_linear_1__MUX_theta_state_inst_n246,
         all_mux_linear_1__MUX_theta_state_inst_n245,
         all_mux_linear_1__MUX_theta_state_inst_n244,
         all_mux_linear_1__MUX_theta_state_inst_n243,
         all_mux_linear_1__MUX_theta_state_inst_n242,
         all_mux_linear_1__MUX_theta_state_inst_n241,
         all_mux_linear_1__MUX_theta_state_inst_n240,
         all_mux_linear_1__MUX_theta_state_inst_n239,
         all_mux_linear_1__MUX_theta_state_inst_n238,
         all_mux_linear_1__MUX_theta_state_inst_n237,
         all_mux_linear_1__MUX_theta_state_inst_n236,
         all_mux_linear_1__MUX_theta_state_inst_n235,
         all_mux_linear_1__MUX_theta_state_inst_n234,
         all_mux_linear_1__MUX_theta_state_inst_n233,
         all_mux_linear_1__MUX_theta_state_inst_n232,
         all_mux_linear_1__MUX_theta_state_inst_n231,
         all_mux_linear_1__MUX_theta_state_inst_n230,
         all_mux_linear_2__MUX_theta_state_inst_n335,
         all_mux_linear_2__MUX_theta_state_inst_n334,
         all_mux_linear_2__MUX_theta_state_inst_n333,
         all_mux_linear_2__MUX_theta_state_inst_n332,
         all_mux_linear_2__MUX_theta_state_inst_n331,
         all_mux_linear_2__MUX_theta_state_inst_n330,
         all_mux_linear_2__MUX_theta_state_inst_n329,
         all_mux_linear_2__MUX_theta_state_inst_n328,
         all_mux_linear_2__MUX_theta_state_inst_n327,
         all_mux_linear_2__MUX_theta_state_inst_n326,
         all_mux_linear_2__MUX_theta_state_inst_n325,
         all_mux_linear_2__MUX_theta_state_inst_n324,
         all_mux_linear_2__MUX_theta_state_inst_n323,
         all_mux_linear_2__MUX_theta_state_inst_n322,
         all_mux_linear_2__MUX_theta_state_inst_n321,
         all_mux_linear_2__MUX_theta_state_inst_n320,
         all_mux_linear_2__MUX_theta_state_inst_n319,
         all_mux_linear_2__MUX_theta_state_inst_n318,
         all_mux_linear_2__MUX_theta_state_inst_n317,
         all_mux_linear_2__MUX_theta_state_inst_n316,
         all_mux_linear_2__MUX_theta_state_inst_n315,
         all_mux_linear_2__MUX_theta_state_inst_n314,
         all_mux_linear_2__MUX_theta_state_inst_n313,
         all_mux_linear_2__MUX_theta_state_inst_n312,
         all_mux_linear_2__MUX_theta_state_inst_n311,
         all_mux_linear_2__MUX_theta_state_inst_n310,
         all_mux_linear_2__MUX_theta_state_inst_n309,
         all_mux_linear_2__MUX_theta_state_inst_n308,
         all_mux_linear_2__MUX_theta_state_inst_n307,
         all_mux_linear_2__MUX_theta_state_inst_n306,
         all_mux_linear_2__MUX_theta_state_inst_n305,
         all_mux_linear_2__MUX_theta_state_inst_n304,
         all_mux_linear_2__MUX_theta_state_inst_n303,
         all_mux_linear_2__MUX_theta_state_inst_n302,
         all_mux_linear_2__MUX_theta_state_inst_n301,
         all_mux_linear_2__MUX_theta_state_inst_n300,
         all_mux_linear_2__MUX_theta_state_inst_n299,
         all_mux_linear_2__MUX_theta_state_inst_n298,
         all_mux_linear_2__MUX_theta_state_inst_n297,
         all_mux_linear_2__MUX_theta_state_inst_n296,
         all_mux_linear_2__MUX_theta_state_inst_n295,
         all_mux_linear_2__MUX_theta_state_inst_n294,
         all_mux_linear_2__MUX_theta_state_inst_n293,
         all_mux_linear_2__MUX_theta_state_inst_n292,
         all_mux_linear_2__MUX_theta_state_inst_n291,
         all_mux_linear_2__MUX_theta_state_inst_n290,
         all_mux_linear_2__MUX_theta_state_inst_n289,
         all_mux_linear_2__MUX_theta_state_inst_n288,
         all_mux_linear_2__MUX_theta_state_inst_n287,
         all_mux_linear_2__MUX_theta_state_inst_n286,
         all_mux_linear_2__MUX_theta_state_inst_n285,
         all_mux_linear_2__MUX_theta_state_inst_n284,
         all_mux_linear_2__MUX_theta_state_inst_n283,
         all_mux_linear_2__MUX_theta_state_inst_n282,
         all_mux_linear_2__MUX_theta_state_inst_n281,
         all_mux_linear_2__MUX_theta_state_inst_n280,
         all_mux_linear_2__MUX_theta_state_inst_n279,
         all_mux_linear_2__MUX_theta_state_inst_n278,
         all_mux_linear_2__MUX_theta_state_inst_n277,
         all_mux_linear_2__MUX_theta_state_inst_n276,
         all_mux_linear_2__MUX_theta_state_inst_n275,
         all_mux_linear_2__MUX_theta_state_inst_n274,
         all_mux_linear_2__MUX_theta_state_inst_n273,
         all_mux_linear_2__MUX_theta_state_inst_n272,
         all_mux_linear_2__MUX_theta_state_inst_n271,
         all_mux_linear_2__MUX_theta_state_inst_n270,
         all_mux_linear_2__MUX_theta_state_inst_n269,
         all_mux_linear_2__MUX_theta_state_inst_n268,
         all_mux_linear_2__MUX_theta_state_inst_n267,
         all_mux_linear_2__MUX_theta_state_inst_n266,
         all_mux_linear_2__MUX_theta_state_inst_n265,
         all_mux_linear_2__MUX_theta_state_inst_n264,
         all_mux_linear_2__MUX_theta_state_inst_n263,
         all_mux_linear_2__MUX_theta_state_inst_n262,
         all_mux_linear_2__MUX_theta_state_inst_n261,
         all_mux_linear_2__MUX_theta_state_inst_n260,
         all_mux_linear_2__MUX_theta_state_inst_n259,
         all_mux_linear_2__MUX_theta_state_inst_n258,
         all_mux_linear_2__MUX_theta_state_inst_n257,
         all_mux_linear_2__MUX_theta_state_inst_n256,
         all_mux_linear_2__MUX_theta_state_inst_n255,
         all_mux_linear_2__MUX_theta_state_inst_n254,
         all_mux_linear_2__MUX_theta_state_inst_n253,
         all_mux_linear_2__MUX_theta_state_inst_n252,
         all_mux_linear_2__MUX_theta_state_inst_n251,
         all_mux_linear_2__MUX_theta_state_inst_n250,
         all_mux_linear_2__MUX_theta_state_inst_n249,
         all_mux_linear_2__MUX_theta_state_inst_n248,
         all_mux_linear_2__MUX_theta_state_inst_n247,
         all_mux_linear_2__MUX_theta_state_inst_n246,
         all_mux_linear_2__MUX_theta_state_inst_n245,
         all_mux_linear_2__MUX_theta_state_inst_n244,
         all_mux_linear_2__MUX_theta_state_inst_n243,
         all_mux_linear_2__MUX_theta_state_inst_n242,
         all_mux_linear_2__MUX_theta_state_inst_n241,
         all_mux_linear_2__MUX_theta_state_inst_n240,
         all_mux_linear_2__MUX_theta_state_inst_n239,
         all_mux_linear_2__MUX_theta_state_inst_n238,
         all_mux_linear_2__MUX_theta_state_inst_n237,
         all_mux_linear_2__MUX_theta_state_inst_n236,
         all_mux_linear_2__MUX_theta_state_inst_n235,
         all_mux_linear_2__MUX_theta_state_inst_n234,
         all_mux_linear_2__MUX_theta_state_inst_n233,
         all_mux_linear_2__MUX_theta_state_inst_n232,
         all_mux_linear_2__MUX_theta_state_inst_n231,
         all_mux_linear_2__MUX_theta_state_inst_n230,
         all_mux_linear_2__MUX_theta_state_inst_n229,
         all_mux_linear_3__MUX_theta_state_inst_n335,
         all_mux_linear_3__MUX_theta_state_inst_n334,
         all_mux_linear_3__MUX_theta_state_inst_n333,
         all_mux_linear_3__MUX_theta_state_inst_n332,
         all_mux_linear_3__MUX_theta_state_inst_n331,
         all_mux_linear_3__MUX_theta_state_inst_n330,
         all_mux_linear_3__MUX_theta_state_inst_n329,
         all_mux_linear_3__MUX_theta_state_inst_n328,
         all_mux_linear_3__MUX_theta_state_inst_n327,
         all_mux_linear_3__MUX_theta_state_inst_n326,
         all_mux_linear_3__MUX_theta_state_inst_n325,
         all_mux_linear_3__MUX_theta_state_inst_n324,
         all_mux_linear_3__MUX_theta_state_inst_n323,
         all_mux_linear_3__MUX_theta_state_inst_n322,
         all_mux_linear_3__MUX_theta_state_inst_n321,
         all_mux_linear_3__MUX_theta_state_inst_n320,
         all_mux_linear_3__MUX_theta_state_inst_n319,
         all_mux_linear_3__MUX_theta_state_inst_n318,
         all_mux_linear_3__MUX_theta_state_inst_n317,
         all_mux_linear_3__MUX_theta_state_inst_n316,
         all_mux_linear_3__MUX_theta_state_inst_n315,
         all_mux_linear_3__MUX_theta_state_inst_n314,
         all_mux_linear_3__MUX_theta_state_inst_n313,
         all_mux_linear_3__MUX_theta_state_inst_n312,
         all_mux_linear_3__MUX_theta_state_inst_n311,
         all_mux_linear_3__MUX_theta_state_inst_n310,
         all_mux_linear_3__MUX_theta_state_inst_n309,
         all_mux_linear_3__MUX_theta_state_inst_n308,
         all_mux_linear_3__MUX_theta_state_inst_n307,
         all_mux_linear_3__MUX_theta_state_inst_n306,
         all_mux_linear_3__MUX_theta_state_inst_n305,
         all_mux_linear_3__MUX_theta_state_inst_n304,
         all_mux_linear_3__MUX_theta_state_inst_n303,
         all_mux_linear_3__MUX_theta_state_inst_n302,
         all_mux_linear_3__MUX_theta_state_inst_n301,
         all_mux_linear_3__MUX_theta_state_inst_n300,
         all_mux_linear_3__MUX_theta_state_inst_n299,
         all_mux_linear_3__MUX_theta_state_inst_n298,
         all_mux_linear_3__MUX_theta_state_inst_n297,
         all_mux_linear_3__MUX_theta_state_inst_n296,
         all_mux_linear_3__MUX_theta_state_inst_n295,
         all_mux_linear_3__MUX_theta_state_inst_n294,
         all_mux_linear_3__MUX_theta_state_inst_n293,
         all_mux_linear_3__MUX_theta_state_inst_n292,
         all_mux_linear_3__MUX_theta_state_inst_n291,
         all_mux_linear_3__MUX_theta_state_inst_n290,
         all_mux_linear_3__MUX_theta_state_inst_n289,
         all_mux_linear_3__MUX_theta_state_inst_n288,
         all_mux_linear_3__MUX_theta_state_inst_n287,
         all_mux_linear_3__MUX_theta_state_inst_n286,
         all_mux_linear_3__MUX_theta_state_inst_n285,
         all_mux_linear_3__MUX_theta_state_inst_n284,
         all_mux_linear_3__MUX_theta_state_inst_n283,
         all_mux_linear_3__MUX_theta_state_inst_n282,
         all_mux_linear_3__MUX_theta_state_inst_n281,
         all_mux_linear_3__MUX_theta_state_inst_n280,
         all_mux_linear_3__MUX_theta_state_inst_n279,
         all_mux_linear_3__MUX_theta_state_inst_n278,
         all_mux_linear_3__MUX_theta_state_inst_n277,
         all_mux_linear_3__MUX_theta_state_inst_n276,
         all_mux_linear_3__MUX_theta_state_inst_n275,
         all_mux_linear_3__MUX_theta_state_inst_n274,
         all_mux_linear_3__MUX_theta_state_inst_n273,
         all_mux_linear_3__MUX_theta_state_inst_n272,
         all_mux_linear_3__MUX_theta_state_inst_n271,
         all_mux_linear_3__MUX_theta_state_inst_n270,
         all_mux_linear_3__MUX_theta_state_inst_n269,
         all_mux_linear_3__MUX_theta_state_inst_n268,
         all_mux_linear_3__MUX_theta_state_inst_n267,
         all_mux_linear_3__MUX_theta_state_inst_n266,
         all_mux_linear_3__MUX_theta_state_inst_n265,
         all_mux_linear_3__MUX_theta_state_inst_n264,
         all_mux_linear_3__MUX_theta_state_inst_n263,
         all_mux_linear_3__MUX_theta_state_inst_n262,
         all_mux_linear_3__MUX_theta_state_inst_n261,
         all_mux_linear_3__MUX_theta_state_inst_n260,
         all_mux_linear_3__MUX_theta_state_inst_n259,
         all_mux_linear_3__MUX_theta_state_inst_n258,
         all_mux_linear_3__MUX_theta_state_inst_n257,
         all_mux_linear_3__MUX_theta_state_inst_n256,
         all_mux_linear_3__MUX_theta_state_inst_n255,
         all_mux_linear_3__MUX_theta_state_inst_n254,
         all_mux_linear_3__MUX_theta_state_inst_n253,
         all_mux_linear_3__MUX_theta_state_inst_n252,
         all_mux_linear_3__MUX_theta_state_inst_n251,
         all_mux_linear_3__MUX_theta_state_inst_n250,
         all_mux_linear_3__MUX_theta_state_inst_n249,
         all_mux_linear_3__MUX_theta_state_inst_n248,
         all_mux_linear_3__MUX_theta_state_inst_n247,
         all_mux_linear_3__MUX_theta_state_inst_n246,
         all_mux_linear_3__MUX_theta_state_inst_n245,
         all_mux_linear_3__MUX_theta_state_inst_n244,
         all_mux_linear_3__MUX_theta_state_inst_n243,
         all_mux_linear_3__MUX_theta_state_inst_n242,
         all_mux_linear_3__MUX_theta_state_inst_n241,
         all_mux_linear_3__MUX_theta_state_inst_n240,
         all_mux_linear_3__MUX_theta_state_inst_n239,
         all_mux_linear_3__MUX_theta_state_inst_n238,
         all_mux_linear_3__MUX_theta_state_inst_n237,
         all_mux_linear_3__MUX_theta_state_inst_n236,
         all_mux_linear_3__MUX_theta_state_inst_n235,
         all_mux_linear_3__MUX_theta_state_inst_n234,
         all_mux_linear_3__MUX_theta_state_inst_n233,
         all_mux_linear_3__MUX_theta_state_inst_n232,
         all_mux_linear_3__MUX_theta_state_inst_n231,
         all_mux_linear_3__MUX_theta_state_inst_n230,
         all_mux_linear_3__MUX_theta_state_inst_n229,
         all_mux_linear_4__MUX_theta_state_inst_n318,
         all_mux_linear_4__MUX_theta_state_inst_n317,
         all_mux_linear_4__MUX_theta_state_inst_n316,
         all_mux_linear_4__MUX_theta_state_inst_n315,
         all_mux_linear_4__MUX_theta_state_inst_n314,
         all_mux_linear_4__MUX_theta_state_inst_n313,
         all_mux_linear_4__MUX_theta_state_inst_n312,
         all_mux_linear_4__MUX_theta_state_inst_n311,
         all_mux_linear_4__MUX_theta_state_inst_n310,
         all_mux_linear_4__MUX_theta_state_inst_n309,
         all_mux_linear_4__MUX_theta_state_inst_n308,
         all_mux_linear_4__MUX_theta_state_inst_n307,
         all_mux_linear_4__MUX_theta_state_inst_n306,
         all_mux_linear_4__MUX_theta_state_inst_n305,
         all_mux_linear_4__MUX_theta_state_inst_n304,
         all_mux_linear_4__MUX_theta_state_inst_n303,
         all_mux_linear_4__MUX_theta_state_inst_n302,
         all_mux_linear_4__MUX_theta_state_inst_n301,
         all_mux_linear_4__MUX_theta_state_inst_n300,
         all_mux_linear_4__MUX_theta_state_inst_n299,
         all_mux_linear_4__MUX_theta_state_inst_n298,
         all_mux_linear_4__MUX_theta_state_inst_n297,
         all_mux_linear_4__MUX_theta_state_inst_n296,
         all_mux_linear_4__MUX_theta_state_inst_n295,
         all_mux_linear_4__MUX_theta_state_inst_n294,
         all_mux_linear_4__MUX_theta_state_inst_n293,
         all_mux_linear_4__MUX_theta_state_inst_n292,
         all_mux_linear_4__MUX_theta_state_inst_n291,
         all_mux_linear_4__MUX_theta_state_inst_n290,
         all_mux_linear_4__MUX_theta_state_inst_n289,
         all_mux_linear_4__MUX_theta_state_inst_n288,
         all_mux_linear_4__MUX_theta_state_inst_n287,
         all_mux_linear_4__MUX_theta_state_inst_n286,
         all_mux_linear_4__MUX_theta_state_inst_n285,
         all_mux_linear_4__MUX_theta_state_inst_n284,
         all_mux_linear_4__MUX_theta_state_inst_n283,
         all_mux_linear_4__MUX_theta_state_inst_n282,
         all_mux_linear_4__MUX_theta_state_inst_n281,
         all_mux_linear_4__MUX_theta_state_inst_n280,
         all_mux_linear_4__MUX_theta_state_inst_n279,
         all_mux_linear_4__MUX_theta_state_inst_n278,
         all_mux_linear_4__MUX_theta_state_inst_n277,
         all_mux_linear_4__MUX_theta_state_inst_n276,
         all_mux_linear_4__MUX_theta_state_inst_n275,
         all_mux_linear_4__MUX_theta_state_inst_n274,
         all_mux_linear_4__MUX_theta_state_inst_n273,
         all_mux_linear_4__MUX_theta_state_inst_n272,
         all_mux_linear_4__MUX_theta_state_inst_n271,
         all_mux_linear_4__MUX_theta_state_inst_n270,
         all_mux_linear_4__MUX_theta_state_inst_n269,
         all_mux_linear_4__MUX_theta_state_inst_n268,
         all_mux_linear_4__MUX_theta_state_inst_n267,
         all_mux_linear_4__MUX_theta_state_inst_n266,
         all_mux_linear_4__MUX_theta_state_inst_n265,
         all_mux_linear_4__MUX_theta_state_inst_n264,
         all_mux_linear_4__MUX_theta_state_inst_n263,
         all_mux_linear_4__MUX_theta_state_inst_n262,
         all_mux_linear_4__MUX_theta_state_inst_n261,
         all_mux_linear_4__MUX_theta_state_inst_n260,
         all_mux_linear_4__MUX_theta_state_inst_n259,
         all_mux_linear_4__MUX_theta_state_inst_n258,
         all_mux_linear_4__MUX_theta_state_inst_n257,
         all_mux_linear_4__MUX_theta_state_inst_n256,
         all_mux_linear_4__MUX_theta_state_inst_n255,
         all_mux_linear_4__MUX_theta_state_inst_n254,
         all_mux_linear_4__MUX_theta_state_inst_n253,
         all_mux_linear_4__MUX_theta_state_inst_n252,
         all_mux_linear_4__MUX_theta_state_inst_n251,
         all_mux_linear_4__MUX_theta_state_inst_n250,
         all_mux_linear_4__MUX_theta_state_inst_n249,
         all_mux_linear_4__MUX_theta_state_inst_n248,
         all_mux_linear_4__MUX_theta_state_inst_n247,
         all_mux_linear_4__MUX_theta_state_inst_n246,
         all_mux_linear_4__MUX_theta_state_inst_n245,
         all_mux_linear_4__MUX_theta_state_inst_n244,
         all_mux_linear_4__MUX_theta_state_inst_n243,
         all_mux_linear_4__MUX_theta_state_inst_n242,
         all_mux_linear_4__MUX_theta_state_inst_n241,
         all_mux_linear_4__MUX_theta_state_inst_n240,
         all_mux_linear_4__MUX_theta_state_inst_n239,
         all_mux_linear_4__MUX_theta_state_inst_n238,
         all_mux_linear_4__MUX_theta_state_inst_n237,
         all_mux_linear_4__MUX_theta_state_inst_n236,
         all_mux_linear_4__MUX_theta_state_inst_n235,
         all_mux_linear_4__MUX_theta_state_inst_n234,
         all_mux_linear_4__MUX_theta_state_inst_n233,
         all_mux_linear_4__MUX_theta_state_inst_n232,
         all_mux_linear_4__MUX_theta_state_inst_n231,
         all_mux_linear_4__MUX_theta_state_inst_n230,
         all_mux_linear_5__MUX_theta_state_inst_n336,
         all_mux_linear_5__MUX_theta_state_inst_n335,
         all_mux_linear_5__MUX_theta_state_inst_n334,
         all_mux_linear_5__MUX_theta_state_inst_n333,
         all_mux_linear_5__MUX_theta_state_inst_n332,
         all_mux_linear_5__MUX_theta_state_inst_n331,
         all_mux_linear_5__MUX_theta_state_inst_n330,
         all_mux_linear_5__MUX_theta_state_inst_n329,
         all_mux_linear_5__MUX_theta_state_inst_n328,
         all_mux_linear_5__MUX_theta_state_inst_n327,
         all_mux_linear_5__MUX_theta_state_inst_n326,
         all_mux_linear_5__MUX_theta_state_inst_n325,
         all_mux_linear_5__MUX_theta_state_inst_n324,
         all_mux_linear_5__MUX_theta_state_inst_n323,
         all_mux_linear_5__MUX_theta_state_inst_n322,
         all_mux_linear_5__MUX_theta_state_inst_n321,
         all_mux_linear_5__MUX_theta_state_inst_n320,
         all_mux_linear_5__MUX_theta_state_inst_n319,
         all_mux_linear_5__MUX_theta_state_inst_n318,
         all_mux_linear_5__MUX_theta_state_inst_n317,
         all_mux_linear_5__MUX_theta_state_inst_n316,
         all_mux_linear_5__MUX_theta_state_inst_n315,
         all_mux_linear_5__MUX_theta_state_inst_n314,
         all_mux_linear_5__MUX_theta_state_inst_n313,
         all_mux_linear_5__MUX_theta_state_inst_n312,
         all_mux_linear_5__MUX_theta_state_inst_n311,
         all_mux_linear_5__MUX_theta_state_inst_n310,
         all_mux_linear_5__MUX_theta_state_inst_n309,
         all_mux_linear_5__MUX_theta_state_inst_n308,
         all_mux_linear_5__MUX_theta_state_inst_n307,
         all_mux_linear_5__MUX_theta_state_inst_n306,
         all_mux_linear_5__MUX_theta_state_inst_n305,
         all_mux_linear_5__MUX_theta_state_inst_n304,
         all_mux_linear_5__MUX_theta_state_inst_n303,
         all_mux_linear_5__MUX_theta_state_inst_n302,
         all_mux_linear_5__MUX_theta_state_inst_n301,
         all_mux_linear_5__MUX_theta_state_inst_n300,
         all_mux_linear_5__MUX_theta_state_inst_n299,
         all_mux_linear_5__MUX_theta_state_inst_n298,
         all_mux_linear_5__MUX_theta_state_inst_n297,
         all_mux_linear_5__MUX_theta_state_inst_n296,
         all_mux_linear_5__MUX_theta_state_inst_n295,
         all_mux_linear_5__MUX_theta_state_inst_n294,
         all_mux_linear_5__MUX_theta_state_inst_n293,
         all_mux_linear_5__MUX_theta_state_inst_n292,
         all_mux_linear_5__MUX_theta_state_inst_n291,
         all_mux_linear_5__MUX_theta_state_inst_n290,
         all_mux_linear_5__MUX_theta_state_inst_n289,
         all_mux_linear_5__MUX_theta_state_inst_n288,
         all_mux_linear_5__MUX_theta_state_inst_n287,
         all_mux_linear_5__MUX_theta_state_inst_n286,
         all_mux_linear_5__MUX_theta_state_inst_n285,
         all_mux_linear_5__MUX_theta_state_inst_n284,
         all_mux_linear_5__MUX_theta_state_inst_n283,
         all_mux_linear_5__MUX_theta_state_inst_n282,
         all_mux_linear_5__MUX_theta_state_inst_n281,
         all_mux_linear_5__MUX_theta_state_inst_n280,
         all_mux_linear_5__MUX_theta_state_inst_n279,
         all_mux_linear_5__MUX_theta_state_inst_n278,
         all_mux_linear_5__MUX_theta_state_inst_n277,
         all_mux_linear_5__MUX_theta_state_inst_n276,
         all_mux_linear_5__MUX_theta_state_inst_n275,
         all_mux_linear_5__MUX_theta_state_inst_n274,
         all_mux_linear_5__MUX_theta_state_inst_n273,
         all_mux_linear_5__MUX_theta_state_inst_n272,
         all_mux_linear_5__MUX_theta_state_inst_n271,
         all_mux_linear_5__MUX_theta_state_inst_n270,
         all_mux_linear_5__MUX_theta_state_inst_n269,
         all_mux_linear_5__MUX_theta_state_inst_n268,
         all_mux_linear_5__MUX_theta_state_inst_n267,
         all_mux_linear_5__MUX_theta_state_inst_n266,
         all_mux_linear_5__MUX_theta_state_inst_n265,
         all_mux_linear_5__MUX_theta_state_inst_n264,
         all_mux_linear_5__MUX_theta_state_inst_n263,
         all_mux_linear_5__MUX_theta_state_inst_n262,
         all_mux_linear_5__MUX_theta_state_inst_n261,
         all_mux_linear_5__MUX_theta_state_inst_n260,
         all_mux_linear_5__MUX_theta_state_inst_n259,
         all_mux_linear_5__MUX_theta_state_inst_n258,
         all_mux_linear_5__MUX_theta_state_inst_n257,
         all_mux_linear_5__MUX_theta_state_inst_n256,
         all_mux_linear_5__MUX_theta_state_inst_n255,
         all_mux_linear_5__MUX_theta_state_inst_n254,
         all_mux_linear_5__MUX_theta_state_inst_n253,
         all_mux_linear_5__MUX_theta_state_inst_n252,
         all_mux_linear_5__MUX_theta_state_inst_n251,
         all_mux_linear_5__MUX_theta_state_inst_n250,
         all_mux_linear_5__MUX_theta_state_inst_n249,
         all_mux_linear_5__MUX_theta_state_inst_n248,
         all_mux_linear_5__MUX_theta_state_inst_n247,
         all_mux_linear_5__MUX_theta_state_inst_n246,
         all_mux_linear_5__MUX_theta_state_inst_n245,
         all_mux_linear_5__MUX_theta_state_inst_n244,
         all_mux_linear_5__MUX_theta_state_inst_n243,
         all_mux_linear_5__MUX_theta_state_inst_n242,
         all_mux_linear_5__MUX_theta_state_inst_n241,
         all_mux_linear_5__MUX_theta_state_inst_n240,
         all_mux_linear_5__MUX_theta_state_inst_n239,
         all_mux_linear_5__MUX_theta_state_inst_n238,
         all_mux_linear_5__MUX_theta_state_inst_n237,
         all_mux_linear_5__MUX_theta_state_inst_n236,
         all_mux_linear_5__MUX_theta_state_inst_n235,
         all_mux_linear_5__MUX_theta_state_inst_n234,
         all_mux_linear_5__MUX_theta_state_inst_n233,
         all_mux_linear_5__MUX_theta_state_inst_n232,
         all_mux_linear_5__MUX_theta_state_inst_n231,
         all_mux_linear_5__MUX_theta_state_inst_n230,
         all_mux_linear_6__MUX_theta_state_inst_n335,
         all_mux_linear_6__MUX_theta_state_inst_n334,
         all_mux_linear_6__MUX_theta_state_inst_n333,
         all_mux_linear_6__MUX_theta_state_inst_n332,
         all_mux_linear_6__MUX_theta_state_inst_n331,
         all_mux_linear_6__MUX_theta_state_inst_n330,
         all_mux_linear_6__MUX_theta_state_inst_n329,
         all_mux_linear_6__MUX_theta_state_inst_n328,
         all_mux_linear_6__MUX_theta_state_inst_n327,
         all_mux_linear_6__MUX_theta_state_inst_n326,
         all_mux_linear_6__MUX_theta_state_inst_n325,
         all_mux_linear_6__MUX_theta_state_inst_n324,
         all_mux_linear_6__MUX_theta_state_inst_n323,
         all_mux_linear_6__MUX_theta_state_inst_n322,
         all_mux_linear_6__MUX_theta_state_inst_n321,
         all_mux_linear_6__MUX_theta_state_inst_n320,
         all_mux_linear_6__MUX_theta_state_inst_n319,
         all_mux_linear_6__MUX_theta_state_inst_n318,
         all_mux_linear_6__MUX_theta_state_inst_n317,
         all_mux_linear_6__MUX_theta_state_inst_n316,
         all_mux_linear_6__MUX_theta_state_inst_n315,
         all_mux_linear_6__MUX_theta_state_inst_n314,
         all_mux_linear_6__MUX_theta_state_inst_n313,
         all_mux_linear_6__MUX_theta_state_inst_n312,
         all_mux_linear_6__MUX_theta_state_inst_n311,
         all_mux_linear_6__MUX_theta_state_inst_n310,
         all_mux_linear_6__MUX_theta_state_inst_n309,
         all_mux_linear_6__MUX_theta_state_inst_n308,
         all_mux_linear_6__MUX_theta_state_inst_n307,
         all_mux_linear_6__MUX_theta_state_inst_n306,
         all_mux_linear_6__MUX_theta_state_inst_n305,
         all_mux_linear_6__MUX_theta_state_inst_n304,
         all_mux_linear_6__MUX_theta_state_inst_n303,
         all_mux_linear_6__MUX_theta_state_inst_n302,
         all_mux_linear_6__MUX_theta_state_inst_n301,
         all_mux_linear_6__MUX_theta_state_inst_n300,
         all_mux_linear_6__MUX_theta_state_inst_n299,
         all_mux_linear_6__MUX_theta_state_inst_n298,
         all_mux_linear_6__MUX_theta_state_inst_n297,
         all_mux_linear_6__MUX_theta_state_inst_n296,
         all_mux_linear_6__MUX_theta_state_inst_n295,
         all_mux_linear_6__MUX_theta_state_inst_n294,
         all_mux_linear_6__MUX_theta_state_inst_n293,
         all_mux_linear_6__MUX_theta_state_inst_n292,
         all_mux_linear_6__MUX_theta_state_inst_n291,
         all_mux_linear_6__MUX_theta_state_inst_n290,
         all_mux_linear_6__MUX_theta_state_inst_n289,
         all_mux_linear_6__MUX_theta_state_inst_n288,
         all_mux_linear_6__MUX_theta_state_inst_n287,
         all_mux_linear_6__MUX_theta_state_inst_n286,
         all_mux_linear_6__MUX_theta_state_inst_n285,
         all_mux_linear_6__MUX_theta_state_inst_n284,
         all_mux_linear_6__MUX_theta_state_inst_n283,
         all_mux_linear_6__MUX_theta_state_inst_n282,
         all_mux_linear_6__MUX_theta_state_inst_n281,
         all_mux_linear_6__MUX_theta_state_inst_n280,
         all_mux_linear_6__MUX_theta_state_inst_n279,
         all_mux_linear_6__MUX_theta_state_inst_n278,
         all_mux_linear_6__MUX_theta_state_inst_n277,
         all_mux_linear_6__MUX_theta_state_inst_n276,
         all_mux_linear_6__MUX_theta_state_inst_n275,
         all_mux_linear_6__MUX_theta_state_inst_n274,
         all_mux_linear_6__MUX_theta_state_inst_n273,
         all_mux_linear_6__MUX_theta_state_inst_n272,
         all_mux_linear_6__MUX_theta_state_inst_n271,
         all_mux_linear_6__MUX_theta_state_inst_n270,
         all_mux_linear_6__MUX_theta_state_inst_n269,
         all_mux_linear_6__MUX_theta_state_inst_n268,
         all_mux_linear_6__MUX_theta_state_inst_n267,
         all_mux_linear_6__MUX_theta_state_inst_n266,
         all_mux_linear_6__MUX_theta_state_inst_n265,
         all_mux_linear_6__MUX_theta_state_inst_n264,
         all_mux_linear_6__MUX_theta_state_inst_n263,
         all_mux_linear_6__MUX_theta_state_inst_n262,
         all_mux_linear_6__MUX_theta_state_inst_n261,
         all_mux_linear_6__MUX_theta_state_inst_n260,
         all_mux_linear_6__MUX_theta_state_inst_n259,
         all_mux_linear_6__MUX_theta_state_inst_n258,
         all_mux_linear_6__MUX_theta_state_inst_n257,
         all_mux_linear_6__MUX_theta_state_inst_n256,
         all_mux_linear_6__MUX_theta_state_inst_n255,
         all_mux_linear_6__MUX_theta_state_inst_n254,
         all_mux_linear_6__MUX_theta_state_inst_n253,
         all_mux_linear_6__MUX_theta_state_inst_n252,
         all_mux_linear_6__MUX_theta_state_inst_n251,
         all_mux_linear_6__MUX_theta_state_inst_n250,
         all_mux_linear_6__MUX_theta_state_inst_n249,
         all_mux_linear_6__MUX_theta_state_inst_n248,
         all_mux_linear_6__MUX_theta_state_inst_n247,
         all_mux_linear_6__MUX_theta_state_inst_n246,
         all_mux_linear_6__MUX_theta_state_inst_n245,
         all_mux_linear_6__MUX_theta_state_inst_n244,
         all_mux_linear_6__MUX_theta_state_inst_n243,
         all_mux_linear_6__MUX_theta_state_inst_n242,
         all_mux_linear_6__MUX_theta_state_inst_n241,
         all_mux_linear_6__MUX_theta_state_inst_n240,
         all_mux_linear_6__MUX_theta_state_inst_n239,
         all_mux_linear_6__MUX_theta_state_inst_n238,
         all_mux_linear_6__MUX_theta_state_inst_n237,
         all_mux_linear_6__MUX_theta_state_inst_n236,
         all_mux_linear_6__MUX_theta_state_inst_n235,
         all_mux_linear_6__MUX_theta_state_inst_n234,
         all_mux_linear_6__MUX_theta_state_inst_n233,
         all_mux_linear_6__MUX_theta_state_inst_n232,
         all_mux_linear_6__MUX_theta_state_inst_n231,
         all_mux_linear_6__MUX_theta_state_inst_n230,
         all_mux_linear_6__MUX_theta_state_inst_n229,
         all_mux_linear_7__MUX_theta_state_inst_n336,
         all_mux_linear_7__MUX_theta_state_inst_n335,
         all_mux_linear_7__MUX_theta_state_inst_n334,
         all_mux_linear_7__MUX_theta_state_inst_n333,
         all_mux_linear_7__MUX_theta_state_inst_n332,
         all_mux_linear_7__MUX_theta_state_inst_n331,
         all_mux_linear_7__MUX_theta_state_inst_n330,
         all_mux_linear_7__MUX_theta_state_inst_n329,
         all_mux_linear_7__MUX_theta_state_inst_n328,
         all_mux_linear_7__MUX_theta_state_inst_n327,
         all_mux_linear_7__MUX_theta_state_inst_n326,
         all_mux_linear_7__MUX_theta_state_inst_n325,
         all_mux_linear_7__MUX_theta_state_inst_n324,
         all_mux_linear_7__MUX_theta_state_inst_n323,
         all_mux_linear_7__MUX_theta_state_inst_n322,
         all_mux_linear_7__MUX_theta_state_inst_n321,
         all_mux_linear_7__MUX_theta_state_inst_n320,
         all_mux_linear_7__MUX_theta_state_inst_n319,
         all_mux_linear_7__MUX_theta_state_inst_n318,
         all_mux_linear_7__MUX_theta_state_inst_n317,
         all_mux_linear_7__MUX_theta_state_inst_n316,
         all_mux_linear_7__MUX_theta_state_inst_n315,
         all_mux_linear_7__MUX_theta_state_inst_n314,
         all_mux_linear_7__MUX_theta_state_inst_n313,
         all_mux_linear_7__MUX_theta_state_inst_n312,
         all_mux_linear_7__MUX_theta_state_inst_n311,
         all_mux_linear_7__MUX_theta_state_inst_n310,
         all_mux_linear_7__MUX_theta_state_inst_n309,
         all_mux_linear_7__MUX_theta_state_inst_n308,
         all_mux_linear_7__MUX_theta_state_inst_n307,
         all_mux_linear_7__MUX_theta_state_inst_n306,
         all_mux_linear_7__MUX_theta_state_inst_n305,
         all_mux_linear_7__MUX_theta_state_inst_n304,
         all_mux_linear_7__MUX_theta_state_inst_n303,
         all_mux_linear_7__MUX_theta_state_inst_n302,
         all_mux_linear_7__MUX_theta_state_inst_n301,
         all_mux_linear_7__MUX_theta_state_inst_n300,
         all_mux_linear_7__MUX_theta_state_inst_n299,
         all_mux_linear_7__MUX_theta_state_inst_n298,
         all_mux_linear_7__MUX_theta_state_inst_n297,
         all_mux_linear_7__MUX_theta_state_inst_n296,
         all_mux_linear_7__MUX_theta_state_inst_n295,
         all_mux_linear_7__MUX_theta_state_inst_n294,
         all_mux_linear_7__MUX_theta_state_inst_n293,
         all_mux_linear_7__MUX_theta_state_inst_n292,
         all_mux_linear_7__MUX_theta_state_inst_n291,
         all_mux_linear_7__MUX_theta_state_inst_n290,
         all_mux_linear_7__MUX_theta_state_inst_n289,
         all_mux_linear_7__MUX_theta_state_inst_n288,
         all_mux_linear_7__MUX_theta_state_inst_n287,
         all_mux_linear_7__MUX_theta_state_inst_n286,
         all_mux_linear_7__MUX_theta_state_inst_n285,
         all_mux_linear_7__MUX_theta_state_inst_n284,
         all_mux_linear_7__MUX_theta_state_inst_n283,
         all_mux_linear_7__MUX_theta_state_inst_n282,
         all_mux_linear_7__MUX_theta_state_inst_n281,
         all_mux_linear_7__MUX_theta_state_inst_n280,
         all_mux_linear_7__MUX_theta_state_inst_n279,
         all_mux_linear_7__MUX_theta_state_inst_n278,
         all_mux_linear_7__MUX_theta_state_inst_n277,
         all_mux_linear_7__MUX_theta_state_inst_n276,
         all_mux_linear_7__MUX_theta_state_inst_n275,
         all_mux_linear_7__MUX_theta_state_inst_n274,
         all_mux_linear_7__MUX_theta_state_inst_n273,
         all_mux_linear_7__MUX_theta_state_inst_n272,
         all_mux_linear_7__MUX_theta_state_inst_n271,
         all_mux_linear_7__MUX_theta_state_inst_n270,
         all_mux_linear_7__MUX_theta_state_inst_n269,
         all_mux_linear_7__MUX_theta_state_inst_n268,
         all_mux_linear_7__MUX_theta_state_inst_n267,
         all_mux_linear_7__MUX_theta_state_inst_n266,
         all_mux_linear_7__MUX_theta_state_inst_n265,
         all_mux_linear_7__MUX_theta_state_inst_n264,
         all_mux_linear_7__MUX_theta_state_inst_n263,
         all_mux_linear_7__MUX_theta_state_inst_n262,
         all_mux_linear_7__MUX_theta_state_inst_n261,
         all_mux_linear_7__MUX_theta_state_inst_n260,
         all_mux_linear_7__MUX_theta_state_inst_n259,
         all_mux_linear_7__MUX_theta_state_inst_n258,
         all_mux_linear_7__MUX_theta_state_inst_n257,
         all_mux_linear_7__MUX_theta_state_inst_n256,
         all_mux_linear_7__MUX_theta_state_inst_n255,
         all_mux_linear_7__MUX_theta_state_inst_n254,
         all_mux_linear_7__MUX_theta_state_inst_n253,
         all_mux_linear_7__MUX_theta_state_inst_n252,
         all_mux_linear_7__MUX_theta_state_inst_n251,
         all_mux_linear_7__MUX_theta_state_inst_n250,
         all_mux_linear_7__MUX_theta_state_inst_n249,
         all_mux_linear_7__MUX_theta_state_inst_n248,
         all_mux_linear_7__MUX_theta_state_inst_n247,
         all_mux_linear_7__MUX_theta_state_inst_n246,
         all_mux_linear_7__MUX_theta_state_inst_n245,
         all_mux_linear_7__MUX_theta_state_inst_n244,
         all_mux_linear_7__MUX_theta_state_inst_n243,
         all_mux_linear_7__MUX_theta_state_inst_n242,
         all_mux_linear_7__MUX_theta_state_inst_n241,
         all_mux_linear_7__MUX_theta_state_inst_n240,
         all_mux_linear_7__MUX_theta_state_inst_n239,
         all_mux_linear_7__MUX_theta_state_inst_n238,
         all_mux_linear_7__MUX_theta_state_inst_n237,
         all_mux_linear_7__MUX_theta_state_inst_n236,
         all_mux_linear_7__MUX_theta_state_inst_n235,
         all_mux_linear_7__MUX_theta_state_inst_n234,
         all_mux_linear_7__MUX_theta_state_inst_n233,
         all_mux_linear_7__MUX_theta_state_inst_n232,
         all_mux_linear_7__MUX_theta_state_inst_n231,
         all_mux_linear_7__MUX_theta_state_inst_n230,
         all_mux_linear_8__MUX_theta_state_inst_n318,
         all_mux_linear_8__MUX_theta_state_inst_n317,
         all_mux_linear_8__MUX_theta_state_inst_n316,
         all_mux_linear_8__MUX_theta_state_inst_n315,
         all_mux_linear_8__MUX_theta_state_inst_n314,
         all_mux_linear_8__MUX_theta_state_inst_n313,
         all_mux_linear_8__MUX_theta_state_inst_n312,
         all_mux_linear_8__MUX_theta_state_inst_n311,
         all_mux_linear_8__MUX_theta_state_inst_n310,
         all_mux_linear_8__MUX_theta_state_inst_n309,
         all_mux_linear_8__MUX_theta_state_inst_n308,
         all_mux_linear_8__MUX_theta_state_inst_n307,
         all_mux_linear_8__MUX_theta_state_inst_n306,
         all_mux_linear_8__MUX_theta_state_inst_n305,
         all_mux_linear_8__MUX_theta_state_inst_n304,
         all_mux_linear_8__MUX_theta_state_inst_n303,
         all_mux_linear_8__MUX_theta_state_inst_n302,
         all_mux_linear_8__MUX_theta_state_inst_n301,
         all_mux_linear_8__MUX_theta_state_inst_n300,
         all_mux_linear_8__MUX_theta_state_inst_n299,
         all_mux_linear_8__MUX_theta_state_inst_n298,
         all_mux_linear_8__MUX_theta_state_inst_n297,
         all_mux_linear_8__MUX_theta_state_inst_n296,
         all_mux_linear_8__MUX_theta_state_inst_n295,
         all_mux_linear_8__MUX_theta_state_inst_n294,
         all_mux_linear_8__MUX_theta_state_inst_n293,
         all_mux_linear_8__MUX_theta_state_inst_n292,
         all_mux_linear_8__MUX_theta_state_inst_n291,
         all_mux_linear_8__MUX_theta_state_inst_n290,
         all_mux_linear_8__MUX_theta_state_inst_n289,
         all_mux_linear_8__MUX_theta_state_inst_n288,
         all_mux_linear_8__MUX_theta_state_inst_n287,
         all_mux_linear_8__MUX_theta_state_inst_n286,
         all_mux_linear_8__MUX_theta_state_inst_n285,
         all_mux_linear_8__MUX_theta_state_inst_n284,
         all_mux_linear_8__MUX_theta_state_inst_n283,
         all_mux_linear_8__MUX_theta_state_inst_n282,
         all_mux_linear_8__MUX_theta_state_inst_n281,
         all_mux_linear_8__MUX_theta_state_inst_n280,
         all_mux_linear_8__MUX_theta_state_inst_n279,
         all_mux_linear_8__MUX_theta_state_inst_n278,
         all_mux_linear_8__MUX_theta_state_inst_n277,
         all_mux_linear_8__MUX_theta_state_inst_n276,
         all_mux_linear_8__MUX_theta_state_inst_n275,
         all_mux_linear_8__MUX_theta_state_inst_n274,
         all_mux_linear_8__MUX_theta_state_inst_n273,
         all_mux_linear_8__MUX_theta_state_inst_n272,
         all_mux_linear_8__MUX_theta_state_inst_n271,
         all_mux_linear_8__MUX_theta_state_inst_n270,
         all_mux_linear_8__MUX_theta_state_inst_n269,
         all_mux_linear_8__MUX_theta_state_inst_n268,
         all_mux_linear_8__MUX_theta_state_inst_n267,
         all_mux_linear_8__MUX_theta_state_inst_n266,
         all_mux_linear_8__MUX_theta_state_inst_n265,
         all_mux_linear_8__MUX_theta_state_inst_n264,
         all_mux_linear_8__MUX_theta_state_inst_n263,
         all_mux_linear_8__MUX_theta_state_inst_n262,
         all_mux_linear_8__MUX_theta_state_inst_n261,
         all_mux_linear_8__MUX_theta_state_inst_n260,
         all_mux_linear_8__MUX_theta_state_inst_n259,
         all_mux_linear_8__MUX_theta_state_inst_n258,
         all_mux_linear_8__MUX_theta_state_inst_n257,
         all_mux_linear_8__MUX_theta_state_inst_n256,
         all_mux_linear_8__MUX_theta_state_inst_n255,
         all_mux_linear_8__MUX_theta_state_inst_n254,
         all_mux_linear_8__MUX_theta_state_inst_n253,
         all_mux_linear_8__MUX_theta_state_inst_n252,
         all_mux_linear_8__MUX_theta_state_inst_n251,
         all_mux_linear_8__MUX_theta_state_inst_n250,
         all_mux_linear_8__MUX_theta_state_inst_n249,
         all_mux_linear_8__MUX_theta_state_inst_n248,
         all_mux_linear_8__MUX_theta_state_inst_n247,
         all_mux_linear_8__MUX_theta_state_inst_n246,
         all_mux_linear_8__MUX_theta_state_inst_n245,
         all_mux_linear_8__MUX_theta_state_inst_n244,
         all_mux_linear_8__MUX_theta_state_inst_n243,
         all_mux_linear_8__MUX_theta_state_inst_n242,
         all_mux_linear_8__MUX_theta_state_inst_n241,
         all_mux_linear_8__MUX_theta_state_inst_n240,
         all_mux_linear_8__MUX_theta_state_inst_n239,
         all_mux_linear_8__MUX_theta_state_inst_n238,
         all_mux_linear_8__MUX_theta_state_inst_n237,
         all_mux_linear_8__MUX_theta_state_inst_n236,
         all_mux_linear_8__MUX_theta_state_inst_n235,
         all_mux_linear_8__MUX_theta_state_inst_n234,
         all_mux_linear_8__MUX_theta_state_inst_n233,
         all_mux_linear_8__MUX_theta_state_inst_n232,
         all_mux_linear_8__MUX_theta_state_inst_n231,
         all_mux_linear_8__MUX_theta_state_inst_n230,
         COMPRESSION_BITS_0__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_0__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_0__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_1__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_1__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_1__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_2__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_2__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_2__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_3__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_3__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_3__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_4__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_4__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_4__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_5__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_5__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_5__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_6__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_6__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_6__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_7__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_7__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_7__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_8__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_8__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_8__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_9__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_9__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_9__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_10__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_10__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_10__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_11__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_11__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_11__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_12__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_12__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_12__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_13__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_13__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_13__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_14__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_14__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_14__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_15__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_15__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_15__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_16__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_16__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_16__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_17__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_17__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_17__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_18__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_18__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_18__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_19__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_19__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_19__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_20__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_20__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_20__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_21__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_21__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_21__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_22__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_22__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_22__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_23__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_23__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_23__BIT_SHARES_2__Copression_n3,
         COMPRESSION_BITS_24__BIT_SHARES_0__Copression_n3,
         COMPRESSION_BITS_24__BIT_SHARES_1__Copression_n3,
         COMPRESSION_BITS_24__BIT_SHARES_2__Copression_n3, CHI_ChiOut_0_,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n2,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3,
         CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3,
         KECCAK_CONTROL_n62, KECCAK_CONTROL_n61, KECCAK_CONTROL_n60,
         KECCAK_CONTROL_n59, KECCAK_CONTROL_n58, KECCAK_CONTROL_n57,
         KECCAK_CONTROL_n56, KECCAK_CONTROL_n55, KECCAK_CONTROL_n54,
         KECCAK_CONTROL_n53, KECCAK_CONTROL_n52, KECCAK_CONTROL_n51,
         KECCAK_CONTROL_n50, KECCAK_CONTROL_n49, KECCAK_CONTROL_n48,
         KECCAK_CONTROL_n47, KECCAK_CONTROL_n46, KECCAK_CONTROL_n45,
         KECCAK_CONTROL_n44, KECCAK_CONTROL_n43, KECCAK_CONTROL_n42,
         KECCAK_CONTROL_n41, KECCAK_CONTROL_n40, KECCAK_CONTROL_n39,
         KECCAK_CONTROL_n38, KECCAK_CONTROL_n37, KECCAK_CONTROL_n36,
         KECCAK_CONTROL_n35, KECCAK_CONTROL_n34, KECCAK_CONTROL_n32,
         KECCAK_CONTROL_n31, KECCAK_CONTROL_n27, KECCAK_CONTROL_n26,
         KECCAK_CONTROL_n6, KECCAK_CONTROL_n29, KECCAK_CONTROL_n28,
         KECCAK_CONTROL_n15, KECCAK_CONTROL_n14, KECCAK_CONTROL_n5,
         KECCAK_CONTROL_N32, KECCAK_CONTROL_RoundCountxDP_0_,
         KECCAK_CONTROL_RoundCountxDP_1_, KECCAK_CONTROL_RoundCountxDP_2_,
         KECCAK_CONTROL_RoundCountxDP_3_, KECCAK_CONTROL_RoundCountxDP_4_,
         KECCAK_CONTROL_RC_GEN_n3, KECCAK_CONTROL_RC_GEN_n2;
  wire   [224:0] SlicesFromChi;
  wire   [224:0] StateOut;
  wire   [24:0] all_mux_linear_0__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_1__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_2__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_3__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_4__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_5__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_6__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_7__MUX_theta_state_inst_StateIn;
  wire   [24:0] all_mux_linear_8__MUX_theta_state_inst_StateIn;

  BUF_X1 U2 ( .A(Lastround), .Z(n4) );
  BUF_X1 U3 ( .A(Lastround), .Z(n2) );
  BUF_X1 U4 ( .A(Lastround), .Z(n3) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U116 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n218), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n217), .A(
        all_mux_linear_0__MUX_theta_state_inst_n216), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U115 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[9]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n218), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n215), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n216) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U114 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n214), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n217), .A(
        all_mux_linear_0__MUX_theta_state_inst_n213), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U113 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[8]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n214), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n215), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n213) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U112 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n212), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n217), .A(
        all_mux_linear_0__MUX_theta_state_inst_n211), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U111 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[7]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n212), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n215), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n211) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U110 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n210), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n217), .A(
        all_mux_linear_0__MUX_theta_state_inst_n209), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U109 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[6]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n210), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n215), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n209) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U108 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n208), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n217), .A(
        all_mux_linear_0__MUX_theta_state_inst_n207), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U107 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[5]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n208), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n215), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n207) );
  NOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U106 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n206), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n215) );
  NAND2_X1 all_mux_linear_0__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n131), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n206), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n217) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U104 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n205), .B(
        all_mux_linear_0__MUX_theta_state_inst_n204), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n206) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U103 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n203), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n202), .A(
        all_mux_linear_0__MUX_theta_state_inst_n201), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[4]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U102 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[4]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n200), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n203), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n201) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U101 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n199), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n202), .A(
        all_mux_linear_0__MUX_theta_state_inst_n198), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[3]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U100 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[3]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n200), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n199), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n198) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U99 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n197), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n202), .A(
        all_mux_linear_0__MUX_theta_state_inst_n196), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[2]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U98 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[2]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n200), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n197), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n196) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U97 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n195), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n194), .A(
        all_mux_linear_0__MUX_theta_state_inst_n193), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[24]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U96 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[24]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n195), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n192), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n193) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n191), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n194), .A(
        all_mux_linear_0__MUX_theta_state_inst_n190), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[23]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[23]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n191), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n192), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n190) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U93 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n189), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n194), .A(
        all_mux_linear_0__MUX_theta_state_inst_n188), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[22]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U92 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[22]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n189), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n192), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n188) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n187), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n194), .A(
        all_mux_linear_0__MUX_theta_state_inst_n186), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[21]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[21]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n187), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n192), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n186) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U89 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n185), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n194), .A(
        all_mux_linear_0__MUX_theta_state_inst_n184), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[20]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U88 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[20]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n185), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n192), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n184) );
  NOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U87 ( .A1(n3), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n183), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n192) );
  NAND2_X1 all_mux_linear_0__MUX_theta_state_inst_U86 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n131), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n183), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n194) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U85 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n182), .B(
        all_mux_linear_0__MUX_theta_state_inst_n204), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n183) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n181), .B(
        all_mux_linear_0__MUX_theta_state_inst_n180), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n204) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U83 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n179), .B(
        all_mux_linear_0__MUX_theta_state_inst_n178), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n180) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U82 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n177), .B(
        all_mux_linear_0__MUX_theta_state_inst_n203), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n178) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U81 ( .A1(Reset), .A2(
        InData[4]), .B1(SlicesFromChi[4]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n203) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U80 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n199), .B(
        all_mux_linear_0__MUX_theta_state_inst_n197), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n179) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U79 ( .A1(Reset), .A2(
        InData[2]), .B1(SlicesFromChi[2]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n197) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U78 ( .A1(Reset), .A2(
        InData[3]), .B1(SlicesFromChi[3]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n199) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n177), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n202), .A(
        all_mux_linear_0__MUX_theta_state_inst_n176), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[1]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[1]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n200), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n177), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n176) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U75 ( .A1(Reset), .A2(
        InData[1]), .B1(SlicesFromChi[1]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n177) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U74 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n175), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n174), .A(
        all_mux_linear_0__MUX_theta_state_inst_n173), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[19]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U73 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[19]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n175), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n172), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n173) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U72 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n171), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n174), .A(
        all_mux_linear_0__MUX_theta_state_inst_n170), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[18]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U71 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[18]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n171), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n172), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n170) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U70 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n169), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n174), .A(
        all_mux_linear_0__MUX_theta_state_inst_n168), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[17]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U69 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[17]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n169), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n172), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n168) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U68 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n167), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n174), .A(
        all_mux_linear_0__MUX_theta_state_inst_n166), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[16]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U67 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[16]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n167), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n172), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n166) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n165), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n174), .A(
        all_mux_linear_0__MUX_theta_state_inst_n164), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[15]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[15]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n165), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n172), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n164) );
  NOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U64 ( .A1(n3), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n163), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n172) );
  NAND2_X1 all_mux_linear_0__MUX_theta_state_inst_U63 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n131), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n163), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n174) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U62 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n162), .B(
        all_mux_linear_0__MUX_theta_state_inst_n205), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n163) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U61 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n161), .B(
        all_mux_linear_0__MUX_theta_state_inst_n160), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n205) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U60 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n159), .B(
        all_mux_linear_0__MUX_theta_state_inst_n158), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n160) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n157), .B(
        all_mux_linear_0__MUX_theta_state_inst_n156), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n158) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n155), .B(
        all_mux_linear_0__MUX_theta_state_inst_n154), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n159) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U57 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n155), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n153), .A(
        all_mux_linear_0__MUX_theta_state_inst_n152), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[14]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U56 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[14]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n151), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n155), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n152) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U55 ( .A1(Reset), .A2(
        InData[14]), .B1(SlicesFromChi[14]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n155) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n154), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n153), .A(
        all_mux_linear_0__MUX_theta_state_inst_n150), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[13]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[13]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n151), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n154), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n150) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U52 ( .A1(Reset), .A2(
        InData[13]), .B1(SlicesFromChi[13]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n154) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U51 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n156), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n153), .A(
        all_mux_linear_0__MUX_theta_state_inst_n149), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[12]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U50 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[12]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n151), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n156), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n149) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U49 ( .A1(Reset), .A2(
        InData[12]), .B1(SlicesFromChi[12]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n156) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U48 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n157), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n153), .A(
        all_mux_linear_0__MUX_theta_state_inst_n148), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[11]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U47 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[11]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n151), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n157), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n148) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U46 ( .A1(Reset), .A2(
        InData[11]), .B1(SlicesFromChi[11]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n157) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U45 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n161), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n153), .A(
        all_mux_linear_0__MUX_theta_state_inst_n147), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[10]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U44 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n130), .A2(SlicesFromChi[10]), 
        .B1(all_mux_linear_0__MUX_theta_state_inst_n161), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n151), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n147) );
  NOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U43 ( .A1(n3), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n146), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n151) );
  NAND2_X1 all_mux_linear_0__MUX_theta_state_inst_U42 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n131), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n146), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n153) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U41 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n145), .B(
        all_mux_linear_0__MUX_theta_state_inst_n182), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n146) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U40 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n175), .B(
        all_mux_linear_0__MUX_theta_state_inst_n144), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n182) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U39 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n143), .B(
        all_mux_linear_0__MUX_theta_state_inst_n142), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n144) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U38 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n167), .B(
        all_mux_linear_0__MUX_theta_state_inst_n165), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n142) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U37 ( .A1(Reset), .A2(
        InData[15]), .B1(SlicesFromChi[15]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n165) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U36 ( .A1(Reset), .A2(
        InData[16]), .B1(SlicesFromChi[16]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n167) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n171), .B(
        all_mux_linear_0__MUX_theta_state_inst_n169), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n143) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U34 ( .A1(Reset), .A2(
        InData[17]), .B1(SlicesFromChi[17]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n169) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U33 ( .A1(Reset), .A2(
        InData[18]), .B1(SlicesFromChi[18]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n171) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U32 ( .A1(Reset), .A2(
        InData[19]), .B1(SlicesFromChi[19]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n132), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n175) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U31 ( .A1(Reset), .A2(
        InData[10]), .B1(SlicesFromChi[10]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n161) );
  OAI21_X1 all_mux_linear_0__MUX_theta_state_inst_U30 ( .B1(
        all_mux_linear_0__MUX_theta_state_inst_n181), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n202), .A(
        all_mux_linear_0__MUX_theta_state_inst_n141), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[0]) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[0]), 
        .A2(all_mux_linear_0__MUX_theta_state_inst_n130), .B1(
        all_mux_linear_0__MUX_theta_state_inst_n181), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n200), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n141) );
  NOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U28 ( .A1(n3), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n140), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n200) );
  NAND2_X1 all_mux_linear_0__MUX_theta_state_inst_U27 ( .A1(
        all_mux_linear_0__MUX_theta_state_inst_n131), .A2(
        all_mux_linear_0__MUX_theta_state_inst_n140), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n202) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U26 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n162), .B(
        all_mux_linear_0__MUX_theta_state_inst_n145), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n140) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U25 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n212), .B(
        all_mux_linear_0__MUX_theta_state_inst_n139), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n145) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n138), .B(
        all_mux_linear_0__MUX_theta_state_inst_n137), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n139) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U23 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n210), .B(
        all_mux_linear_0__MUX_theta_state_inst_n208), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n137) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U22 ( .A1(Reset), .A2(
        InData[5]), .B1(SlicesFromChi[5]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n208) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U21 ( .A1(Reset), .A2(
        InData[6]), .B1(SlicesFromChi[6]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n210) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U20 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n214), .B(
        all_mux_linear_0__MUX_theta_state_inst_n218), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n138) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U19 ( .A1(Reset), .A2(
        InData[9]), .B1(SlicesFromChi[9]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n218) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U18 ( .A1(Reset), .A2(
        InData[8]), .B1(SlicesFromChi[8]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n214) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U17 ( .A1(Reset), .A2(
        InData[7]), .B1(SlicesFromChi[7]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n212) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U16 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n195), .B(
        all_mux_linear_0__MUX_theta_state_inst_n136), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n162) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U15 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n135), .B(
        all_mux_linear_0__MUX_theta_state_inst_n134), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n136) );
  XNOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U14 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n187), .B(
        all_mux_linear_0__MUX_theta_state_inst_n185), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n134) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U13 ( .A1(Reset), .A2(
        InData[20]), .B1(SlicesFromChi[20]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n185) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U12 ( .A1(Reset), .A2(
        InData[21]), .B1(SlicesFromChi[21]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n187) );
  XOR2_X1 all_mux_linear_0__MUX_theta_state_inst_U11 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n191), .B(
        all_mux_linear_0__MUX_theta_state_inst_n189), .Z(
        all_mux_linear_0__MUX_theta_state_inst_n135) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U10 ( .A1(Reset), .A2(
        InData[22]), .B1(SlicesFromChi[22]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n189) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U9 ( .A1(Reset), .A2(
        InData[23]), .B1(SlicesFromChi[23]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n191) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U8 ( .A1(Reset), .A2(
        InData[24]), .B1(SlicesFromChi[24]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n195) );
  AOI22_X1 all_mux_linear_0__MUX_theta_state_inst_U7 ( .A1(Reset), .A2(
        InData[0]), .B1(SlicesFromChi[0]), .B2(
        all_mux_linear_0__MUX_theta_state_inst_n133), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n181) );
  INV_X2 all_mux_linear_0__MUX_theta_state_inst_U6 ( .A(
        all_mux_linear_0__MUX_theta_state_inst_n131), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n130) );
  INV_X1 all_mux_linear_0__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n133) );
  INV_X1 all_mux_linear_0__MUX_theta_state_inst_U4 ( .A(Reset), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n132) );
  INV_X1 all_mux_linear_0__MUX_theta_state_inst_U3 ( .A(n3), .ZN(
        all_mux_linear_0__MUX_theta_state_inst_n131) );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[9]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[5]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[6]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[7]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[8]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[0]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[1]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[2]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[3]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[4]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[10]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[11]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[12]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[13]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[14]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[15]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[16]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[17]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[18]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[19]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[20]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[21]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[22]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[23]), .QN() );
  DFF_X1 all_mux_linear_0__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_0__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[24]), .QN() );
  OAI21_X1 all_mux_linear_1__MUX_theta_state_inst_U134 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n335), .A(
        all_mux_linear_1__MUX_theta_state_inst_n334), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_1__MUX_theta_state_inst_U133 ( .A1(n2), .A2(
        SlicesFromChi[34]), .B1(all_mux_linear_1__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_1__MUX_theta_state_inst_n335), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n334) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U132 ( .A1(SlicesFromChi[34]), .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n335) );
  OAI21_X1 all_mux_linear_1__MUX_theta_state_inst_U131 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n332), .A(
        all_mux_linear_1__MUX_theta_state_inst_n331), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_1__MUX_theta_state_inst_U130 ( .A1(n2), .A2(
        SlicesFromChi[33]), .B1(all_mux_linear_1__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_1__MUX_theta_state_inst_n332), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n331) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U129 ( .A1(SlicesFromChi[33]), .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n332) );
  OAI21_X1 all_mux_linear_1__MUX_theta_state_inst_U128 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n330), .A(
        all_mux_linear_1__MUX_theta_state_inst_n329), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_1__MUX_theta_state_inst_U127 ( .A1(n2), .A2(
        SlicesFromChi[32]), .B1(all_mux_linear_1__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_1__MUX_theta_state_inst_n330), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n329) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U126 ( .A1(SlicesFromChi[32]), .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n330) );
  OAI21_X1 all_mux_linear_1__MUX_theta_state_inst_U125 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n328), .A(
        all_mux_linear_1__MUX_theta_state_inst_n327), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_1__MUX_theta_state_inst_U124 ( .A1(n2), .A2(
        SlicesFromChi[31]), .B1(all_mux_linear_1__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_1__MUX_theta_state_inst_n328), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n327) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U123 ( .A1(SlicesFromChi[31]), .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n328) );
  OAI21_X1 all_mux_linear_1__MUX_theta_state_inst_U122 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n326), .A(
        all_mux_linear_1__MUX_theta_state_inst_n325), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_1__MUX_theta_state_inst_U121 ( .A1(n2), .A2(
        SlicesFromChi[30]), .B1(all_mux_linear_1__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_1__MUX_theta_state_inst_n326), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n325) );
  AND2_X1 all_mux_linear_1__MUX_theta_state_inst_U120 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n336), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n333) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U119 ( .A1(SlicesFromChi[30]), .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n326) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U118 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n324), .B(
        all_mux_linear_1__MUX_theta_state_inst_n323), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n336) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U117 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n322), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n320), .A(
        all_mux_linear_1__MUX_theta_state_inst_n319), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[4]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U116 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n322), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n319) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U115 ( .A(SlicesFromChi[29]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n320) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U114 ( .A1(SlicesFromChi[29]), .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n322) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U113 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n318), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n317), .A(
        all_mux_linear_1__MUX_theta_state_inst_n316), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[3]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U112 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n318), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n316) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U111 ( .A(SlicesFromChi[28]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n317) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U110 ( .A1(SlicesFromChi[28]), .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n318) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U109 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n315), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n314), .A(
        all_mux_linear_1__MUX_theta_state_inst_n313), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[2]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U108 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n315), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n313) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U107 ( .A1(SlicesFromChi[27]), .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n315) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U106 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n312), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n310), .A(
        all_mux_linear_1__MUX_theta_state_inst_n309), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[24]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n312), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n309) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U104 ( .A(SlicesFromChi[49]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n310) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U103 ( .A1(SlicesFromChi[49]), .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n312) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U102 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n308), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n307), .A(
        all_mux_linear_1__MUX_theta_state_inst_n306), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[23]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U101 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n308), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n306) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U100 ( .A(SlicesFromChi[48]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n307) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U99 ( .A1(SlicesFromChi[48]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n308) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U98 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n305), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n304), .A(
        all_mux_linear_1__MUX_theta_state_inst_n303), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[22]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U97 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n305), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n303) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U96 ( .A1(SlicesFromChi[47]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n305) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n302), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n301), .A(
        all_mux_linear_1__MUX_theta_state_inst_n300), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[21]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n302), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n300) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U93 ( .A(SlicesFromChi[46]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n301) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U92 ( .A1(SlicesFromChi[46]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n302) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n299), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n298), .A(
        all_mux_linear_1__MUX_theta_state_inst_n297), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[20]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n299), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n297) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U89 ( .A(SlicesFromChi[45]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n298) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U88 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n295), .B(
        all_mux_linear_1__MUX_theta_state_inst_n294), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n324) );
  XOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U87 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n293), .B(
        all_mux_linear_1__MUX_theta_state_inst_n292), .Z(
        all_mux_linear_1__MUX_theta_state_inst_n294) );
  OAI211_X1 all_mux_linear_1__MUX_theta_state_inst_U86 ( .C1(SlicesFromChi[29]), .C2(all_mux_linear_1__MUX_theta_state_inst_n291), .A(
        all_mux_linear_1__MUX_theta_state_inst_n233), .B(
        all_mux_linear_1__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n295) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U85 ( .A1(SlicesFromChi[29]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n291), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n290) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n314), .B(SlicesFromChi[28]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n291) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U83 ( .A(SlicesFromChi[27]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n314) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U82 ( .A1(SlicesFromChi[45]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n299) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U81 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n292), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n289), .A(
        all_mux_linear_1__MUX_theta_state_inst_n288), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[1]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U80 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n292), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n288) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U79 ( .A(SlicesFromChi[26]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n289) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U78 ( .A1(SlicesFromChi[26]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n292) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n287), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n285), .A(
        all_mux_linear_1__MUX_theta_state_inst_n284), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[19]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n287), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n284) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U75 ( .A(SlicesFromChi[44]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n285) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U74 ( .A1(SlicesFromChi[44]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n287) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U73 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n283), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n282), .A(
        all_mux_linear_1__MUX_theta_state_inst_n281), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[18]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U72 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n283), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n281) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U71 ( .A(SlicesFromChi[43]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n282) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U70 ( .A1(SlicesFromChi[43]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n283) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U69 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n280), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n279), .A(
        all_mux_linear_1__MUX_theta_state_inst_n278), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[17]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U68 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n280), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n278) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U67 ( .A1(SlicesFromChi[42]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n280) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n277), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n276), .A(
        all_mux_linear_1__MUX_theta_state_inst_n275), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[16]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n277), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n275) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U64 ( .A(SlicesFromChi[41]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n276) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U63 ( .A1(SlicesFromChi[41]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n277) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U62 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n274), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n273), .A(
        all_mux_linear_1__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[15]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U61 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n274), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n272) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U60 ( .A(SlicesFromChi[40]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n273) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n270), .B(
        all_mux_linear_1__MUX_theta_state_inst_n269), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n323) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n268), .B(
        all_mux_linear_1__MUX_theta_state_inst_n267), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n269) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U57 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n266), .B(
        all_mux_linear_1__MUX_theta_state_inst_n265), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n268) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U56 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n264), .B(
        all_mux_linear_1__MUX_theta_state_inst_n263), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n270) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U55 ( .A1(SlicesFromChi[40]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n274) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n267), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n261), .A(
        all_mux_linear_1__MUX_theta_state_inst_n260), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[14]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n267), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n260) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U52 ( .A(SlicesFromChi[39]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n261) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U51 ( .A1(SlicesFromChi[39]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n267) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U50 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n259), .A(
        all_mux_linear_1__MUX_theta_state_inst_n258), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[13]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U49 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n265), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n258) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U48 ( .A(SlicesFromChi[38]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n259) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U47 ( .A1(SlicesFromChi[38]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n265) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U46 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n266), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n257), .A(
        all_mux_linear_1__MUX_theta_state_inst_n256), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[12]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U45 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n266), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n256) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U44 ( .A(SlicesFromChi[37]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n257) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U43 ( .A1(SlicesFromChi[37]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n266) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U42 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n263), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n255), .A(
        all_mux_linear_1__MUX_theta_state_inst_n254), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[11]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U41 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n263), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n254) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U40 ( .A(SlicesFromChi[36]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n255) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U39 ( .A1(SlicesFromChi[36]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n263) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U38 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n264), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n253), .A(
        all_mux_linear_1__MUX_theta_state_inst_n252), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[10]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U37 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n264), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n252) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U36 ( .A(SlicesFromChi[35]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n253) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n250), .B(
        all_mux_linear_1__MUX_theta_state_inst_n249), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n296) );
  OAI211_X1 all_mux_linear_1__MUX_theta_state_inst_U34 ( .C1(SlicesFromChi[40]), .C2(all_mux_linear_1__MUX_theta_state_inst_n248), .A(
        all_mux_linear_1__MUX_theta_state_inst_n233), .B(
        all_mux_linear_1__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n249) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U33 ( .A1(SlicesFromChi[40]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n247) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U32 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n279), .B(SlicesFromChi[43]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n248) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U31 ( .A(SlicesFromChi[42]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n279) );
  OAI211_X1 all_mux_linear_1__MUX_theta_state_inst_U30 ( .C1(SlicesFromChi[41]), .C2(SlicesFromChi[44]), .A(all_mux_linear_1__MUX_theta_state_inst_n232), .B(
        all_mux_linear_1__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n250) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[44]), 
        .A2(SlicesFromChi[41]), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n246) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U28 ( .A1(SlicesFromChi[35]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n264) );
  OAI221_X1 all_mux_linear_1__MUX_theta_state_inst_U27 ( .B1(
        all_mux_linear_1__MUX_theta_state_inst_n293), .B2(
        all_mux_linear_1__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_1__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_1__MUX_theta_state_inst_n245), .A(
        all_mux_linear_1__MUX_theta_state_inst_n244), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[0]) );
  NAND3_X1 all_mux_linear_1__MUX_theta_state_inst_U26 ( .A1(
        all_mux_linear_1__MUX_theta_state_inst_n293), .A2(
        all_mux_linear_1__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_1__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n244) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U25 ( .A(SlicesFromChi[25]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n245) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n243), .B(
        all_mux_linear_1__MUX_theta_state_inst_n242), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n251) );
  AOI211_X1 all_mux_linear_1__MUX_theta_state_inst_U23 ( .C1(SlicesFromChi[31]), .C2(SlicesFromChi[32]), .A(Reset), .B(
        all_mux_linear_1__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n242) );
  NOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U22 ( .A1(SlicesFromChi[31]), 
        .A2(SlicesFromChi[32]), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n241) );
  OAI211_X1 all_mux_linear_1__MUX_theta_state_inst_U21 ( .C1(SlicesFromChi[30]), .C2(all_mux_linear_1__MUX_theta_state_inst_n240), .A(
        all_mux_linear_1__MUX_theta_state_inst_n232), .B(
        all_mux_linear_1__MUX_theta_state_inst_n239), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n243) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U20 ( .A1(SlicesFromChi[30]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n239) );
  XOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U19 ( .A(SlicesFromChi[34]), 
        .B(SlicesFromChi[33]), .Z(all_mux_linear_1__MUX_theta_state_inst_n240)
         );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U18 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n238), .B(
        all_mux_linear_1__MUX_theta_state_inst_n237), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n271) );
  AOI211_X1 all_mux_linear_1__MUX_theta_state_inst_U17 ( .C1(SlicesFromChi[46]), .C2(SlicesFromChi[49]), .A(Reset), .B(
        all_mux_linear_1__MUX_theta_state_inst_n236), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n237) );
  NOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U16 ( .A1(SlicesFromChi[46]), 
        .A2(SlicesFromChi[49]), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n236) );
  OAI211_X1 all_mux_linear_1__MUX_theta_state_inst_U15 ( .C1(SlicesFromChi[45]), .C2(all_mux_linear_1__MUX_theta_state_inst_n235), .A(
        all_mux_linear_1__MUX_theta_state_inst_n232), .B(
        all_mux_linear_1__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n238) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U14 ( .A1(SlicesFromChi[45]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n235), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n234) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U13 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n304), .B(SlicesFromChi[48]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n235) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U12 ( .A(SlicesFromChi[47]), 
        .ZN(all_mux_linear_1__MUX_theta_state_inst_n304) );
  NAND2_X1 all_mux_linear_1__MUX_theta_state_inst_U11 ( .A1(SlicesFromChi[25]), 
        .A2(all_mux_linear_1__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n293) );
  XOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U10 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n271), .B(
        all_mux_linear_1__MUX_theta_state_inst_n251), .Z(
        all_mux_linear_1__MUX_theta_state_inst_n321) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U9 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n271), .B(
        all_mux_linear_1__MUX_theta_state_inst_n323), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n286) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U8 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n324), .B(
        all_mux_linear_1__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n311) );
  XNOR2_X1 all_mux_linear_1__MUX_theta_state_inst_U7 ( .A(
        all_mux_linear_1__MUX_theta_state_inst_n251), .B(
        all_mux_linear_1__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n262) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U6 ( .A(Reset), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n233) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U4 ( .A(n2), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n231) );
  INV_X1 all_mux_linear_1__MUX_theta_state_inst_U3 ( .A(n2), .ZN(
        all_mux_linear_1__MUX_theta_state_inst_n230) );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[25]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[26]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[27]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[28]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[29]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[30]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[31]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[32]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[33]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[34]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[35]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[36]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[37]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[38]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[39]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[40]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[41]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[42]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[43]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[44]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[45]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[46]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[47]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[48]), .QN() );
  DFF_X1 all_mux_linear_1__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_1__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[49]), .QN() );
  OAI21_X1 all_mux_linear_2__MUX_theta_state_inst_U134 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n334), .A(
        all_mux_linear_2__MUX_theta_state_inst_n333), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_2__MUX_theta_state_inst_U133 ( .A1(n3), .A2(
        SlicesFromChi[59]), .B1(all_mux_linear_2__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_2__MUX_theta_state_inst_n334), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n333) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U132 ( .A1(SlicesFromChi[59]), .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n334) );
  OAI21_X1 all_mux_linear_2__MUX_theta_state_inst_U131 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n331), .A(
        all_mux_linear_2__MUX_theta_state_inst_n330), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_2__MUX_theta_state_inst_U130 ( .A1(n3), .A2(
        SlicesFromChi[58]), .B1(all_mux_linear_2__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_2__MUX_theta_state_inst_n331), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n330) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U129 ( .A1(SlicesFromChi[58]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n331) );
  OAI21_X1 all_mux_linear_2__MUX_theta_state_inst_U128 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n329), .A(
        all_mux_linear_2__MUX_theta_state_inst_n328), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_2__MUX_theta_state_inst_U127 ( .A1(n3), .A2(
        SlicesFromChi[57]), .B1(all_mux_linear_2__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_2__MUX_theta_state_inst_n329), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n328) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U126 ( .A1(SlicesFromChi[57]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n329) );
  OAI21_X1 all_mux_linear_2__MUX_theta_state_inst_U125 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n327), .A(
        all_mux_linear_2__MUX_theta_state_inst_n326), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_2__MUX_theta_state_inst_U124 ( .A1(n3), .A2(
        SlicesFromChi[56]), .B1(all_mux_linear_2__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_2__MUX_theta_state_inst_n327), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n326) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U123 ( .A1(SlicesFromChi[56]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n327) );
  OAI21_X1 all_mux_linear_2__MUX_theta_state_inst_U122 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n325), .A(
        all_mux_linear_2__MUX_theta_state_inst_n324), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_2__MUX_theta_state_inst_U121 ( .A1(n3), .A2(
        SlicesFromChi[55]), .B1(all_mux_linear_2__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_2__MUX_theta_state_inst_n325), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n324) );
  AND2_X1 all_mux_linear_2__MUX_theta_state_inst_U120 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n335), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n332) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U119 ( .A1(SlicesFromChi[55]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n325) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U118 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n323), .B(
        all_mux_linear_2__MUX_theta_state_inst_n322), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n335) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U117 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n321), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n319), .A(
        all_mux_linear_2__MUX_theta_state_inst_n318), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[4]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U116 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n321), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n318) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U115 ( .A(SlicesFromChi[54]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n319) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U114 ( .A1(SlicesFromChi[54]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n321) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U113 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n317), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n316), .A(
        all_mux_linear_2__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[3]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U112 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n317), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n315) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U111 ( .A(SlicesFromChi[53]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n316) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U110 ( .A1(SlicesFromChi[53]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n317) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U109 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n313), .A(
        all_mux_linear_2__MUX_theta_state_inst_n312), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[2]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U108 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n314), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n312) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U107 ( .A1(SlicesFromChi[52]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n314) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U106 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n311), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n309), .A(
        all_mux_linear_2__MUX_theta_state_inst_n308), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[24]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n311), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n308) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U104 ( .A(SlicesFromChi[74]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n309) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U103 ( .A1(SlicesFromChi[74]), .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n311) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U102 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n307), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n306), .A(
        all_mux_linear_2__MUX_theta_state_inst_n305), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[23]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U101 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n307), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n305) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U100 ( .A(SlicesFromChi[73]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n306) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U99 ( .A1(SlicesFromChi[73]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n307) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U98 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n304), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n303), .A(
        all_mux_linear_2__MUX_theta_state_inst_n302), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[22]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U97 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n304), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n302) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U96 ( .A1(SlicesFromChi[72]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n304) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n301), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n300), .A(
        all_mux_linear_2__MUX_theta_state_inst_n299), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[21]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n301), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n299) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U93 ( .A(SlicesFromChi[71]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n300) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U92 ( .A1(SlicesFromChi[71]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n301) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n298), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n297), .A(
        all_mux_linear_2__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[20]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n298), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n296) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U89 ( .A(SlicesFromChi[70]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n297) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U88 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n294), .B(
        all_mux_linear_2__MUX_theta_state_inst_n293), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n323) );
  XOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U87 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n292), .B(
        all_mux_linear_2__MUX_theta_state_inst_n291), .Z(
        all_mux_linear_2__MUX_theta_state_inst_n293) );
  OAI211_X1 all_mux_linear_2__MUX_theta_state_inst_U86 ( .C1(SlicesFromChi[54]), .C2(all_mux_linear_2__MUX_theta_state_inst_n290), .A(
        all_mux_linear_2__MUX_theta_state_inst_n232), .B(
        all_mux_linear_2__MUX_theta_state_inst_n289), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n294) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U85 ( .A1(SlicesFromChi[54]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n289) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n313), .B(SlicesFromChi[53]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n290) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U83 ( .A(SlicesFromChi[52]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n313) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U82 ( .A1(SlicesFromChi[70]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n298) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U81 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n288), .A(
        all_mux_linear_2__MUX_theta_state_inst_n287), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[1]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U80 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n291), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n287) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U79 ( .A(SlicesFromChi[51]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n288) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U78 ( .A1(SlicesFromChi[51]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n291) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n286), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n284), .A(
        all_mux_linear_2__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[19]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n286), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n283) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U75 ( .A(SlicesFromChi[69]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n284) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U74 ( .A1(SlicesFromChi[69]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n286) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U73 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n282), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n281), .A(
        all_mux_linear_2__MUX_theta_state_inst_n280), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[18]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U72 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n282), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n280) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U71 ( .A(SlicesFromChi[68]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n281) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U70 ( .A1(SlicesFromChi[68]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n282) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U69 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n279), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n278), .A(
        all_mux_linear_2__MUX_theta_state_inst_n277), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[17]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U68 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n279), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n277) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U67 ( .A1(SlicesFromChi[67]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n279) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n276), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n275), .A(
        all_mux_linear_2__MUX_theta_state_inst_n274), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[16]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n276), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n274) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U64 ( .A(SlicesFromChi[66]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n275) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U63 ( .A1(SlicesFromChi[66]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n276) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U62 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n273), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n272), .A(
        all_mux_linear_2__MUX_theta_state_inst_n271), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[15]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U61 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n273), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n271) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U60 ( .A(SlicesFromChi[65]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n272) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n269), .B(
        all_mux_linear_2__MUX_theta_state_inst_n268), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n322) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n267), .B(
        all_mux_linear_2__MUX_theta_state_inst_n266), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n268) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U57 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n265), .B(
        all_mux_linear_2__MUX_theta_state_inst_n264), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n267) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U56 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n263), .B(
        all_mux_linear_2__MUX_theta_state_inst_n262), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n269) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U55 ( .A1(SlicesFromChi[65]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n273) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n266), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n260), .A(
        all_mux_linear_2__MUX_theta_state_inst_n259), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[14]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n266), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n259) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U52 ( .A(SlicesFromChi[64]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n260) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U51 ( .A1(SlicesFromChi[64]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n266) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U50 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n264), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n258), .A(
        all_mux_linear_2__MUX_theta_state_inst_n257), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[13]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U49 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n264), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n257) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U48 ( .A(SlicesFromChi[63]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n258) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U47 ( .A1(SlicesFromChi[63]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n264) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U46 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n256), .A(
        all_mux_linear_2__MUX_theta_state_inst_n255), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[12]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U45 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n265), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n255) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U44 ( .A(SlicesFromChi[62]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n256) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U43 ( .A1(SlicesFromChi[62]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n265) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U42 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n262), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n254), .A(
        all_mux_linear_2__MUX_theta_state_inst_n253), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[11]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U41 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n262), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n253) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U40 ( .A(SlicesFromChi[61]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n254) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U39 ( .A1(SlicesFromChi[61]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n262) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U38 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n263), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n252), .A(
        all_mux_linear_2__MUX_theta_state_inst_n251), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[10]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U37 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n263), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n251) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U36 ( .A(SlicesFromChi[60]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n252) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n249), .B(
        all_mux_linear_2__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n295) );
  OAI211_X1 all_mux_linear_2__MUX_theta_state_inst_U34 ( .C1(SlicesFromChi[65]), .C2(all_mux_linear_2__MUX_theta_state_inst_n247), .A(
        all_mux_linear_2__MUX_theta_state_inst_n232), .B(
        all_mux_linear_2__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n248) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U33 ( .A1(SlicesFromChi[65]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n246) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U32 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n278), .B(SlicesFromChi[68]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n247) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U31 ( .A(SlicesFromChi[67]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n278) );
  OAI211_X1 all_mux_linear_2__MUX_theta_state_inst_U30 ( .C1(SlicesFromChi[66]), .C2(SlicesFromChi[69]), .A(all_mux_linear_2__MUX_theta_state_inst_n231), .B(
        all_mux_linear_2__MUX_theta_state_inst_n245), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n249) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[69]), 
        .A2(SlicesFromChi[66]), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n245) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U28 ( .A1(SlicesFromChi[60]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n263) );
  OAI221_X1 all_mux_linear_2__MUX_theta_state_inst_U27 ( .B1(
        all_mux_linear_2__MUX_theta_state_inst_n292), .B2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_2__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_2__MUX_theta_state_inst_n244), .A(
        all_mux_linear_2__MUX_theta_state_inst_n243), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[0]) );
  NAND3_X1 all_mux_linear_2__MUX_theta_state_inst_U26 ( .A1(
        all_mux_linear_2__MUX_theta_state_inst_n292), .A2(
        all_mux_linear_2__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_2__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n243) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U25 ( .A(SlicesFromChi[50]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n244) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n242), .B(
        all_mux_linear_2__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n250) );
  AOI211_X1 all_mux_linear_2__MUX_theta_state_inst_U23 ( .C1(SlicesFromChi[56]), .C2(SlicesFromChi[57]), .A(Reset), .B(
        all_mux_linear_2__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n241) );
  NOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U22 ( .A1(SlicesFromChi[56]), 
        .A2(SlicesFromChi[57]), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n240) );
  OAI211_X1 all_mux_linear_2__MUX_theta_state_inst_U21 ( .C1(SlicesFromChi[55]), .C2(all_mux_linear_2__MUX_theta_state_inst_n239), .A(
        all_mux_linear_2__MUX_theta_state_inst_n231), .B(
        all_mux_linear_2__MUX_theta_state_inst_n238), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n242) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U20 ( .A1(SlicesFromChi[55]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n239), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n238) );
  XOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U19 ( .A(SlicesFromChi[59]), 
        .B(SlicesFromChi[58]), .Z(all_mux_linear_2__MUX_theta_state_inst_n239)
         );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U18 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n237), .B(
        all_mux_linear_2__MUX_theta_state_inst_n236), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n270) );
  AOI211_X1 all_mux_linear_2__MUX_theta_state_inst_U17 ( .C1(SlicesFromChi[71]), .C2(SlicesFromChi[74]), .A(Reset), .B(
        all_mux_linear_2__MUX_theta_state_inst_n235), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n236) );
  NOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U16 ( .A1(SlicesFromChi[71]), 
        .A2(SlicesFromChi[74]), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n235) );
  OAI211_X1 all_mux_linear_2__MUX_theta_state_inst_U15 ( .C1(SlicesFromChi[70]), .C2(all_mux_linear_2__MUX_theta_state_inst_n234), .A(
        all_mux_linear_2__MUX_theta_state_inst_n231), .B(
        all_mux_linear_2__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n237) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U14 ( .A1(SlicesFromChi[70]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n233) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U13 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n303), .B(SlicesFromChi[73]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n234) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U12 ( .A(SlicesFromChi[72]), 
        .ZN(all_mux_linear_2__MUX_theta_state_inst_n303) );
  NAND2_X1 all_mux_linear_2__MUX_theta_state_inst_U11 ( .A1(SlicesFromChi[50]), 
        .A2(all_mux_linear_2__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n292) );
  XOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U10 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n270), .B(
        all_mux_linear_2__MUX_theta_state_inst_n250), .Z(
        all_mux_linear_2__MUX_theta_state_inst_n320) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U9 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n270), .B(
        all_mux_linear_2__MUX_theta_state_inst_n322), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n285) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U8 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n323), .B(
        all_mux_linear_2__MUX_theta_state_inst_n295), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n310) );
  XNOR2_X1 all_mux_linear_2__MUX_theta_state_inst_U7 ( .A(
        all_mux_linear_2__MUX_theta_state_inst_n250), .B(
        all_mux_linear_2__MUX_theta_state_inst_n295), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n261) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U6 ( .A(Reset), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n231) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U4 ( .A(n3), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n230) );
  INV_X1 all_mux_linear_2__MUX_theta_state_inst_U3 ( .A(n3), .ZN(
        all_mux_linear_2__MUX_theta_state_inst_n229) );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[50]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[51]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[52]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[53]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[54]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[55]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[56]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[57]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[58]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[59]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[60]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[61]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[62]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[63]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[64]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[65]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[66]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[67]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[68]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[69]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[70]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[71]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[72]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[73]), .QN() );
  DFF_X1 all_mux_linear_2__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_2__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[74]), .QN() );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U134 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n334), .A(
        all_mux_linear_3__MUX_theta_state_inst_n333), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U133 ( .A1(n2), .A2(
        SlicesFromChi[84]), .B1(all_mux_linear_3__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_3__MUX_theta_state_inst_n334), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n333) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U132 ( .A1(SlicesFromChi[84]), .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n334) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U131 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n331), .A(
        all_mux_linear_3__MUX_theta_state_inst_n330), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U130 ( .A1(n2), .A2(
        SlicesFromChi[83]), .B1(all_mux_linear_3__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_3__MUX_theta_state_inst_n331), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n330) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U129 ( .A1(SlicesFromChi[83]), .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n331) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U128 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n329), .A(
        all_mux_linear_3__MUX_theta_state_inst_n328), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U127 ( .A1(n2), .A2(
        SlicesFromChi[82]), .B1(all_mux_linear_3__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_3__MUX_theta_state_inst_n329), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n328) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U126 ( .A1(SlicesFromChi[82]), .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n329) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U125 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n327), .A(
        all_mux_linear_3__MUX_theta_state_inst_n326), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U124 ( .A1(n2), .A2(
        SlicesFromChi[81]), .B1(all_mux_linear_3__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_3__MUX_theta_state_inst_n327), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n326) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U123 ( .A1(SlicesFromChi[81]), .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n327) );
  OAI21_X1 all_mux_linear_3__MUX_theta_state_inst_U122 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n325), .A(
        all_mux_linear_3__MUX_theta_state_inst_n324), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_3__MUX_theta_state_inst_U121 ( .A1(n2), .A2(
        SlicesFromChi[80]), .B1(all_mux_linear_3__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_3__MUX_theta_state_inst_n325), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n324) );
  AND2_X1 all_mux_linear_3__MUX_theta_state_inst_U120 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n335), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n332) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U119 ( .A1(SlicesFromChi[80]), .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n325) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U118 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n323), .B(
        all_mux_linear_3__MUX_theta_state_inst_n322), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n335) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U117 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n321), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n319), .A(
        all_mux_linear_3__MUX_theta_state_inst_n318), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[4]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U116 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n321), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n318) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U115 ( .A(SlicesFromChi[79]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n319) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U114 ( .A1(SlicesFromChi[79]), .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n321) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U113 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n317), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n316), .A(
        all_mux_linear_3__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[3]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U112 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n317), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n315) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U111 ( .A(SlicesFromChi[78]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n316) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U110 ( .A1(SlicesFromChi[78]), .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n317) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U109 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n313), .A(
        all_mux_linear_3__MUX_theta_state_inst_n312), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[2]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U108 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n314), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n312) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U107 ( .A1(SlicesFromChi[77]), .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n314) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U106 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n311), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n309), .A(
        all_mux_linear_3__MUX_theta_state_inst_n308), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[24]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n311), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n308) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U104 ( .A(SlicesFromChi[99]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n309) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U103 ( .A1(SlicesFromChi[99]), .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n311) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U102 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n307), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n306), .A(
        all_mux_linear_3__MUX_theta_state_inst_n305), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[23]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U101 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n307), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n305) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U100 ( .A(SlicesFromChi[98]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n306) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U99 ( .A1(SlicesFromChi[98]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n307) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U98 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n304), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n303), .A(
        all_mux_linear_3__MUX_theta_state_inst_n302), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[22]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U97 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n304), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n302) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U96 ( .A1(SlicesFromChi[97]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n304) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n301), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n300), .A(
        all_mux_linear_3__MUX_theta_state_inst_n299), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[21]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n301), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n299) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U93 ( .A(SlicesFromChi[96]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n300) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U92 ( .A1(SlicesFromChi[96]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n301) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n298), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n297), .A(
        all_mux_linear_3__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[20]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n298), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n296) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U89 ( .A(SlicesFromChi[95]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n297) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U88 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n294), .B(
        all_mux_linear_3__MUX_theta_state_inst_n293), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n323) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U87 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n292), .B(
        all_mux_linear_3__MUX_theta_state_inst_n291), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n293) );
  OAI211_X1 all_mux_linear_3__MUX_theta_state_inst_U86 ( .C1(SlicesFromChi[79]), .C2(all_mux_linear_3__MUX_theta_state_inst_n290), .A(
        all_mux_linear_3__MUX_theta_state_inst_n232), .B(
        all_mux_linear_3__MUX_theta_state_inst_n289), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n294) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U85 ( .A1(SlicesFromChi[79]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n289) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n313), .B(SlicesFromChi[78]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n290) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U83 ( .A(SlicesFromChi[77]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n313) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U82 ( .A1(SlicesFromChi[95]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n298) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U81 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n288), .A(
        all_mux_linear_3__MUX_theta_state_inst_n287), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[1]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U80 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n291), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n287) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U79 ( .A(SlicesFromChi[76]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n288) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U78 ( .A1(SlicesFromChi[76]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n291) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n286), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n284), .A(
        all_mux_linear_3__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[19]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n286), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n283) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U75 ( .A(SlicesFromChi[94]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n284) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U74 ( .A1(SlicesFromChi[94]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n286) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U73 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n282), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n281), .A(
        all_mux_linear_3__MUX_theta_state_inst_n280), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[18]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U72 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n282), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n280) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U71 ( .A(SlicesFromChi[93]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n281) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U70 ( .A1(SlicesFromChi[93]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n282) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U69 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n279), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n278), .A(
        all_mux_linear_3__MUX_theta_state_inst_n277), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[17]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U68 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n279), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n277) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U67 ( .A1(SlicesFromChi[92]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n279) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n276), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n275), .A(
        all_mux_linear_3__MUX_theta_state_inst_n274), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[16]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n276), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n274) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U64 ( .A(SlicesFromChi[91]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n275) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U63 ( .A1(SlicesFromChi[91]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n276) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U62 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n273), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n272), .A(
        all_mux_linear_3__MUX_theta_state_inst_n271), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[15]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U61 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n273), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n271) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U60 ( .A(SlicesFromChi[90]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n272) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n269), .B(
        all_mux_linear_3__MUX_theta_state_inst_n268), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n322) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n267), .B(
        all_mux_linear_3__MUX_theta_state_inst_n266), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n268) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U57 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n265), .B(
        all_mux_linear_3__MUX_theta_state_inst_n264), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n267) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U56 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n263), .B(
        all_mux_linear_3__MUX_theta_state_inst_n262), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n269) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U55 ( .A1(SlicesFromChi[90]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n273) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n266), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n260), .A(
        all_mux_linear_3__MUX_theta_state_inst_n259), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[14]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n266), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n259) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U52 ( .A(SlicesFromChi[89]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n260) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U51 ( .A1(SlicesFromChi[89]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n266) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U50 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n264), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n258), .A(
        all_mux_linear_3__MUX_theta_state_inst_n257), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[13]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U49 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n264), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n257) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U48 ( .A(SlicesFromChi[88]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n258) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U47 ( .A1(SlicesFromChi[88]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n264) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U46 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n256), .A(
        all_mux_linear_3__MUX_theta_state_inst_n255), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[12]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U45 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n265), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n255) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U44 ( .A(SlicesFromChi[87]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n256) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U43 ( .A1(SlicesFromChi[87]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n265) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U42 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n262), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n254), .A(
        all_mux_linear_3__MUX_theta_state_inst_n253), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[11]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U41 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n262), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n253) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U40 ( .A(SlicesFromChi[86]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n254) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U39 ( .A1(SlicesFromChi[86]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n262) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U38 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n263), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n252), .A(
        all_mux_linear_3__MUX_theta_state_inst_n251), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[10]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U37 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n263), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n251) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U36 ( .A(SlicesFromChi[85]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n252) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n249), .B(
        all_mux_linear_3__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n295) );
  OAI211_X1 all_mux_linear_3__MUX_theta_state_inst_U34 ( .C1(SlicesFromChi[90]), .C2(all_mux_linear_3__MUX_theta_state_inst_n247), .A(
        all_mux_linear_3__MUX_theta_state_inst_n232), .B(
        all_mux_linear_3__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n248) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U33 ( .A1(SlicesFromChi[90]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n246) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U32 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n278), .B(SlicesFromChi[93]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n247) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U31 ( .A(SlicesFromChi[92]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n278) );
  OAI211_X1 all_mux_linear_3__MUX_theta_state_inst_U30 ( .C1(SlicesFromChi[91]), .C2(SlicesFromChi[94]), .A(all_mux_linear_3__MUX_theta_state_inst_n231), .B(
        all_mux_linear_3__MUX_theta_state_inst_n245), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n249) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[94]), 
        .A2(SlicesFromChi[91]), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n245) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U28 ( .A1(SlicesFromChi[85]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n263) );
  OAI221_X1 all_mux_linear_3__MUX_theta_state_inst_U27 ( .B1(
        all_mux_linear_3__MUX_theta_state_inst_n292), .B2(
        all_mux_linear_3__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_3__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_3__MUX_theta_state_inst_n244), .A(
        all_mux_linear_3__MUX_theta_state_inst_n243), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[0]) );
  NAND3_X1 all_mux_linear_3__MUX_theta_state_inst_U26 ( .A1(
        all_mux_linear_3__MUX_theta_state_inst_n292), .A2(
        all_mux_linear_3__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_3__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n243) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U25 ( .A(SlicesFromChi[75]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n244) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n242), .B(
        all_mux_linear_3__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n250) );
  AOI211_X1 all_mux_linear_3__MUX_theta_state_inst_U23 ( .C1(SlicesFromChi[81]), .C2(SlicesFromChi[82]), .A(Reset), .B(
        all_mux_linear_3__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n241) );
  NOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U22 ( .A1(SlicesFromChi[81]), 
        .A2(SlicesFromChi[82]), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n240) );
  OAI211_X1 all_mux_linear_3__MUX_theta_state_inst_U21 ( .C1(SlicesFromChi[80]), .C2(all_mux_linear_3__MUX_theta_state_inst_n239), .A(
        all_mux_linear_3__MUX_theta_state_inst_n231), .B(
        all_mux_linear_3__MUX_theta_state_inst_n238), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n242) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U20 ( .A1(SlicesFromChi[80]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n239), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n238) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U19 ( .A(SlicesFromChi[84]), 
        .B(SlicesFromChi[83]), .Z(all_mux_linear_3__MUX_theta_state_inst_n239)
         );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U18 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n237), .B(
        all_mux_linear_3__MUX_theta_state_inst_n236), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n270) );
  AOI211_X1 all_mux_linear_3__MUX_theta_state_inst_U17 ( .C1(SlicesFromChi[96]), .C2(SlicesFromChi[99]), .A(Reset), .B(
        all_mux_linear_3__MUX_theta_state_inst_n235), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n236) );
  NOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U16 ( .A1(SlicesFromChi[96]), 
        .A2(SlicesFromChi[99]), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n235) );
  OAI211_X1 all_mux_linear_3__MUX_theta_state_inst_U15 ( .C1(SlicesFromChi[95]), .C2(all_mux_linear_3__MUX_theta_state_inst_n234), .A(
        all_mux_linear_3__MUX_theta_state_inst_n231), .B(
        all_mux_linear_3__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n237) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U14 ( .A1(SlicesFromChi[95]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n233) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U13 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n303), .B(SlicesFromChi[98]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n234) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U12 ( .A(SlicesFromChi[97]), 
        .ZN(all_mux_linear_3__MUX_theta_state_inst_n303) );
  NAND2_X1 all_mux_linear_3__MUX_theta_state_inst_U11 ( .A1(SlicesFromChi[75]), 
        .A2(all_mux_linear_3__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n292) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U10 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n250), .B(
        all_mux_linear_3__MUX_theta_state_inst_n295), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n261) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U9 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n323), .B(
        all_mux_linear_3__MUX_theta_state_inst_n295), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n310) );
  XOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U8 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n270), .B(
        all_mux_linear_3__MUX_theta_state_inst_n250), .Z(
        all_mux_linear_3__MUX_theta_state_inst_n320) );
  XNOR2_X1 all_mux_linear_3__MUX_theta_state_inst_U7 ( .A(
        all_mux_linear_3__MUX_theta_state_inst_n270), .B(
        all_mux_linear_3__MUX_theta_state_inst_n322), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n285) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U6 ( .A(Reset), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n231) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U4 ( .A(n2), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n230) );
  INV_X1 all_mux_linear_3__MUX_theta_state_inst_U3 ( .A(n2), .ZN(
        all_mux_linear_3__MUX_theta_state_inst_n229) );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[75]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[76]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[77]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[78]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[79]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[80]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[81]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[82]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[83]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[84]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[85]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[86]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[87]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[88]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[89]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[90]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[91]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[92]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[93]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[94]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[95]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[96]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[97]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[98]), .QN() );
  DFF_X1 all_mux_linear_3__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_3__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[99]), .QN() );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U116 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n318), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n317), .A(
        all_mux_linear_4__MUX_theta_state_inst_n316), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U115 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[109]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n318), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n316) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U114 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n317), .A(
        all_mux_linear_4__MUX_theta_state_inst_n313), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U113 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[108]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n313) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U112 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n312), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n317), .A(
        all_mux_linear_4__MUX_theta_state_inst_n311), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U111 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[107]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n312), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n311) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U110 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n310), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n317), .A(
        all_mux_linear_4__MUX_theta_state_inst_n309), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U109 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[106]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n310), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n309) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U108 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n308), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n317), .A(
        all_mux_linear_4__MUX_theta_state_inst_n307), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U107 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[105]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n308), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n307) );
  NOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U106 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_4__MUX_theta_state_inst_n306), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n315) );
  NAND2_X1 all_mux_linear_4__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_4__MUX_theta_state_inst_n306), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n317) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U104 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n305), .B(
        all_mux_linear_4__MUX_theta_state_inst_n304), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n306) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U103 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n303), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n302), .A(
        all_mux_linear_4__MUX_theta_state_inst_n301), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[4]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U102 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[104]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n303), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n301) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U101 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n299), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n302), .A(
        all_mux_linear_4__MUX_theta_state_inst_n298), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[3]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U100 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[103]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n299), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n298) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U99 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n297), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n302), .A(
        all_mux_linear_4__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[2]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U98 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[102]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n297), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n296) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U97 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n295), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n294), .A(
        all_mux_linear_4__MUX_theta_state_inst_n293), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[24]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U96 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[124]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n295), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n293) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n294), .A(
        all_mux_linear_4__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[23]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[123]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n290) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U93 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n289), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n294), .A(
        all_mux_linear_4__MUX_theta_state_inst_n288), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[22]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U92 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[122]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n289), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n288) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n287), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n294), .A(
        all_mux_linear_4__MUX_theta_state_inst_n286), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[21]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[121]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n287), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n286) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U89 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n285), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n294), .A(
        all_mux_linear_4__MUX_theta_state_inst_n284), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[20]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U88 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[120]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n285), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n284) );
  NOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U87 ( .A1(n2), .A2(
        all_mux_linear_4__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n292) );
  NAND2_X1 all_mux_linear_4__MUX_theta_state_inst_U86 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_4__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n294) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U85 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n282), .B(
        all_mux_linear_4__MUX_theta_state_inst_n304), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n283) );
  XOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n281), .B(
        all_mux_linear_4__MUX_theta_state_inst_n280), .Z(
        all_mux_linear_4__MUX_theta_state_inst_n304) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U83 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n279), .B(
        all_mux_linear_4__MUX_theta_state_inst_n278), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n280) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U82 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n277), .B(
        all_mux_linear_4__MUX_theta_state_inst_n303), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n278) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U81 ( .A1(Reset), .A2(
        InData[29]), .B1(SlicesFromChi[104]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n303) );
  XOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U80 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n299), .B(
        all_mux_linear_4__MUX_theta_state_inst_n297), .Z(
        all_mux_linear_4__MUX_theta_state_inst_n279) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U79 ( .A1(Reset), .A2(
        InData[27]), .B1(SlicesFromChi[102]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n297) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U78 ( .A1(Reset), .A2(
        InData[28]), .B1(SlicesFromChi[103]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n299) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n277), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n302), .A(
        all_mux_linear_4__MUX_theta_state_inst_n276), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[1]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[101]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n277), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n276) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U75 ( .A1(Reset), .A2(
        InData[26]), .B1(SlicesFromChi[101]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n277) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U74 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n275), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n274), .A(
        all_mux_linear_4__MUX_theta_state_inst_n273), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[19]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U73 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[119]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n275), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n273) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U72 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n271), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n274), .A(
        all_mux_linear_4__MUX_theta_state_inst_n270), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[18]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U71 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[118]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n271), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n270) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U70 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n269), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n274), .A(
        all_mux_linear_4__MUX_theta_state_inst_n268), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[17]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U69 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[117]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n269), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n268) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U68 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n267), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n274), .A(
        all_mux_linear_4__MUX_theta_state_inst_n266), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[16]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U67 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[116]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n267), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n266) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n274), .A(
        all_mux_linear_4__MUX_theta_state_inst_n264), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[15]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[115]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n264) );
  NOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U64 ( .A1(n2), .A2(
        all_mux_linear_4__MUX_theta_state_inst_n263), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n272) );
  NAND2_X1 all_mux_linear_4__MUX_theta_state_inst_U63 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_4__MUX_theta_state_inst_n263), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n274) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U62 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n262), .B(
        all_mux_linear_4__MUX_theta_state_inst_n305), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n263) );
  XOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U61 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n261), .B(
        all_mux_linear_4__MUX_theta_state_inst_n260), .Z(
        all_mux_linear_4__MUX_theta_state_inst_n305) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U60 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n259), .B(
        all_mux_linear_4__MUX_theta_state_inst_n258), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n260) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n257), .B(
        all_mux_linear_4__MUX_theta_state_inst_n256), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n258) );
  XOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n255), .B(
        all_mux_linear_4__MUX_theta_state_inst_n254), .Z(
        all_mux_linear_4__MUX_theta_state_inst_n259) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U57 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n255), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n253), .A(
        all_mux_linear_4__MUX_theta_state_inst_n252), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[14]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U56 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[114]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n255), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n252) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U55 ( .A1(Reset), .A2(
        InData[39]), .B1(SlicesFromChi[114]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n255) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n254), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n253), .A(
        all_mux_linear_4__MUX_theta_state_inst_n250), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[13]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[113]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n254), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n250) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U52 ( .A1(Reset), .A2(
        InData[38]), .B1(SlicesFromChi[113]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n254) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U51 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n256), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n253), .A(
        all_mux_linear_4__MUX_theta_state_inst_n249), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[12]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U50 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[112]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n256), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n249) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U49 ( .A1(Reset), .A2(
        InData[37]), .B1(SlicesFromChi[112]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n256) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U48 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n257), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n253), .A(
        all_mux_linear_4__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[11]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U47 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[111]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n257), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n248) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U46 ( .A1(Reset), .A2(
        InData[36]), .B1(SlicesFromChi[111]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n257) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U45 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n261), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n253), .A(
        all_mux_linear_4__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[10]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U44 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n230), .A2(SlicesFromChi[110]), 
        .B1(all_mux_linear_4__MUX_theta_state_inst_n261), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n251), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n247) );
  NOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U43 ( .A1(n2), .A2(
        all_mux_linear_4__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n251) );
  NAND2_X1 all_mux_linear_4__MUX_theta_state_inst_U42 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_4__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n253) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U41 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n245), .B(
        all_mux_linear_4__MUX_theta_state_inst_n282), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n246) );
  XOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U40 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n275), .B(
        all_mux_linear_4__MUX_theta_state_inst_n244), .Z(
        all_mux_linear_4__MUX_theta_state_inst_n282) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U39 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n243), .B(
        all_mux_linear_4__MUX_theta_state_inst_n242), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n244) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U38 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n267), .B(
        all_mux_linear_4__MUX_theta_state_inst_n265), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n242) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U37 ( .A1(Reset), .A2(
        InData[40]), .B1(SlicesFromChi[115]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n265) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U36 ( .A1(Reset), .A2(
        InData[41]), .B1(SlicesFromChi[116]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n267) );
  XOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n271), .B(
        all_mux_linear_4__MUX_theta_state_inst_n269), .Z(
        all_mux_linear_4__MUX_theta_state_inst_n243) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U34 ( .A1(Reset), .A2(
        InData[42]), .B1(SlicesFromChi[117]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n269) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U33 ( .A1(Reset), .A2(
        InData[43]), .B1(SlicesFromChi[118]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n271) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U32 ( .A1(Reset), .A2(
        InData[44]), .B1(SlicesFromChi[119]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n275) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U31 ( .A1(Reset), .A2(
        InData[35]), .B1(SlicesFromChi[110]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n261) );
  OAI21_X1 all_mux_linear_4__MUX_theta_state_inst_U30 ( .B1(
        all_mux_linear_4__MUX_theta_state_inst_n281), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n302), .A(
        all_mux_linear_4__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[0]) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[100]), .A2(all_mux_linear_4__MUX_theta_state_inst_n230), .B1(
        all_mux_linear_4__MUX_theta_state_inst_n281), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n300), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n241) );
  NOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U28 ( .A1(n2), .A2(
        all_mux_linear_4__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n300) );
  NAND2_X1 all_mux_linear_4__MUX_theta_state_inst_U27 ( .A1(
        all_mux_linear_4__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_4__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n302) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U26 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n262), .B(
        all_mux_linear_4__MUX_theta_state_inst_n245), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n240) );
  XOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U25 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n312), .B(
        all_mux_linear_4__MUX_theta_state_inst_n239), .Z(
        all_mux_linear_4__MUX_theta_state_inst_n245) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n238), .B(
        all_mux_linear_4__MUX_theta_state_inst_n237), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n239) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U23 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n310), .B(
        all_mux_linear_4__MUX_theta_state_inst_n308), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n237) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U22 ( .A1(Reset), .A2(
        InData[30]), .B1(SlicesFromChi[105]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n308) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U21 ( .A1(Reset), .A2(
        InData[31]), .B1(SlicesFromChi[106]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n310) );
  XOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U20 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n314), .B(
        all_mux_linear_4__MUX_theta_state_inst_n318), .Z(
        all_mux_linear_4__MUX_theta_state_inst_n238) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U19 ( .A1(Reset), .A2(
        InData[34]), .B1(SlicesFromChi[109]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n318) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U18 ( .A1(Reset), .A2(
        InData[33]), .B1(SlicesFromChi[108]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n314) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U17 ( .A1(Reset), .A2(
        InData[32]), .B1(SlicesFromChi[107]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n312) );
  XOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U16 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n295), .B(
        all_mux_linear_4__MUX_theta_state_inst_n236), .Z(
        all_mux_linear_4__MUX_theta_state_inst_n262) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U15 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n235), .B(
        all_mux_linear_4__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n236) );
  XNOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U14 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n287), .B(
        all_mux_linear_4__MUX_theta_state_inst_n285), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n234) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U13 ( .A1(Reset), .A2(
        InData[45]), .B1(SlicesFromChi[120]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n285) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U12 ( .A1(Reset), .A2(
        InData[46]), .B1(SlicesFromChi[121]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n287) );
  XOR2_X1 all_mux_linear_4__MUX_theta_state_inst_U11 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n291), .B(
        all_mux_linear_4__MUX_theta_state_inst_n289), .Z(
        all_mux_linear_4__MUX_theta_state_inst_n235) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U10 ( .A1(Reset), .A2(
        InData[47]), .B1(SlicesFromChi[122]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n289) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U9 ( .A1(Reset), .A2(
        InData[48]), .B1(SlicesFromChi[123]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n291) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U8 ( .A1(Reset), .A2(
        InData[49]), .B1(SlicesFromChi[124]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n295) );
  AOI22_X1 all_mux_linear_4__MUX_theta_state_inst_U7 ( .A1(Reset), .A2(
        InData[25]), .B1(SlicesFromChi[100]), .B2(
        all_mux_linear_4__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n281) );
  INV_X2 all_mux_linear_4__MUX_theta_state_inst_U6 ( .A(
        all_mux_linear_4__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n230) );
  INV_X1 all_mux_linear_4__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n233) );
  INV_X1 all_mux_linear_4__MUX_theta_state_inst_U4 ( .A(Reset), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_4__MUX_theta_state_inst_U3 ( .A(n2), .ZN(
        all_mux_linear_4__MUX_theta_state_inst_n231) );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[100]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[101]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[102]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[103]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[104]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[105]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[106]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[107]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[108]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[109]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[110]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[111]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[112]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[113]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[114]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[115]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[116]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[117]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[118]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[119]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[120]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[121]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[122]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[123]), .QN() );
  DFF_X1 all_mux_linear_4__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_4__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[124]), .QN() );
  OAI21_X1 all_mux_linear_5__MUX_theta_state_inst_U134 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n335), .A(
        all_mux_linear_5__MUX_theta_state_inst_n334), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_5__MUX_theta_state_inst_U133 ( .A1(n3), .A2(
        SlicesFromChi[134]), .B1(all_mux_linear_5__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_5__MUX_theta_state_inst_n335), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n334) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U132 ( .A1(
        SlicesFromChi[134]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n335) );
  OAI21_X1 all_mux_linear_5__MUX_theta_state_inst_U131 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n332), .A(
        all_mux_linear_5__MUX_theta_state_inst_n331), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_5__MUX_theta_state_inst_U130 ( .A1(n3), .A2(
        SlicesFromChi[133]), .B1(all_mux_linear_5__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_5__MUX_theta_state_inst_n332), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n331) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U129 ( .A1(
        SlicesFromChi[133]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n332) );
  OAI21_X1 all_mux_linear_5__MUX_theta_state_inst_U128 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n330), .A(
        all_mux_linear_5__MUX_theta_state_inst_n329), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_5__MUX_theta_state_inst_U127 ( .A1(n3), .A2(
        SlicesFromChi[132]), .B1(all_mux_linear_5__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_5__MUX_theta_state_inst_n330), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n329) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U126 ( .A1(
        SlicesFromChi[132]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n330) );
  OAI21_X1 all_mux_linear_5__MUX_theta_state_inst_U125 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n328), .A(
        all_mux_linear_5__MUX_theta_state_inst_n327), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_5__MUX_theta_state_inst_U124 ( .A1(n3), .A2(
        SlicesFromChi[131]), .B1(all_mux_linear_5__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_5__MUX_theta_state_inst_n328), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n327) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U123 ( .A1(
        SlicesFromChi[131]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n328) );
  OAI21_X1 all_mux_linear_5__MUX_theta_state_inst_U122 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n326), .A(
        all_mux_linear_5__MUX_theta_state_inst_n325), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_5__MUX_theta_state_inst_U121 ( .A1(n3), .A2(
        SlicesFromChi[130]), .B1(all_mux_linear_5__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_5__MUX_theta_state_inst_n326), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n325) );
  AND2_X1 all_mux_linear_5__MUX_theta_state_inst_U120 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n336), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n333) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U119 ( .A1(
        SlicesFromChi[130]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n326) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U118 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n324), .B(
        all_mux_linear_5__MUX_theta_state_inst_n323), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n336) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U117 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n322), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n320), .A(
        all_mux_linear_5__MUX_theta_state_inst_n319), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[4]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U116 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n322), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n319) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U115 ( .A(SlicesFromChi[129]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n320) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U114 ( .A1(
        SlicesFromChi[129]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n322) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U113 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n318), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n317), .A(
        all_mux_linear_5__MUX_theta_state_inst_n316), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[3]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U112 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n318), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n316) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U111 ( .A(SlicesFromChi[128]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n317) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U110 ( .A1(
        SlicesFromChi[128]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n318) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U109 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n315), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n314), .A(
        all_mux_linear_5__MUX_theta_state_inst_n313), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[2]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U108 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n315), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n313) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U107 ( .A1(
        SlicesFromChi[127]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n315) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U106 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n312), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n310), .A(
        all_mux_linear_5__MUX_theta_state_inst_n309), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[24]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n312), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n309) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U104 ( .A(SlicesFromChi[149]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n310) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U103 ( .A1(
        SlicesFromChi[149]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n312) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U102 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n308), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n307), .A(
        all_mux_linear_5__MUX_theta_state_inst_n306), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[23]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U101 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n308), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n306) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U100 ( .A(SlicesFromChi[148]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n307) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U99 ( .A1(SlicesFromChi[148]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n308) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U98 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n305), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n304), .A(
        all_mux_linear_5__MUX_theta_state_inst_n303), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[22]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U97 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n305), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n303) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U96 ( .A1(SlicesFromChi[147]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n305) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n302), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n301), .A(
        all_mux_linear_5__MUX_theta_state_inst_n300), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[21]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n302), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n300) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U93 ( .A(SlicesFromChi[146]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n301) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U92 ( .A1(SlicesFromChi[146]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n302) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n299), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n298), .A(
        all_mux_linear_5__MUX_theta_state_inst_n297), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[20]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n299), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n297) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U89 ( .A(SlicesFromChi[145]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n298) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U88 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n295), .B(
        all_mux_linear_5__MUX_theta_state_inst_n294), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n324) );
  XOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U87 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n293), .B(
        all_mux_linear_5__MUX_theta_state_inst_n292), .Z(
        all_mux_linear_5__MUX_theta_state_inst_n294) );
  OAI211_X1 all_mux_linear_5__MUX_theta_state_inst_U86 ( .C1(
        SlicesFromChi[129]), .C2(all_mux_linear_5__MUX_theta_state_inst_n291), 
        .A(all_mux_linear_5__MUX_theta_state_inst_n233), .B(
        all_mux_linear_5__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n295) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U85 ( .A1(SlicesFromChi[129]), .A2(all_mux_linear_5__MUX_theta_state_inst_n291), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n290) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n314), .B(SlicesFromChi[128]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n291) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U83 ( .A(SlicesFromChi[127]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n314) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U82 ( .A1(SlicesFromChi[145]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n299) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U81 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n292), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n289), .A(
        all_mux_linear_5__MUX_theta_state_inst_n288), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[1]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U80 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n292), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n288) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U79 ( .A(SlicesFromChi[126]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n289) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U78 ( .A1(SlicesFromChi[126]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n292) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n287), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n285), .A(
        all_mux_linear_5__MUX_theta_state_inst_n284), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[19]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n287), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n284) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U75 ( .A(SlicesFromChi[144]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n285) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U74 ( .A1(SlicesFromChi[144]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n287) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U73 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n283), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n282), .A(
        all_mux_linear_5__MUX_theta_state_inst_n281), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[18]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U72 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n283), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n281) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U71 ( .A(SlicesFromChi[143]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n282) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U70 ( .A1(SlicesFromChi[143]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n283) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U69 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n280), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n279), .A(
        all_mux_linear_5__MUX_theta_state_inst_n278), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[17]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U68 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n280), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n278) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U67 ( .A1(SlicesFromChi[142]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n280) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n277), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n276), .A(
        all_mux_linear_5__MUX_theta_state_inst_n275), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[16]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n277), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n275) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U64 ( .A(SlicesFromChi[141]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n276) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U63 ( .A1(SlicesFromChi[141]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n277) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U62 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n274), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n273), .A(
        all_mux_linear_5__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[15]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U61 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n274), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n272) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U60 ( .A(SlicesFromChi[140]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n273) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n270), .B(
        all_mux_linear_5__MUX_theta_state_inst_n269), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n323) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n268), .B(
        all_mux_linear_5__MUX_theta_state_inst_n267), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n269) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U57 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n266), .B(
        all_mux_linear_5__MUX_theta_state_inst_n265), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n268) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U56 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n264), .B(
        all_mux_linear_5__MUX_theta_state_inst_n263), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n270) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U55 ( .A1(SlicesFromChi[140]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n274) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n267), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n261), .A(
        all_mux_linear_5__MUX_theta_state_inst_n260), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[14]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n267), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n260) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U52 ( .A(SlicesFromChi[139]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n261) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U51 ( .A1(SlicesFromChi[139]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n267) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U50 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n259), .A(
        all_mux_linear_5__MUX_theta_state_inst_n258), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[13]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U49 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n265), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n258) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U48 ( .A(SlicesFromChi[138]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n259) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U47 ( .A1(SlicesFromChi[138]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n265) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U46 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n266), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n257), .A(
        all_mux_linear_5__MUX_theta_state_inst_n256), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[12]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U45 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n266), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n256) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U44 ( .A(SlicesFromChi[137]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n257) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U43 ( .A1(SlicesFromChi[137]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n266) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U42 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n263), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n255), .A(
        all_mux_linear_5__MUX_theta_state_inst_n254), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[11]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U41 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n263), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n254) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U40 ( .A(SlicesFromChi[136]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n255) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U39 ( .A1(SlicesFromChi[136]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n263) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U38 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n264), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n253), .A(
        all_mux_linear_5__MUX_theta_state_inst_n252), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[10]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U37 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n264), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n252) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U36 ( .A(SlicesFromChi[135]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n253) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n250), .B(
        all_mux_linear_5__MUX_theta_state_inst_n249), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n296) );
  OAI211_X1 all_mux_linear_5__MUX_theta_state_inst_U34 ( .C1(
        SlicesFromChi[140]), .C2(all_mux_linear_5__MUX_theta_state_inst_n248), 
        .A(all_mux_linear_5__MUX_theta_state_inst_n233), .B(
        all_mux_linear_5__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n249) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U33 ( .A1(SlicesFromChi[140]), .A2(all_mux_linear_5__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n247) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U32 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n279), .B(SlicesFromChi[143]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n248) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U31 ( .A(SlicesFromChi[142]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n279) );
  OAI211_X1 all_mux_linear_5__MUX_theta_state_inst_U30 ( .C1(
        SlicesFromChi[141]), .C2(SlicesFromChi[144]), .A(
        all_mux_linear_5__MUX_theta_state_inst_n232), .B(
        all_mux_linear_5__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n250) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[144]), .A2(SlicesFromChi[141]), .ZN(all_mux_linear_5__MUX_theta_state_inst_n246) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U28 ( .A1(SlicesFromChi[135]), .A2(all_mux_linear_5__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n264) );
  OAI221_X1 all_mux_linear_5__MUX_theta_state_inst_U27 ( .B1(
        all_mux_linear_5__MUX_theta_state_inst_n293), .B2(
        all_mux_linear_5__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_5__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_5__MUX_theta_state_inst_n245), .A(
        all_mux_linear_5__MUX_theta_state_inst_n244), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[0]) );
  NAND3_X1 all_mux_linear_5__MUX_theta_state_inst_U26 ( .A1(
        all_mux_linear_5__MUX_theta_state_inst_n293), .A2(
        all_mux_linear_5__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_5__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n244) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U25 ( .A(SlicesFromChi[125]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n245) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n243), .B(
        all_mux_linear_5__MUX_theta_state_inst_n242), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n251) );
  AOI211_X1 all_mux_linear_5__MUX_theta_state_inst_U23 ( .C1(
        SlicesFromChi[131]), .C2(SlicesFromChi[132]), .A(Reset), .B(
        all_mux_linear_5__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n242) );
  NOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U22 ( .A1(SlicesFromChi[131]), 
        .A2(SlicesFromChi[132]), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n241) );
  OAI211_X1 all_mux_linear_5__MUX_theta_state_inst_U21 ( .C1(
        SlicesFromChi[130]), .C2(all_mux_linear_5__MUX_theta_state_inst_n240), 
        .A(all_mux_linear_5__MUX_theta_state_inst_n232), .B(
        all_mux_linear_5__MUX_theta_state_inst_n239), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n243) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U20 ( .A1(SlicesFromChi[130]), .A2(all_mux_linear_5__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n239) );
  XOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U19 ( .A(SlicesFromChi[134]), 
        .B(SlicesFromChi[133]), .Z(all_mux_linear_5__MUX_theta_state_inst_n240) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U18 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n238), .B(
        all_mux_linear_5__MUX_theta_state_inst_n237), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n271) );
  AOI211_X1 all_mux_linear_5__MUX_theta_state_inst_U17 ( .C1(
        SlicesFromChi[146]), .C2(SlicesFromChi[149]), .A(Reset), .B(
        all_mux_linear_5__MUX_theta_state_inst_n236), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n237) );
  NOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U16 ( .A1(SlicesFromChi[146]), 
        .A2(SlicesFromChi[149]), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n236) );
  OAI211_X1 all_mux_linear_5__MUX_theta_state_inst_U15 ( .C1(
        SlicesFromChi[145]), .C2(all_mux_linear_5__MUX_theta_state_inst_n235), 
        .A(all_mux_linear_5__MUX_theta_state_inst_n232), .B(
        all_mux_linear_5__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n238) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U14 ( .A1(SlicesFromChi[145]), .A2(all_mux_linear_5__MUX_theta_state_inst_n235), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n234) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U13 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n304), .B(SlicesFromChi[148]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n235) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U12 ( .A(SlicesFromChi[147]), 
        .ZN(all_mux_linear_5__MUX_theta_state_inst_n304) );
  NAND2_X1 all_mux_linear_5__MUX_theta_state_inst_U11 ( .A1(SlicesFromChi[125]), .A2(all_mux_linear_5__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n293) );
  XOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U10 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n271), .B(
        all_mux_linear_5__MUX_theta_state_inst_n251), .Z(
        all_mux_linear_5__MUX_theta_state_inst_n321) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U9 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n271), .B(
        all_mux_linear_5__MUX_theta_state_inst_n323), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n286) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U8 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n251), .B(
        all_mux_linear_5__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n262) );
  XNOR2_X1 all_mux_linear_5__MUX_theta_state_inst_U7 ( .A(
        all_mux_linear_5__MUX_theta_state_inst_n324), .B(
        all_mux_linear_5__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n311) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U6 ( .A(Reset), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U5 ( .A(n3), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n231) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U4 ( .A(n3), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n230) );
  INV_X1 all_mux_linear_5__MUX_theta_state_inst_U3 ( .A(Reset), .ZN(
        all_mux_linear_5__MUX_theta_state_inst_n233) );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[125]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[126]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[127]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[128]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[129]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[130]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[131]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[132]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[133]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[134]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[135]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[136]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[137]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[138]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[139]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[140]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[141]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[142]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[143]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[144]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[145]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[146]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[147]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[148]), .QN() );
  DFF_X1 all_mux_linear_5__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_5__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[149]), .QN() );
  OAI21_X1 all_mux_linear_6__MUX_theta_state_inst_U134 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n334), .A(
        all_mux_linear_6__MUX_theta_state_inst_n333), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_6__MUX_theta_state_inst_U133 ( .A1(n4), .A2(
        SlicesFromChi[159]), .B1(all_mux_linear_6__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_6__MUX_theta_state_inst_n334), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n333) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U132 ( .A1(
        SlicesFromChi[159]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n334) );
  OAI21_X1 all_mux_linear_6__MUX_theta_state_inst_U131 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n331), .A(
        all_mux_linear_6__MUX_theta_state_inst_n330), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_6__MUX_theta_state_inst_U130 ( .A1(n4), .A2(
        SlicesFromChi[158]), .B1(all_mux_linear_6__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_6__MUX_theta_state_inst_n331), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n330) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U129 ( .A1(
        SlicesFromChi[158]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n331) );
  OAI21_X1 all_mux_linear_6__MUX_theta_state_inst_U128 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n329), .A(
        all_mux_linear_6__MUX_theta_state_inst_n328), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_6__MUX_theta_state_inst_U127 ( .A1(n4), .A2(
        SlicesFromChi[157]), .B1(all_mux_linear_6__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_6__MUX_theta_state_inst_n329), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n328) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U126 ( .A1(
        SlicesFromChi[157]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n329) );
  OAI21_X1 all_mux_linear_6__MUX_theta_state_inst_U125 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n327), .A(
        all_mux_linear_6__MUX_theta_state_inst_n326), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_6__MUX_theta_state_inst_U124 ( .A1(n4), .A2(
        SlicesFromChi[156]), .B1(all_mux_linear_6__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_6__MUX_theta_state_inst_n327), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n326) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U123 ( .A1(
        SlicesFromChi[156]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n327) );
  OAI21_X1 all_mux_linear_6__MUX_theta_state_inst_U122 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n335), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n325), .A(
        all_mux_linear_6__MUX_theta_state_inst_n324), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_6__MUX_theta_state_inst_U121 ( .A1(n4), .A2(
        SlicesFromChi[155]), .B1(all_mux_linear_6__MUX_theta_state_inst_n332), 
        .B2(all_mux_linear_6__MUX_theta_state_inst_n325), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n324) );
  AND2_X1 all_mux_linear_6__MUX_theta_state_inst_U120 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n335), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n332) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U119 ( .A1(
        SlicesFromChi[155]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n325) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U118 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n323), .B(
        all_mux_linear_6__MUX_theta_state_inst_n322), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n335) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U117 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n321), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n319), .A(
        all_mux_linear_6__MUX_theta_state_inst_n318), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[4]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U116 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n321), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n318) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U115 ( .A(SlicesFromChi[154]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n319) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U114 ( .A1(
        SlicesFromChi[154]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n321) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U113 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n317), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n316), .A(
        all_mux_linear_6__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[3]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U112 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n317), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n315) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U111 ( .A(SlicesFromChi[153]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n316) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U110 ( .A1(
        SlicesFromChi[153]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n317) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U109 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n313), .A(
        all_mux_linear_6__MUX_theta_state_inst_n312), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[2]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U108 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n314), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n312) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U107 ( .A1(
        SlicesFromChi[152]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n314) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U106 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n311), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n309), .A(
        all_mux_linear_6__MUX_theta_state_inst_n308), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[24]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n311), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n308) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U104 ( .A(SlicesFromChi[174]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n309) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U103 ( .A1(
        SlicesFromChi[174]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n311) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U102 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n307), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n306), .A(
        all_mux_linear_6__MUX_theta_state_inst_n305), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[23]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U101 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n307), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n305) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U100 ( .A(SlicesFromChi[173]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n306) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U99 ( .A1(SlicesFromChi[173]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n307) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U98 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n304), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n303), .A(
        all_mux_linear_6__MUX_theta_state_inst_n302), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[22]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U97 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n304), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n302) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U96 ( .A1(SlicesFromChi[172]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n304) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n301), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n300), .A(
        all_mux_linear_6__MUX_theta_state_inst_n299), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[21]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n301), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n299) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U93 ( .A(SlicesFromChi[171]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n300) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U92 ( .A1(SlicesFromChi[171]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n301) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n298), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n310), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n297), .A(
        all_mux_linear_6__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[20]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n298), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n310), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n296) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U89 ( .A(SlicesFromChi[170]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n297) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U88 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n294), .B(
        all_mux_linear_6__MUX_theta_state_inst_n293), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n323) );
  XOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U87 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n292), .B(
        all_mux_linear_6__MUX_theta_state_inst_n291), .Z(
        all_mux_linear_6__MUX_theta_state_inst_n293) );
  OAI211_X1 all_mux_linear_6__MUX_theta_state_inst_U86 ( .C1(
        SlicesFromChi[154]), .C2(all_mux_linear_6__MUX_theta_state_inst_n290), 
        .A(all_mux_linear_6__MUX_theta_state_inst_n232), .B(
        all_mux_linear_6__MUX_theta_state_inst_n289), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n294) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U85 ( .A1(SlicesFromChi[154]), .A2(all_mux_linear_6__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n289) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n313), .B(SlicesFromChi[153]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n290) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U83 ( .A(SlicesFromChi[152]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n313) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U82 ( .A1(SlicesFromChi[170]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n298) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U81 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n288), .A(
        all_mux_linear_6__MUX_theta_state_inst_n287), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[1]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U80 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n291), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n287) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U79 ( .A(SlicesFromChi[151]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n288) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U78 ( .A1(SlicesFromChi[151]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n291) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n286), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n284), .A(
        all_mux_linear_6__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[19]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n286), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n283) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U75 ( .A(SlicesFromChi[169]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n284) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U74 ( .A1(SlicesFromChi[169]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n286) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U73 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n282), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n281), .A(
        all_mux_linear_6__MUX_theta_state_inst_n280), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[18]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U72 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n282), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n280) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U71 ( .A(SlicesFromChi[168]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n281) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U70 ( .A1(SlicesFromChi[168]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n282) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U69 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n279), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n278), .A(
        all_mux_linear_6__MUX_theta_state_inst_n277), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[17]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U68 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n279), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n277) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U67 ( .A1(SlicesFromChi[167]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n279) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n276), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n229), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n275), .A(
        all_mux_linear_6__MUX_theta_state_inst_n274), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[16]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n276), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n274) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U64 ( .A(SlicesFromChi[166]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n275) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U63 ( .A1(SlicesFromChi[166]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n276) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U62 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n273), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n285), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n272), .A(
        all_mux_linear_6__MUX_theta_state_inst_n271), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[15]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U61 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n273), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n285), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n271) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U60 ( .A(SlicesFromChi[165]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n272) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n269), .B(
        all_mux_linear_6__MUX_theta_state_inst_n268), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n322) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n267), .B(
        all_mux_linear_6__MUX_theta_state_inst_n266), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n268) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U57 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n265), .B(
        all_mux_linear_6__MUX_theta_state_inst_n264), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n267) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U56 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n263), .B(
        all_mux_linear_6__MUX_theta_state_inst_n262), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n269) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U55 ( .A1(SlicesFromChi[165]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n273) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n266), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n260), .A(
        all_mux_linear_6__MUX_theta_state_inst_n259), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[14]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n266), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n259) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U52 ( .A(SlicesFromChi[164]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n260) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U51 ( .A1(SlicesFromChi[164]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n266) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U50 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n264), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n258), .A(
        all_mux_linear_6__MUX_theta_state_inst_n257), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[13]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U49 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n264), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n257) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U48 ( .A(SlicesFromChi[163]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n258) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U47 ( .A1(SlicesFromChi[163]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n264) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U46 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n256), .A(
        all_mux_linear_6__MUX_theta_state_inst_n255), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[12]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U45 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n265), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n255) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U44 ( .A(SlicesFromChi[162]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n256) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U43 ( .A1(SlicesFromChi[162]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n265) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U42 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n262), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n254), .A(
        all_mux_linear_6__MUX_theta_state_inst_n253), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[11]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U41 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n262), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n253) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U40 ( .A(SlicesFromChi[161]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n254) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U39 ( .A1(SlicesFromChi[161]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n262) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U38 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n263), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n261), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n252), .A(
        all_mux_linear_6__MUX_theta_state_inst_n251), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[10]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U37 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n263), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n261), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n251) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U36 ( .A(SlicesFromChi[160]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n252) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n249), .B(
        all_mux_linear_6__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n295) );
  OAI211_X1 all_mux_linear_6__MUX_theta_state_inst_U34 ( .C1(
        SlicesFromChi[165]), .C2(all_mux_linear_6__MUX_theta_state_inst_n247), 
        .A(all_mux_linear_6__MUX_theta_state_inst_n232), .B(
        all_mux_linear_6__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n248) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U33 ( .A1(SlicesFromChi[165]), .A2(all_mux_linear_6__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n246) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U32 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n278), .B(SlicesFromChi[168]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n247) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U31 ( .A(SlicesFromChi[167]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n278) );
  OAI211_X1 all_mux_linear_6__MUX_theta_state_inst_U30 ( .C1(
        SlicesFromChi[166]), .C2(SlicesFromChi[169]), .A(
        all_mux_linear_6__MUX_theta_state_inst_n231), .B(
        all_mux_linear_6__MUX_theta_state_inst_n245), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n249) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[169]), .A2(SlicesFromChi[166]), .ZN(all_mux_linear_6__MUX_theta_state_inst_n245) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U28 ( .A1(SlicesFromChi[160]), .A2(all_mux_linear_6__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n263) );
  OAI221_X1 all_mux_linear_6__MUX_theta_state_inst_U27 ( .B1(
        all_mux_linear_6__MUX_theta_state_inst_n292), .B2(
        all_mux_linear_6__MUX_theta_state_inst_n320), .C1(
        all_mux_linear_6__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_6__MUX_theta_state_inst_n244), .A(
        all_mux_linear_6__MUX_theta_state_inst_n243), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[0]) );
  NAND3_X1 all_mux_linear_6__MUX_theta_state_inst_U26 ( .A1(
        all_mux_linear_6__MUX_theta_state_inst_n292), .A2(
        all_mux_linear_6__MUX_theta_state_inst_n320), .A3(
        all_mux_linear_6__MUX_theta_state_inst_n229), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n243) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U25 ( .A(SlicesFromChi[150]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n244) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n242), .B(
        all_mux_linear_6__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n250) );
  AOI211_X1 all_mux_linear_6__MUX_theta_state_inst_U23 ( .C1(
        SlicesFromChi[156]), .C2(SlicesFromChi[157]), .A(Reset), .B(
        all_mux_linear_6__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n241) );
  NOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U22 ( .A1(SlicesFromChi[156]), 
        .A2(SlicesFromChi[157]), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n240) );
  OAI211_X1 all_mux_linear_6__MUX_theta_state_inst_U21 ( .C1(
        SlicesFromChi[155]), .C2(all_mux_linear_6__MUX_theta_state_inst_n239), 
        .A(all_mux_linear_6__MUX_theta_state_inst_n231), .B(
        all_mux_linear_6__MUX_theta_state_inst_n238), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n242) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U20 ( .A1(SlicesFromChi[155]), .A2(all_mux_linear_6__MUX_theta_state_inst_n239), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n238) );
  XOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U19 ( .A(SlicesFromChi[159]), 
        .B(SlicesFromChi[158]), .Z(all_mux_linear_6__MUX_theta_state_inst_n239) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U18 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n237), .B(
        all_mux_linear_6__MUX_theta_state_inst_n236), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n270) );
  AOI211_X1 all_mux_linear_6__MUX_theta_state_inst_U17 ( .C1(
        SlicesFromChi[171]), .C2(SlicesFromChi[174]), .A(Reset), .B(
        all_mux_linear_6__MUX_theta_state_inst_n235), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n236) );
  NOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U16 ( .A1(SlicesFromChi[171]), 
        .A2(SlicesFromChi[174]), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n235) );
  OAI211_X1 all_mux_linear_6__MUX_theta_state_inst_U15 ( .C1(
        SlicesFromChi[170]), .C2(all_mux_linear_6__MUX_theta_state_inst_n234), 
        .A(all_mux_linear_6__MUX_theta_state_inst_n231), .B(
        all_mux_linear_6__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n237) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U14 ( .A1(SlicesFromChi[170]), .A2(all_mux_linear_6__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n233) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U13 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n303), .B(SlicesFromChi[173]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n234) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U12 ( .A(SlicesFromChi[172]), 
        .ZN(all_mux_linear_6__MUX_theta_state_inst_n303) );
  NAND2_X1 all_mux_linear_6__MUX_theta_state_inst_U11 ( .A1(SlicesFromChi[150]), .A2(all_mux_linear_6__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n292) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U10 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n323), .B(
        all_mux_linear_6__MUX_theta_state_inst_n295), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n310) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U9 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n250), .B(
        all_mux_linear_6__MUX_theta_state_inst_n295), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n261) );
  XOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U8 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n270), .B(
        all_mux_linear_6__MUX_theta_state_inst_n250), .Z(
        all_mux_linear_6__MUX_theta_state_inst_n320) );
  XNOR2_X1 all_mux_linear_6__MUX_theta_state_inst_U7 ( .A(
        all_mux_linear_6__MUX_theta_state_inst_n270), .B(
        all_mux_linear_6__MUX_theta_state_inst_n322), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n285) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U6 ( .A(Reset), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n231) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U4 ( .A(n4), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n230) );
  INV_X1 all_mux_linear_6__MUX_theta_state_inst_U3 ( .A(n4), .ZN(
        all_mux_linear_6__MUX_theta_state_inst_n229) );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[150]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[151]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[152]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[153]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[154]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[155]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[156]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[157]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[158]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[159]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[160]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[161]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[162]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[163]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[164]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[165]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[166]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[167]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[168]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[169]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[170]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[171]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[172]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[173]), .QN() );
  DFF_X1 all_mux_linear_6__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_6__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[174]), .QN() );
  OAI21_X1 all_mux_linear_7__MUX_theta_state_inst_U134 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n335), .A(
        all_mux_linear_7__MUX_theta_state_inst_n334), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_7__MUX_theta_state_inst_U133 ( .A1(n4), .A2(
        SlicesFromChi[184]), .B1(all_mux_linear_7__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_7__MUX_theta_state_inst_n335), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n334) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U132 ( .A1(
        SlicesFromChi[184]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n335) );
  OAI21_X1 all_mux_linear_7__MUX_theta_state_inst_U131 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n332), .A(
        all_mux_linear_7__MUX_theta_state_inst_n331), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_7__MUX_theta_state_inst_U130 ( .A1(n4), .A2(
        SlicesFromChi[183]), .B1(all_mux_linear_7__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_7__MUX_theta_state_inst_n332), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n331) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U129 ( .A1(
        SlicesFromChi[183]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n332) );
  OAI21_X1 all_mux_linear_7__MUX_theta_state_inst_U128 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n330), .A(
        all_mux_linear_7__MUX_theta_state_inst_n329), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_7__MUX_theta_state_inst_U127 ( .A1(n4), .A2(
        SlicesFromChi[182]), .B1(all_mux_linear_7__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_7__MUX_theta_state_inst_n330), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n329) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U126 ( .A1(
        SlicesFromChi[182]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n330) );
  OAI21_X1 all_mux_linear_7__MUX_theta_state_inst_U125 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n328), .A(
        all_mux_linear_7__MUX_theta_state_inst_n327), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_7__MUX_theta_state_inst_U124 ( .A1(n4), .A2(
        SlicesFromChi[181]), .B1(all_mux_linear_7__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_7__MUX_theta_state_inst_n328), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n327) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U123 ( .A1(
        SlicesFromChi[181]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n328) );
  OAI21_X1 all_mux_linear_7__MUX_theta_state_inst_U122 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n336), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n326), .A(
        all_mux_linear_7__MUX_theta_state_inst_n325), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_7__MUX_theta_state_inst_U121 ( .A1(n4), .A2(
        SlicesFromChi[180]), .B1(all_mux_linear_7__MUX_theta_state_inst_n333), 
        .B2(all_mux_linear_7__MUX_theta_state_inst_n326), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n325) );
  AND2_X1 all_mux_linear_7__MUX_theta_state_inst_U120 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n336), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n333) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U119 ( .A1(
        SlicesFromChi[180]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n326) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U118 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n324), .B(
        all_mux_linear_7__MUX_theta_state_inst_n323), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n336) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U117 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n322), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n320), .A(
        all_mux_linear_7__MUX_theta_state_inst_n319), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[4]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U116 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n322), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n319) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U115 ( .A(SlicesFromChi[179]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n320) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U114 ( .A1(
        SlicesFromChi[179]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n322) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U113 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n318), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n317), .A(
        all_mux_linear_7__MUX_theta_state_inst_n316), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[3]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U112 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n318), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n316) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U111 ( .A(SlicesFromChi[178]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n317) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U110 ( .A1(
        SlicesFromChi[178]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n318) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U109 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n315), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n314), .A(
        all_mux_linear_7__MUX_theta_state_inst_n313), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[2]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U108 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n315), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n313) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U107 ( .A1(
        SlicesFromChi[177]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n315) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U106 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n312), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n310), .A(
        all_mux_linear_7__MUX_theta_state_inst_n309), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[24]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n312), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n309) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U104 ( .A(SlicesFromChi[199]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n310) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U103 ( .A1(
        SlicesFromChi[199]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n312) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U102 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n308), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n307), .A(
        all_mux_linear_7__MUX_theta_state_inst_n306), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[23]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U101 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n308), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n306) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U100 ( .A(SlicesFromChi[198]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n307) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U99 ( .A1(SlicesFromChi[198]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n308) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U98 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n305), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n304), .A(
        all_mux_linear_7__MUX_theta_state_inst_n303), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[22]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U97 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n305), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n303) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U96 ( .A1(SlicesFromChi[197]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n305) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n302), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n301), .A(
        all_mux_linear_7__MUX_theta_state_inst_n300), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[21]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n302), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n300) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U93 ( .A(SlicesFromChi[196]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n301) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U92 ( .A1(SlicesFromChi[196]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n302) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n299), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n311), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n298), .A(
        all_mux_linear_7__MUX_theta_state_inst_n297), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[20]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n299), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n311), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n297) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U89 ( .A(SlicesFromChi[195]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n298) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U88 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n295), .B(
        all_mux_linear_7__MUX_theta_state_inst_n294), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n324) );
  XOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U87 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n293), .B(
        all_mux_linear_7__MUX_theta_state_inst_n292), .Z(
        all_mux_linear_7__MUX_theta_state_inst_n294) );
  OAI211_X1 all_mux_linear_7__MUX_theta_state_inst_U86 ( .C1(
        SlicesFromChi[179]), .C2(all_mux_linear_7__MUX_theta_state_inst_n291), 
        .A(all_mux_linear_7__MUX_theta_state_inst_n233), .B(
        all_mux_linear_7__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n295) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U85 ( .A1(SlicesFromChi[179]), .A2(all_mux_linear_7__MUX_theta_state_inst_n291), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n290) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n314), .B(SlicesFromChi[178]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n291) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U83 ( .A(SlicesFromChi[177]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n314) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U82 ( .A1(SlicesFromChi[195]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n299) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U81 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n292), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n289), .A(
        all_mux_linear_7__MUX_theta_state_inst_n288), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[1]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U80 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n292), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n288) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U79 ( .A(SlicesFromChi[176]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n289) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U78 ( .A1(SlicesFromChi[176]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n292) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n287), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n285), .A(
        all_mux_linear_7__MUX_theta_state_inst_n284), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[19]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n287), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n284) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U75 ( .A(SlicesFromChi[194]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n285) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U74 ( .A1(SlicesFromChi[194]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n287) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U73 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n283), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n282), .A(
        all_mux_linear_7__MUX_theta_state_inst_n281), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[18]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U72 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n283), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n230), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n281) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U71 ( .A(SlicesFromChi[193]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n282) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U70 ( .A1(SlicesFromChi[193]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n283) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U69 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n280), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n279), .A(
        all_mux_linear_7__MUX_theta_state_inst_n278), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[17]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U68 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n280), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n278) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U67 ( .A1(SlicesFromChi[192]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n280) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n277), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n276), .A(
        all_mux_linear_7__MUX_theta_state_inst_n275), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[16]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n277), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n275) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U64 ( .A(SlicesFromChi[191]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n276) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U63 ( .A1(SlicesFromChi[191]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n277) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U62 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n274), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n286), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n273), .A(
        all_mux_linear_7__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[15]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U61 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n274), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n286), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n272) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U60 ( .A(SlicesFromChi[190]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n273) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n270), .B(
        all_mux_linear_7__MUX_theta_state_inst_n269), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n323) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n268), .B(
        all_mux_linear_7__MUX_theta_state_inst_n267), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n269) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U57 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n266), .B(
        all_mux_linear_7__MUX_theta_state_inst_n265), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n268) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U56 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n264), .B(
        all_mux_linear_7__MUX_theta_state_inst_n263), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n270) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U55 ( .A1(SlicesFromChi[190]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n274) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n267), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n261), .A(
        all_mux_linear_7__MUX_theta_state_inst_n260), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[14]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n267), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n260) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U52 ( .A(SlicesFromChi[189]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n261) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U51 ( .A1(SlicesFromChi[189]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n267) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U50 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n259), .A(
        all_mux_linear_7__MUX_theta_state_inst_n258), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[13]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U49 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n265), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n258) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U48 ( .A(SlicesFromChi[188]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n259) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U47 ( .A1(SlicesFromChi[188]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n265) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U46 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n266), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n257), .A(
        all_mux_linear_7__MUX_theta_state_inst_n256), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[12]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U45 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n266), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n256) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U44 ( .A(SlicesFromChi[187]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n257) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U43 ( .A1(SlicesFromChi[187]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n266) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U42 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n263), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n231), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n255), .A(
        all_mux_linear_7__MUX_theta_state_inst_n254), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[11]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U41 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n263), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n254) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U40 ( .A(SlicesFromChi[186]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n255) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U39 ( .A1(SlicesFromChi[186]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n263) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U38 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n264), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n262), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n253), .A(
        all_mux_linear_7__MUX_theta_state_inst_n252), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[10]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U37 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n264), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n262), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n252) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U36 ( .A(SlicesFromChi[185]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n253) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n250), .B(
        all_mux_linear_7__MUX_theta_state_inst_n249), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n296) );
  OAI211_X1 all_mux_linear_7__MUX_theta_state_inst_U34 ( .C1(
        SlicesFromChi[190]), .C2(all_mux_linear_7__MUX_theta_state_inst_n248), 
        .A(all_mux_linear_7__MUX_theta_state_inst_n233), .B(
        all_mux_linear_7__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n249) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U33 ( .A1(SlicesFromChi[190]), .A2(all_mux_linear_7__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n247) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U32 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n279), .B(SlicesFromChi[193]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n248) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U31 ( .A(SlicesFromChi[192]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n279) );
  OAI211_X1 all_mux_linear_7__MUX_theta_state_inst_U30 ( .C1(
        SlicesFromChi[191]), .C2(SlicesFromChi[194]), .A(
        all_mux_linear_7__MUX_theta_state_inst_n232), .B(
        all_mux_linear_7__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n250) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[194]), .A2(SlicesFromChi[191]), .ZN(all_mux_linear_7__MUX_theta_state_inst_n246) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U28 ( .A1(SlicesFromChi[185]), .A2(all_mux_linear_7__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n264) );
  OAI221_X1 all_mux_linear_7__MUX_theta_state_inst_U27 ( .B1(
        all_mux_linear_7__MUX_theta_state_inst_n293), .B2(
        all_mux_linear_7__MUX_theta_state_inst_n321), .C1(
        all_mux_linear_7__MUX_theta_state_inst_n230), .C2(
        all_mux_linear_7__MUX_theta_state_inst_n245), .A(
        all_mux_linear_7__MUX_theta_state_inst_n244), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[0]) );
  NAND3_X1 all_mux_linear_7__MUX_theta_state_inst_U26 ( .A1(
        all_mux_linear_7__MUX_theta_state_inst_n293), .A2(
        all_mux_linear_7__MUX_theta_state_inst_n321), .A3(
        all_mux_linear_7__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n244) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U25 ( .A(SlicesFromChi[175]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n245) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n243), .B(
        all_mux_linear_7__MUX_theta_state_inst_n242), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n251) );
  AOI211_X1 all_mux_linear_7__MUX_theta_state_inst_U23 ( .C1(
        SlicesFromChi[181]), .C2(SlicesFromChi[182]), .A(Reset), .B(
        all_mux_linear_7__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n242) );
  NOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U22 ( .A1(SlicesFromChi[181]), 
        .A2(SlicesFromChi[182]), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n241) );
  OAI211_X1 all_mux_linear_7__MUX_theta_state_inst_U21 ( .C1(
        SlicesFromChi[180]), .C2(all_mux_linear_7__MUX_theta_state_inst_n240), 
        .A(all_mux_linear_7__MUX_theta_state_inst_n232), .B(
        all_mux_linear_7__MUX_theta_state_inst_n239), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n243) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U20 ( .A1(SlicesFromChi[180]), .A2(all_mux_linear_7__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n239) );
  XOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U19 ( .A(SlicesFromChi[184]), 
        .B(SlicesFromChi[183]), .Z(all_mux_linear_7__MUX_theta_state_inst_n240) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U18 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n238), .B(
        all_mux_linear_7__MUX_theta_state_inst_n237), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n271) );
  AOI211_X1 all_mux_linear_7__MUX_theta_state_inst_U17 ( .C1(
        SlicesFromChi[196]), .C2(SlicesFromChi[199]), .A(Reset), .B(
        all_mux_linear_7__MUX_theta_state_inst_n236), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n237) );
  NOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U16 ( .A1(SlicesFromChi[196]), 
        .A2(SlicesFromChi[199]), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n236) );
  OAI211_X1 all_mux_linear_7__MUX_theta_state_inst_U15 ( .C1(
        SlicesFromChi[195]), .C2(all_mux_linear_7__MUX_theta_state_inst_n235), 
        .A(all_mux_linear_7__MUX_theta_state_inst_n232), .B(
        all_mux_linear_7__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n238) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U14 ( .A1(SlicesFromChi[195]), .A2(all_mux_linear_7__MUX_theta_state_inst_n235), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n234) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U13 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n304), .B(SlicesFromChi[198]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n235) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U12 ( .A(SlicesFromChi[197]), 
        .ZN(all_mux_linear_7__MUX_theta_state_inst_n304) );
  NAND2_X1 all_mux_linear_7__MUX_theta_state_inst_U11 ( .A1(SlicesFromChi[175]), .A2(all_mux_linear_7__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n293) );
  XOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U10 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n271), .B(
        all_mux_linear_7__MUX_theta_state_inst_n251), .Z(
        all_mux_linear_7__MUX_theta_state_inst_n321) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U9 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n271), .B(
        all_mux_linear_7__MUX_theta_state_inst_n323), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n286) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U8 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n251), .B(
        all_mux_linear_7__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n262) );
  XNOR2_X1 all_mux_linear_7__MUX_theta_state_inst_U7 ( .A(
        all_mux_linear_7__MUX_theta_state_inst_n324), .B(
        all_mux_linear_7__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n311) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U6 ( .A(Reset), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U5 ( .A(n4), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n230) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U4 ( .A(n4), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n231) );
  INV_X1 all_mux_linear_7__MUX_theta_state_inst_U3 ( .A(Reset), .ZN(
        all_mux_linear_7__MUX_theta_state_inst_n233) );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[175]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[176]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[177]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[178]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[179]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[180]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[181]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[182]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[183]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[184]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[185]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[186]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[187]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[188]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[189]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[190]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[191]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[192]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[193]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[194]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[195]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[196]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[197]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[198]), .QN() );
  DFF_X1 all_mux_linear_7__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_7__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[199]), .QN() );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U116 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n318), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n317), .A(
        all_mux_linear_8__MUX_theta_state_inst_n316), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[9]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U115 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[209]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n318), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n316) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U114 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n317), .A(
        all_mux_linear_8__MUX_theta_state_inst_n313), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[8]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U113 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[208]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n314), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n313) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U112 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n312), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n317), .A(
        all_mux_linear_8__MUX_theta_state_inst_n311), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[7]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U111 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[207]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n312), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n311) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U110 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n310), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n317), .A(
        all_mux_linear_8__MUX_theta_state_inst_n309), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[6]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U109 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[206]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n310), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n309) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U108 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n308), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n317), .A(
        all_mux_linear_8__MUX_theta_state_inst_n307), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[5]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U107 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[205]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n308), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n315), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n307) );
  NOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U106 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(
        all_mux_linear_8__MUX_theta_state_inst_n306), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n315) );
  NAND2_X1 all_mux_linear_8__MUX_theta_state_inst_U105 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_8__MUX_theta_state_inst_n306), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n317) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U104 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n305), .B(
        all_mux_linear_8__MUX_theta_state_inst_n304), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n306) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U103 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n303), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n302), .A(
        all_mux_linear_8__MUX_theta_state_inst_n301), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[4]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U102 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[204]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n303), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n301) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U101 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n299), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n302), .A(
        all_mux_linear_8__MUX_theta_state_inst_n298), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[3]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U100 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[203]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n299), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n298) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U99 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n297), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n302), .A(
        all_mux_linear_8__MUX_theta_state_inst_n296), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[2]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U98 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[202]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n297), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n296) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U97 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n295), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n294), .A(
        all_mux_linear_8__MUX_theta_state_inst_n293), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[24]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U96 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[224]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n295), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n293) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U95 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n294), .A(
        all_mux_linear_8__MUX_theta_state_inst_n290), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[23]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U94 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[223]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n291), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n290) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U93 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n289), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n294), .A(
        all_mux_linear_8__MUX_theta_state_inst_n288), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[22]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U92 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[222]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n289), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n288) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U91 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n287), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n294), .A(
        all_mux_linear_8__MUX_theta_state_inst_n286), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[21]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U90 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[221]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n287), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n286) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U89 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n285), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n294), .A(
        all_mux_linear_8__MUX_theta_state_inst_n284), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[20]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U88 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[220]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n285), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n292), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n284) );
  NOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U87 ( .A1(n4), .A2(
        all_mux_linear_8__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n292) );
  NAND2_X1 all_mux_linear_8__MUX_theta_state_inst_U86 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_8__MUX_theta_state_inst_n283), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n294) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U85 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n282), .B(
        all_mux_linear_8__MUX_theta_state_inst_n304), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n283) );
  XOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U84 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n281), .B(
        all_mux_linear_8__MUX_theta_state_inst_n280), .Z(
        all_mux_linear_8__MUX_theta_state_inst_n304) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U83 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n279), .B(
        all_mux_linear_8__MUX_theta_state_inst_n278), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n280) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U82 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n277), .B(
        all_mux_linear_8__MUX_theta_state_inst_n303), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n278) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U81 ( .A1(Reset), .A2(
        InData[54]), .B1(SlicesFromChi[204]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n303) );
  XOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U80 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n299), .B(
        all_mux_linear_8__MUX_theta_state_inst_n297), .Z(
        all_mux_linear_8__MUX_theta_state_inst_n279) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U79 ( .A1(Reset), .A2(
        InData[52]), .B1(SlicesFromChi[202]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n297) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U78 ( .A1(Reset), .A2(
        InData[53]), .B1(SlicesFromChi[203]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n299) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U77 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n277), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n302), .A(
        all_mux_linear_8__MUX_theta_state_inst_n276), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[1]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U76 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[201]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n300), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n277), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n276) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U75 ( .A1(Reset), .A2(
        InData[51]), .B1(SlicesFromChi[201]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n277) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U74 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n275), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n274), .A(
        all_mux_linear_8__MUX_theta_state_inst_n273), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[19]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U73 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[219]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n275), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n273) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U72 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n271), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n274), .A(
        all_mux_linear_8__MUX_theta_state_inst_n270), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[18]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U71 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[218]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n271), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n270) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U70 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n269), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n274), .A(
        all_mux_linear_8__MUX_theta_state_inst_n268), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[17]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U69 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[217]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n269), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n268) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U68 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n267), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n274), .A(
        all_mux_linear_8__MUX_theta_state_inst_n266), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[16]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U67 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[216]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n267), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n266) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U66 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n274), .A(
        all_mux_linear_8__MUX_theta_state_inst_n264), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[15]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U65 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[215]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n265), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n272), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n264) );
  NOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U64 ( .A1(n4), .A2(
        all_mux_linear_8__MUX_theta_state_inst_n263), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n272) );
  NAND2_X1 all_mux_linear_8__MUX_theta_state_inst_U63 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_8__MUX_theta_state_inst_n263), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n274) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U62 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n262), .B(
        all_mux_linear_8__MUX_theta_state_inst_n305), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n263) );
  XOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U61 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n261), .B(
        all_mux_linear_8__MUX_theta_state_inst_n260), .Z(
        all_mux_linear_8__MUX_theta_state_inst_n305) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U60 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n259), .B(
        all_mux_linear_8__MUX_theta_state_inst_n258), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n260) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U59 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n257), .B(
        all_mux_linear_8__MUX_theta_state_inst_n256), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n258) );
  XOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U58 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n255), .B(
        all_mux_linear_8__MUX_theta_state_inst_n254), .Z(
        all_mux_linear_8__MUX_theta_state_inst_n259) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U57 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n255), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n253), .A(
        all_mux_linear_8__MUX_theta_state_inst_n252), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[14]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U56 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[214]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n255), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n252) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U55 ( .A1(Reset), .A2(
        InData[64]), .B1(SlicesFromChi[214]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n255) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U54 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n254), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n253), .A(
        all_mux_linear_8__MUX_theta_state_inst_n250), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[13]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U53 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[213]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n254), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n250) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U52 ( .A1(Reset), .A2(
        InData[63]), .B1(SlicesFromChi[213]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n254) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U51 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n256), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n253), .A(
        all_mux_linear_8__MUX_theta_state_inst_n249), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[12]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U50 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[212]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n256), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n249) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U49 ( .A1(Reset), .A2(
        InData[62]), .B1(SlicesFromChi[212]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n256) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U48 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n257), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n253), .A(
        all_mux_linear_8__MUX_theta_state_inst_n248), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[11]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U47 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[211]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n251), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n257), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n248) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U46 ( .A1(Reset), .A2(
        InData[61]), .B1(SlicesFromChi[211]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n257) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U45 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n261), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n253), .A(
        all_mux_linear_8__MUX_theta_state_inst_n247), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[10]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U44 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n230), .A2(SlicesFromChi[210]), 
        .B1(all_mux_linear_8__MUX_theta_state_inst_n261), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n251), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n247) );
  NOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U43 ( .A1(n4), .A2(
        all_mux_linear_8__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n251) );
  NAND2_X1 all_mux_linear_8__MUX_theta_state_inst_U42 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_8__MUX_theta_state_inst_n246), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n253) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U41 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n245), .B(
        all_mux_linear_8__MUX_theta_state_inst_n282), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n246) );
  XOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U40 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n275), .B(
        all_mux_linear_8__MUX_theta_state_inst_n244), .Z(
        all_mux_linear_8__MUX_theta_state_inst_n282) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U39 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n243), .B(
        all_mux_linear_8__MUX_theta_state_inst_n242), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n244) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U38 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n267), .B(
        all_mux_linear_8__MUX_theta_state_inst_n265), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n242) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U37 ( .A1(Reset), .A2(
        InData[65]), .B1(SlicesFromChi[215]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n265) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U36 ( .A1(Reset), .A2(
        InData[66]), .B1(SlicesFromChi[216]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n267) );
  XOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U35 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n271), .B(
        all_mux_linear_8__MUX_theta_state_inst_n269), .Z(
        all_mux_linear_8__MUX_theta_state_inst_n243) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U34 ( .A1(Reset), .A2(
        InData[67]), .B1(SlicesFromChi[217]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n269) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U33 ( .A1(Reset), .A2(
        InData[68]), .B1(SlicesFromChi[218]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n271) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U32 ( .A1(Reset), .A2(
        InData[69]), .B1(SlicesFromChi[219]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n232), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n275) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U31 ( .A1(Reset), .A2(
        InData[60]), .B1(SlicesFromChi[210]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n261) );
  OAI21_X1 all_mux_linear_8__MUX_theta_state_inst_U30 ( .B1(
        all_mux_linear_8__MUX_theta_state_inst_n281), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n302), .A(
        all_mux_linear_8__MUX_theta_state_inst_n241), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[0]) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U29 ( .A1(SlicesFromChi[200]), .A2(all_mux_linear_8__MUX_theta_state_inst_n230), .B1(
        all_mux_linear_8__MUX_theta_state_inst_n281), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n300), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n241) );
  NOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U28 ( .A1(n4), .A2(
        all_mux_linear_8__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n300) );
  NAND2_X1 all_mux_linear_8__MUX_theta_state_inst_U27 ( .A1(
        all_mux_linear_8__MUX_theta_state_inst_n231), .A2(
        all_mux_linear_8__MUX_theta_state_inst_n240), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n302) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U26 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n262), .B(
        all_mux_linear_8__MUX_theta_state_inst_n245), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n240) );
  XOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U25 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n312), .B(
        all_mux_linear_8__MUX_theta_state_inst_n239), .Z(
        all_mux_linear_8__MUX_theta_state_inst_n245) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U24 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n238), .B(
        all_mux_linear_8__MUX_theta_state_inst_n237), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n239) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U23 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n310), .B(
        all_mux_linear_8__MUX_theta_state_inst_n308), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n237) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U22 ( .A1(Reset), .A2(
        InData[55]), .B1(SlicesFromChi[205]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n308) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U21 ( .A1(Reset), .A2(
        InData[56]), .B1(SlicesFromChi[206]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n310) );
  XOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U20 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n314), .B(
        all_mux_linear_8__MUX_theta_state_inst_n318), .Z(
        all_mux_linear_8__MUX_theta_state_inst_n238) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U19 ( .A1(Reset), .A2(
        InData[59]), .B1(SlicesFromChi[209]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n318) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U18 ( .A1(Reset), .A2(
        InData[58]), .B1(SlicesFromChi[208]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n314) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U17 ( .A1(Reset), .A2(
        InData[57]), .B1(SlicesFromChi[207]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n312) );
  XOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U16 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n295), .B(
        all_mux_linear_8__MUX_theta_state_inst_n236), .Z(
        all_mux_linear_8__MUX_theta_state_inst_n262) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U15 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n235), .B(
        all_mux_linear_8__MUX_theta_state_inst_n234), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n236) );
  XNOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U14 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n287), .B(
        all_mux_linear_8__MUX_theta_state_inst_n285), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n234) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U13 ( .A1(Reset), .A2(
        InData[70]), .B1(SlicesFromChi[220]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n285) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U12 ( .A1(Reset), .A2(
        InData[71]), .B1(SlicesFromChi[221]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n287) );
  XOR2_X1 all_mux_linear_8__MUX_theta_state_inst_U11 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n291), .B(
        all_mux_linear_8__MUX_theta_state_inst_n289), .Z(
        all_mux_linear_8__MUX_theta_state_inst_n235) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U10 ( .A1(Reset), .A2(
        InData[72]), .B1(SlicesFromChi[222]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n289) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U9 ( .A1(Reset), .A2(
        InData[73]), .B1(SlicesFromChi[223]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n291) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U8 ( .A1(Reset), .A2(
        InData[74]), .B1(SlicesFromChi[224]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n295) );
  AOI22_X1 all_mux_linear_8__MUX_theta_state_inst_U7 ( .A1(Reset), .A2(
        InData[50]), .B1(SlicesFromChi[200]), .B2(
        all_mux_linear_8__MUX_theta_state_inst_n233), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n281) );
  INV_X2 all_mux_linear_8__MUX_theta_state_inst_U6 ( .A(
        all_mux_linear_8__MUX_theta_state_inst_n231), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n230) );
  INV_X1 all_mux_linear_8__MUX_theta_state_inst_U5 ( .A(Reset), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n233) );
  INV_X1 all_mux_linear_8__MUX_theta_state_inst_U4 ( .A(Reset), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n232) );
  INV_X1 all_mux_linear_8__MUX_theta_state_inst_U3 ( .A(n4), .ZN(
        all_mux_linear_8__MUX_theta_state_inst_n231) );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_0_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[0]), .CK(Clock), .Q(
        StateOut[200]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_1_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[1]), .CK(Clock), .Q(
        StateOut[201]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_2_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[2]), .CK(Clock), .Q(
        StateOut[202]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_3_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[3]), .CK(Clock), .Q(
        StateOut[203]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_4_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[4]), .CK(Clock), .Q(
        StateOut[204]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_5_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[5]), .CK(Clock), .Q(
        StateOut[205]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_6_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[6]), .CK(Clock), .Q(
        StateOut[206]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_7_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[7]), .CK(Clock), .Q(
        StateOut[207]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_8_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[8]), .CK(Clock), .Q(
        StateOut[208]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_9_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[9]), .CK(Clock), .Q(
        StateOut[209]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_10_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[10]), .CK(Clock), .Q(
        StateOut[210]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_11_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[11]), .CK(Clock), .Q(
        StateOut[211]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_12_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[12]), .CK(Clock), .Q(
        StateOut[212]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_13_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[13]), .CK(Clock), .Q(
        StateOut[213]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_14_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[14]), .CK(Clock), .Q(
        StateOut[214]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_15_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[15]), .CK(Clock), .Q(
        StateOut[215]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_16_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[16]), .CK(Clock), .Q(
        StateOut[216]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_17_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[17]), .CK(Clock), .Q(
        StateOut[217]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_18_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[18]), .CK(Clock), .Q(
        StateOut[218]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_19_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[19]), .CK(Clock), .Q(
        StateOut[219]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_20_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[20]), .CK(Clock), .Q(
        StateOut[220]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_21_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[21]), .CK(Clock), .Q(
        StateOut[221]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_22_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[22]), .CK(Clock), .Q(
        StateOut[222]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_23_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[23]), .CK(Clock), .Q(
        StateOut[223]), .QN() );
  DFF_X1 all_mux_linear_8__MUX_theta_state_inst_StatexDP_reg_24_ ( .D(
        all_mux_linear_8__MUX_theta_state_inst_StateIn[24]), .CK(Clock), .Q(
        StateOut[224]), .QN() );
  XNOR2_X1 COMPRESSION_BITS_0__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_0__BIT_SHARES_0__Copression_n3), .B(StateOut[50]), 
        .ZN(OutData[0]) );
  XNOR2_X1 COMPRESSION_BITS_0__BIT_SHARES_0__Copression_U1 ( .A(StateOut[0]), 
        .B(StateOut[25]), .ZN(COMPRESSION_BITS_0__BIT_SHARES_0__Copression_n3)
         );
  XNOR2_X1 COMPRESSION_BITS_0__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_0__BIT_SHARES_1__Copression_n3), .B(StateOut[125]), 
        .ZN(OutData[25]) );
  XNOR2_X1 COMPRESSION_BITS_0__BIT_SHARES_1__Copression_U1 ( .A(StateOut[75]), 
        .B(StateOut[100]), .ZN(COMPRESSION_BITS_0__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_0__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_0__BIT_SHARES_2__Copression_n3), .B(StateOut[200]), 
        .ZN(OutData[50]) );
  XNOR2_X1 COMPRESSION_BITS_0__BIT_SHARES_2__Copression_U1 ( .A(StateOut[150]), 
        .B(StateOut[175]), .ZN(COMPRESSION_BITS_0__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_1__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_1__BIT_SHARES_0__Copression_n3), .B(StateOut[51]), 
        .ZN(OutData[1]) );
  XNOR2_X1 COMPRESSION_BITS_1__BIT_SHARES_0__Copression_U1 ( .A(StateOut[1]), 
        .B(StateOut[26]), .ZN(COMPRESSION_BITS_1__BIT_SHARES_0__Copression_n3)
         );
  XNOR2_X1 COMPRESSION_BITS_1__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_1__BIT_SHARES_1__Copression_n3), .B(StateOut[126]), 
        .ZN(OutData[26]) );
  XNOR2_X1 COMPRESSION_BITS_1__BIT_SHARES_1__Copression_U1 ( .A(StateOut[76]), 
        .B(StateOut[101]), .ZN(COMPRESSION_BITS_1__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_1__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_1__BIT_SHARES_2__Copression_n3), .B(StateOut[201]), 
        .ZN(OutData[51]) );
  XNOR2_X1 COMPRESSION_BITS_1__BIT_SHARES_2__Copression_U1 ( .A(StateOut[151]), 
        .B(StateOut[176]), .ZN(COMPRESSION_BITS_1__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_2__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_2__BIT_SHARES_0__Copression_n3), .B(StateOut[52]), 
        .ZN(OutData[2]) );
  XNOR2_X1 COMPRESSION_BITS_2__BIT_SHARES_0__Copression_U1 ( .A(StateOut[2]), 
        .B(StateOut[27]), .ZN(COMPRESSION_BITS_2__BIT_SHARES_0__Copression_n3)
         );
  XNOR2_X1 COMPRESSION_BITS_2__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_2__BIT_SHARES_1__Copression_n3), .B(StateOut[127]), 
        .ZN(OutData[27]) );
  XNOR2_X1 COMPRESSION_BITS_2__BIT_SHARES_1__Copression_U1 ( .A(StateOut[77]), 
        .B(StateOut[102]), .ZN(COMPRESSION_BITS_2__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_2__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_2__BIT_SHARES_2__Copression_n3), .B(StateOut[202]), 
        .ZN(OutData[52]) );
  XNOR2_X1 COMPRESSION_BITS_2__BIT_SHARES_2__Copression_U1 ( .A(StateOut[152]), 
        .B(StateOut[177]), .ZN(COMPRESSION_BITS_2__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_3__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_3__BIT_SHARES_0__Copression_n3), .B(StateOut[53]), 
        .ZN(OutData[3]) );
  XNOR2_X1 COMPRESSION_BITS_3__BIT_SHARES_0__Copression_U1 ( .A(StateOut[3]), 
        .B(StateOut[28]), .ZN(COMPRESSION_BITS_3__BIT_SHARES_0__Copression_n3)
         );
  XNOR2_X1 COMPRESSION_BITS_3__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_3__BIT_SHARES_1__Copression_n3), .B(StateOut[128]), 
        .ZN(OutData[28]) );
  XNOR2_X1 COMPRESSION_BITS_3__BIT_SHARES_1__Copression_U1 ( .A(StateOut[78]), 
        .B(StateOut[103]), .ZN(COMPRESSION_BITS_3__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_3__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_3__BIT_SHARES_2__Copression_n3), .B(StateOut[203]), 
        .ZN(OutData[53]) );
  XNOR2_X1 COMPRESSION_BITS_3__BIT_SHARES_2__Copression_U1 ( .A(StateOut[153]), 
        .B(StateOut[178]), .ZN(COMPRESSION_BITS_3__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_4__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_4__BIT_SHARES_0__Copression_n3), .B(StateOut[54]), 
        .ZN(OutData[4]) );
  XNOR2_X1 COMPRESSION_BITS_4__BIT_SHARES_0__Copression_U1 ( .A(StateOut[4]), 
        .B(StateOut[29]), .ZN(COMPRESSION_BITS_4__BIT_SHARES_0__Copression_n3)
         );
  XNOR2_X1 COMPRESSION_BITS_4__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_4__BIT_SHARES_1__Copression_n3), .B(StateOut[129]), 
        .ZN(OutData[29]) );
  XNOR2_X1 COMPRESSION_BITS_4__BIT_SHARES_1__Copression_U1 ( .A(StateOut[79]), 
        .B(StateOut[104]), .ZN(COMPRESSION_BITS_4__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_4__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_4__BIT_SHARES_2__Copression_n3), .B(StateOut[204]), 
        .ZN(OutData[54]) );
  XNOR2_X1 COMPRESSION_BITS_4__BIT_SHARES_2__Copression_U1 ( .A(StateOut[154]), 
        .B(StateOut[179]), .ZN(COMPRESSION_BITS_4__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_5__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_5__BIT_SHARES_0__Copression_n3), .B(StateOut[55]), 
        .ZN(OutData[5]) );
  XNOR2_X1 COMPRESSION_BITS_5__BIT_SHARES_0__Copression_U1 ( .A(StateOut[5]), 
        .B(StateOut[30]), .ZN(COMPRESSION_BITS_5__BIT_SHARES_0__Copression_n3)
         );
  XNOR2_X1 COMPRESSION_BITS_5__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_5__BIT_SHARES_1__Copression_n3), .B(StateOut[130]), 
        .ZN(OutData[30]) );
  XNOR2_X1 COMPRESSION_BITS_5__BIT_SHARES_1__Copression_U1 ( .A(StateOut[80]), 
        .B(StateOut[105]), .ZN(COMPRESSION_BITS_5__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_5__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_5__BIT_SHARES_2__Copression_n3), .B(StateOut[205]), 
        .ZN(OutData[55]) );
  XNOR2_X1 COMPRESSION_BITS_5__BIT_SHARES_2__Copression_U1 ( .A(StateOut[155]), 
        .B(StateOut[180]), .ZN(COMPRESSION_BITS_5__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_6__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_6__BIT_SHARES_0__Copression_n3), .B(StateOut[56]), 
        .ZN(OutData[6]) );
  XNOR2_X1 COMPRESSION_BITS_6__BIT_SHARES_0__Copression_U1 ( .A(StateOut[6]), 
        .B(StateOut[31]), .ZN(COMPRESSION_BITS_6__BIT_SHARES_0__Copression_n3)
         );
  XNOR2_X1 COMPRESSION_BITS_6__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_6__BIT_SHARES_1__Copression_n3), .B(StateOut[131]), 
        .ZN(OutData[31]) );
  XNOR2_X1 COMPRESSION_BITS_6__BIT_SHARES_1__Copression_U1 ( .A(StateOut[81]), 
        .B(StateOut[106]), .ZN(COMPRESSION_BITS_6__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_6__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_6__BIT_SHARES_2__Copression_n3), .B(StateOut[206]), 
        .ZN(OutData[56]) );
  XNOR2_X1 COMPRESSION_BITS_6__BIT_SHARES_2__Copression_U1 ( .A(StateOut[156]), 
        .B(StateOut[181]), .ZN(COMPRESSION_BITS_6__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_7__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_7__BIT_SHARES_0__Copression_n3), .B(StateOut[57]), 
        .ZN(OutData[7]) );
  XNOR2_X1 COMPRESSION_BITS_7__BIT_SHARES_0__Copression_U1 ( .A(StateOut[7]), 
        .B(StateOut[32]), .ZN(COMPRESSION_BITS_7__BIT_SHARES_0__Copression_n3)
         );
  XNOR2_X1 COMPRESSION_BITS_7__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_7__BIT_SHARES_1__Copression_n3), .B(StateOut[132]), 
        .ZN(OutData[32]) );
  XNOR2_X1 COMPRESSION_BITS_7__BIT_SHARES_1__Copression_U1 ( .A(StateOut[82]), 
        .B(StateOut[107]), .ZN(COMPRESSION_BITS_7__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_7__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_7__BIT_SHARES_2__Copression_n3), .B(StateOut[207]), 
        .ZN(OutData[57]) );
  XNOR2_X1 COMPRESSION_BITS_7__BIT_SHARES_2__Copression_U1 ( .A(StateOut[157]), 
        .B(StateOut[182]), .ZN(COMPRESSION_BITS_7__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_8__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_8__BIT_SHARES_0__Copression_n3), .B(StateOut[58]), 
        .ZN(OutData[8]) );
  XNOR2_X1 COMPRESSION_BITS_8__BIT_SHARES_0__Copression_U1 ( .A(StateOut[8]), 
        .B(StateOut[33]), .ZN(COMPRESSION_BITS_8__BIT_SHARES_0__Copression_n3)
         );
  XNOR2_X1 COMPRESSION_BITS_8__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_8__BIT_SHARES_1__Copression_n3), .B(StateOut[133]), 
        .ZN(OutData[33]) );
  XNOR2_X1 COMPRESSION_BITS_8__BIT_SHARES_1__Copression_U1 ( .A(StateOut[83]), 
        .B(StateOut[108]), .ZN(COMPRESSION_BITS_8__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_8__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_8__BIT_SHARES_2__Copression_n3), .B(StateOut[208]), 
        .ZN(OutData[58]) );
  XNOR2_X1 COMPRESSION_BITS_8__BIT_SHARES_2__Copression_U1 ( .A(StateOut[158]), 
        .B(StateOut[183]), .ZN(COMPRESSION_BITS_8__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_9__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_9__BIT_SHARES_0__Copression_n3), .B(StateOut[59]), 
        .ZN(OutData[9]) );
  XNOR2_X1 COMPRESSION_BITS_9__BIT_SHARES_0__Copression_U1 ( .A(StateOut[9]), 
        .B(StateOut[34]), .ZN(COMPRESSION_BITS_9__BIT_SHARES_0__Copression_n3)
         );
  XNOR2_X1 COMPRESSION_BITS_9__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_9__BIT_SHARES_1__Copression_n3), .B(StateOut[134]), 
        .ZN(OutData[34]) );
  XNOR2_X1 COMPRESSION_BITS_9__BIT_SHARES_1__Copression_U1 ( .A(StateOut[84]), 
        .B(StateOut[109]), .ZN(COMPRESSION_BITS_9__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_9__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_9__BIT_SHARES_2__Copression_n3), .B(StateOut[209]), 
        .ZN(OutData[59]) );
  XNOR2_X1 COMPRESSION_BITS_9__BIT_SHARES_2__Copression_U1 ( .A(StateOut[159]), 
        .B(StateOut[184]), .ZN(COMPRESSION_BITS_9__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_10__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_10__BIT_SHARES_0__Copression_n3), .B(StateOut[60]), 
        .ZN(OutData[10]) );
  XNOR2_X1 COMPRESSION_BITS_10__BIT_SHARES_0__Copression_U1 ( .A(StateOut[10]), 
        .B(StateOut[35]), .ZN(COMPRESSION_BITS_10__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_10__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_10__BIT_SHARES_1__Copression_n3), .B(StateOut[135]), 
        .ZN(OutData[35]) );
  XNOR2_X1 COMPRESSION_BITS_10__BIT_SHARES_1__Copression_U1 ( .A(StateOut[85]), 
        .B(StateOut[110]), .ZN(
        COMPRESSION_BITS_10__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_10__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_10__BIT_SHARES_2__Copression_n3), .B(StateOut[210]), 
        .ZN(OutData[60]) );
  XNOR2_X1 COMPRESSION_BITS_10__BIT_SHARES_2__Copression_U1 ( .A(StateOut[160]), .B(StateOut[185]), .ZN(COMPRESSION_BITS_10__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_11__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_11__BIT_SHARES_0__Copression_n3), .B(StateOut[61]), 
        .ZN(OutData[11]) );
  XNOR2_X1 COMPRESSION_BITS_11__BIT_SHARES_0__Copression_U1 ( .A(StateOut[11]), 
        .B(StateOut[36]), .ZN(COMPRESSION_BITS_11__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_11__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_11__BIT_SHARES_1__Copression_n3), .B(StateOut[136]), 
        .ZN(OutData[36]) );
  XNOR2_X1 COMPRESSION_BITS_11__BIT_SHARES_1__Copression_U1 ( .A(StateOut[86]), 
        .B(StateOut[111]), .ZN(
        COMPRESSION_BITS_11__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_11__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_11__BIT_SHARES_2__Copression_n3), .B(StateOut[211]), 
        .ZN(OutData[61]) );
  XNOR2_X1 COMPRESSION_BITS_11__BIT_SHARES_2__Copression_U1 ( .A(StateOut[161]), .B(StateOut[186]), .ZN(COMPRESSION_BITS_11__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_12__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_12__BIT_SHARES_0__Copression_n3), .B(StateOut[62]), 
        .ZN(OutData[12]) );
  XNOR2_X1 COMPRESSION_BITS_12__BIT_SHARES_0__Copression_U1 ( .A(StateOut[12]), 
        .B(StateOut[37]), .ZN(COMPRESSION_BITS_12__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_12__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_12__BIT_SHARES_1__Copression_n3), .B(StateOut[137]), 
        .ZN(OutData[37]) );
  XNOR2_X1 COMPRESSION_BITS_12__BIT_SHARES_1__Copression_U1 ( .A(StateOut[87]), 
        .B(StateOut[112]), .ZN(
        COMPRESSION_BITS_12__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_12__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_12__BIT_SHARES_2__Copression_n3), .B(StateOut[212]), 
        .ZN(OutData[62]) );
  XNOR2_X1 COMPRESSION_BITS_12__BIT_SHARES_2__Copression_U1 ( .A(StateOut[162]), .B(StateOut[187]), .ZN(COMPRESSION_BITS_12__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_13__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_13__BIT_SHARES_0__Copression_n3), .B(StateOut[63]), 
        .ZN(OutData[13]) );
  XNOR2_X1 COMPRESSION_BITS_13__BIT_SHARES_0__Copression_U1 ( .A(StateOut[13]), 
        .B(StateOut[38]), .ZN(COMPRESSION_BITS_13__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_13__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_13__BIT_SHARES_1__Copression_n3), .B(StateOut[138]), 
        .ZN(OutData[38]) );
  XNOR2_X1 COMPRESSION_BITS_13__BIT_SHARES_1__Copression_U1 ( .A(StateOut[88]), 
        .B(StateOut[113]), .ZN(
        COMPRESSION_BITS_13__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_13__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_13__BIT_SHARES_2__Copression_n3), .B(StateOut[213]), 
        .ZN(OutData[63]) );
  XNOR2_X1 COMPRESSION_BITS_13__BIT_SHARES_2__Copression_U1 ( .A(StateOut[163]), .B(StateOut[188]), .ZN(COMPRESSION_BITS_13__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_14__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_14__BIT_SHARES_0__Copression_n3), .B(StateOut[64]), 
        .ZN(OutData[14]) );
  XNOR2_X1 COMPRESSION_BITS_14__BIT_SHARES_0__Copression_U1 ( .A(StateOut[14]), 
        .B(StateOut[39]), .ZN(COMPRESSION_BITS_14__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_14__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_14__BIT_SHARES_1__Copression_n3), .B(StateOut[139]), 
        .ZN(OutData[39]) );
  XNOR2_X1 COMPRESSION_BITS_14__BIT_SHARES_1__Copression_U1 ( .A(StateOut[89]), 
        .B(StateOut[114]), .ZN(
        COMPRESSION_BITS_14__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_14__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_14__BIT_SHARES_2__Copression_n3), .B(StateOut[214]), 
        .ZN(OutData[64]) );
  XNOR2_X1 COMPRESSION_BITS_14__BIT_SHARES_2__Copression_U1 ( .A(StateOut[164]), .B(StateOut[189]), .ZN(COMPRESSION_BITS_14__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_15__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_15__BIT_SHARES_0__Copression_n3), .B(StateOut[165]), 
        .ZN(OutData[15]) );
  XNOR2_X1 COMPRESSION_BITS_15__BIT_SHARES_0__Copression_U1 ( .A(StateOut[15]), 
        .B(StateOut[90]), .ZN(COMPRESSION_BITS_15__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_15__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_15__BIT_SHARES_1__Copression_n3), .B(StateOut[190]), 
        .ZN(OutData[40]) );
  XNOR2_X1 COMPRESSION_BITS_15__BIT_SHARES_1__Copression_U1 ( .A(StateOut[40]), 
        .B(StateOut[115]), .ZN(
        COMPRESSION_BITS_15__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_15__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_15__BIT_SHARES_2__Copression_n3), .B(StateOut[215]), 
        .ZN(OutData[65]) );
  XNOR2_X1 COMPRESSION_BITS_15__BIT_SHARES_2__Copression_U1 ( .A(StateOut[65]), 
        .B(StateOut[140]), .ZN(
        COMPRESSION_BITS_15__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_16__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_16__BIT_SHARES_0__Copression_n3), .B(StateOut[166]), 
        .ZN(OutData[16]) );
  XNOR2_X1 COMPRESSION_BITS_16__BIT_SHARES_0__Copression_U1 ( .A(StateOut[16]), 
        .B(StateOut[91]), .ZN(COMPRESSION_BITS_16__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_16__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_16__BIT_SHARES_1__Copression_n3), .B(StateOut[191]), 
        .ZN(OutData[41]) );
  XNOR2_X1 COMPRESSION_BITS_16__BIT_SHARES_1__Copression_U1 ( .A(StateOut[41]), 
        .B(StateOut[116]), .ZN(
        COMPRESSION_BITS_16__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_16__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_16__BIT_SHARES_2__Copression_n3), .B(StateOut[216]), 
        .ZN(OutData[66]) );
  XNOR2_X1 COMPRESSION_BITS_16__BIT_SHARES_2__Copression_U1 ( .A(StateOut[66]), 
        .B(StateOut[141]), .ZN(
        COMPRESSION_BITS_16__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_17__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_17__BIT_SHARES_0__Copression_n3), .B(StateOut[167]), 
        .ZN(OutData[17]) );
  XNOR2_X1 COMPRESSION_BITS_17__BIT_SHARES_0__Copression_U1 ( .A(StateOut[17]), 
        .B(StateOut[92]), .ZN(COMPRESSION_BITS_17__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_17__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_17__BIT_SHARES_1__Copression_n3), .B(StateOut[192]), 
        .ZN(OutData[42]) );
  XNOR2_X1 COMPRESSION_BITS_17__BIT_SHARES_1__Copression_U1 ( .A(StateOut[42]), 
        .B(StateOut[117]), .ZN(
        COMPRESSION_BITS_17__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_17__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_17__BIT_SHARES_2__Copression_n3), .B(StateOut[217]), 
        .ZN(OutData[67]) );
  XNOR2_X1 COMPRESSION_BITS_17__BIT_SHARES_2__Copression_U1 ( .A(StateOut[67]), 
        .B(StateOut[142]), .ZN(
        COMPRESSION_BITS_17__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_18__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_18__BIT_SHARES_0__Copression_n3), .B(StateOut[168]), 
        .ZN(OutData[18]) );
  XNOR2_X1 COMPRESSION_BITS_18__BIT_SHARES_0__Copression_U1 ( .A(StateOut[18]), 
        .B(StateOut[93]), .ZN(COMPRESSION_BITS_18__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_18__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_18__BIT_SHARES_1__Copression_n3), .B(StateOut[193]), 
        .ZN(OutData[43]) );
  XNOR2_X1 COMPRESSION_BITS_18__BIT_SHARES_1__Copression_U1 ( .A(StateOut[43]), 
        .B(StateOut[118]), .ZN(
        COMPRESSION_BITS_18__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_18__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_18__BIT_SHARES_2__Copression_n3), .B(StateOut[218]), 
        .ZN(OutData[68]) );
  XNOR2_X1 COMPRESSION_BITS_18__BIT_SHARES_2__Copression_U1 ( .A(StateOut[68]), 
        .B(StateOut[143]), .ZN(
        COMPRESSION_BITS_18__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_19__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_19__BIT_SHARES_0__Copression_n3), .B(StateOut[169]), 
        .ZN(OutData[19]) );
  XNOR2_X1 COMPRESSION_BITS_19__BIT_SHARES_0__Copression_U1 ( .A(StateOut[19]), 
        .B(StateOut[94]), .ZN(COMPRESSION_BITS_19__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_19__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_19__BIT_SHARES_1__Copression_n3), .B(StateOut[194]), 
        .ZN(OutData[44]) );
  XNOR2_X1 COMPRESSION_BITS_19__BIT_SHARES_1__Copression_U1 ( .A(StateOut[44]), 
        .B(StateOut[119]), .ZN(
        COMPRESSION_BITS_19__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_19__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_19__BIT_SHARES_2__Copression_n3), .B(StateOut[219]), 
        .ZN(OutData[69]) );
  XNOR2_X1 COMPRESSION_BITS_19__BIT_SHARES_2__Copression_U1 ( .A(StateOut[69]), 
        .B(StateOut[144]), .ZN(
        COMPRESSION_BITS_19__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_20__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_20__BIT_SHARES_0__Copression_n3), .B(StateOut[70]), 
        .ZN(OutData[20]) );
  XNOR2_X1 COMPRESSION_BITS_20__BIT_SHARES_0__Copression_U1 ( .A(StateOut[20]), 
        .B(StateOut[45]), .ZN(COMPRESSION_BITS_20__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_20__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_20__BIT_SHARES_1__Copression_n3), .B(StateOut[145]), 
        .ZN(OutData[45]) );
  XNOR2_X1 COMPRESSION_BITS_20__BIT_SHARES_1__Copression_U1 ( .A(StateOut[95]), 
        .B(StateOut[120]), .ZN(
        COMPRESSION_BITS_20__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_20__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_20__BIT_SHARES_2__Copression_n3), .B(StateOut[220]), 
        .ZN(OutData[70]) );
  XNOR2_X1 COMPRESSION_BITS_20__BIT_SHARES_2__Copression_U1 ( .A(StateOut[170]), .B(StateOut[195]), .ZN(COMPRESSION_BITS_20__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_21__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_21__BIT_SHARES_0__Copression_n3), .B(StateOut[71]), 
        .ZN(OutData[21]) );
  XNOR2_X1 COMPRESSION_BITS_21__BIT_SHARES_0__Copression_U1 ( .A(StateOut[21]), 
        .B(StateOut[46]), .ZN(COMPRESSION_BITS_21__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_21__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_21__BIT_SHARES_1__Copression_n3), .B(StateOut[146]), 
        .ZN(OutData[46]) );
  XNOR2_X1 COMPRESSION_BITS_21__BIT_SHARES_1__Copression_U1 ( .A(StateOut[96]), 
        .B(StateOut[121]), .ZN(
        COMPRESSION_BITS_21__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_21__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_21__BIT_SHARES_2__Copression_n3), .B(StateOut[221]), 
        .ZN(OutData[71]) );
  XNOR2_X1 COMPRESSION_BITS_21__BIT_SHARES_2__Copression_U1 ( .A(StateOut[171]), .B(StateOut[196]), .ZN(COMPRESSION_BITS_21__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_22__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_22__BIT_SHARES_0__Copression_n3), .B(StateOut[72]), 
        .ZN(OutData[22]) );
  XNOR2_X1 COMPRESSION_BITS_22__BIT_SHARES_0__Copression_U1 ( .A(StateOut[22]), 
        .B(StateOut[47]), .ZN(COMPRESSION_BITS_22__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_22__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_22__BIT_SHARES_1__Copression_n3), .B(StateOut[147]), 
        .ZN(OutData[47]) );
  XNOR2_X1 COMPRESSION_BITS_22__BIT_SHARES_1__Copression_U1 ( .A(StateOut[97]), 
        .B(StateOut[122]), .ZN(
        COMPRESSION_BITS_22__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_22__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_22__BIT_SHARES_2__Copression_n3), .B(StateOut[222]), 
        .ZN(OutData[72]) );
  XNOR2_X1 COMPRESSION_BITS_22__BIT_SHARES_2__Copression_U1 ( .A(StateOut[172]), .B(StateOut[197]), .ZN(COMPRESSION_BITS_22__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_23__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_23__BIT_SHARES_0__Copression_n3), .B(StateOut[73]), 
        .ZN(OutData[23]) );
  XNOR2_X1 COMPRESSION_BITS_23__BIT_SHARES_0__Copression_U1 ( .A(StateOut[23]), 
        .B(StateOut[48]), .ZN(COMPRESSION_BITS_23__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_23__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_23__BIT_SHARES_1__Copression_n3), .B(StateOut[148]), 
        .ZN(OutData[48]) );
  XNOR2_X1 COMPRESSION_BITS_23__BIT_SHARES_1__Copression_U1 ( .A(StateOut[98]), 
        .B(StateOut[123]), .ZN(
        COMPRESSION_BITS_23__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_23__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_23__BIT_SHARES_2__Copression_n3), .B(StateOut[223]), 
        .ZN(OutData[73]) );
  XNOR2_X1 COMPRESSION_BITS_23__BIT_SHARES_2__Copression_U1 ( .A(StateOut[173]), .B(StateOut[198]), .ZN(COMPRESSION_BITS_23__BIT_SHARES_2__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_24__BIT_SHARES_0__Copression_U2 ( .A(
        COMPRESSION_BITS_24__BIT_SHARES_0__Copression_n3), .B(StateOut[74]), 
        .ZN(OutData[24]) );
  XNOR2_X1 COMPRESSION_BITS_24__BIT_SHARES_0__Copression_U1 ( .A(StateOut[24]), 
        .B(StateOut[49]), .ZN(COMPRESSION_BITS_24__BIT_SHARES_0__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_24__BIT_SHARES_1__Copression_U2 ( .A(
        COMPRESSION_BITS_24__BIT_SHARES_1__Copression_n3), .B(StateOut[149]), 
        .ZN(OutData[49]) );
  XNOR2_X1 COMPRESSION_BITS_24__BIT_SHARES_1__Copression_U1 ( .A(StateOut[99]), 
        .B(StateOut[124]), .ZN(
        COMPRESSION_BITS_24__BIT_SHARES_1__Copression_n3) );
  XNOR2_X1 COMPRESSION_BITS_24__BIT_SHARES_2__Copression_U2 ( .A(
        COMPRESSION_BITS_24__BIT_SHARES_2__Copression_n3), .B(StateOut[224]), 
        .ZN(OutData[74]) );
  XNOR2_X1 COMPRESSION_BITS_24__BIT_SHARES_2__Copression_U1 ( .A(StateOut[174]), .B(StateOut[199]), .ZN(COMPRESSION_BITS_24__BIT_SHARES_2__Copression_n3) );
  XOR2_X1 CHI_U1 ( .A(CHI_ChiOut_0_), .B(IotaRC_0_), .Z(SlicesFromChi[0]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(OutData[0]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n3), .ZN(CHI_ChiOut_0_) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[12]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n2), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n3) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(OutData[6]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n2) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A(OutData[6]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[5]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A1(OutData[18]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(OutData[12]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U3 ( 
        .A(OutData[12]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7), .ZN(SlicesFromChi[10]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A1(OutData[24]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A(OutData[18]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A(OutData[18]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[15]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A1(OutData[0]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(OutData[24]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U3 ( 
        .A(OutData[24]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7), .ZN(SlicesFromChi[20]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U2 ( 
        .A1(OutData[6]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A(OutData[0]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U3 ( 
        .A(FreshRand[0]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5), .ZN(SlicesFromChi[25]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A1(OutData[37]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A(OutData[6]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[3]), .ZN(SlicesFromChi[30]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[37]), .A2(OutData[18]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7), .ZN(SlicesFromChi[35]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U3 ( 
        .A1(OutData[49]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(OutData[18]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A(FreshRand[6]), .B(OutData[37]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[25]), .A2(OutData[49]), .ZN(SlicesFromChi[40]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[45]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[25]), .A2(OutData[6]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(FreshRand[12]), .B(OutData[49]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U3 ( 
        .A(FreshRand[1]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5), .ZN(SlicesFromChi[50]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U2 ( 
        .A1(OutData[62]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A(OutData[6]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3), .B(FreshRand[4]), .ZN(SlicesFromChi[55]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[62]), .A2(OutData[18]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7), .ZN(SlicesFromChi[60]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U3 ( 
        .A1(OutData[74]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U2 ( 
        .A(OutData[18]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A(FreshRand[7]), .B(OutData[62]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[50]), .A2(OutData[74]), .ZN(SlicesFromChi[65]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5), .ZN(SlicesFromChi[70]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A1(OutData[50]), .A2(OutData[6]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A(FreshRand[13]), .B(OutData[74]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[75]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[31]), .A2(OutData[12]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[0]), .B(OutData[25]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[80]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[43]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[12]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[3]), .B(OutData[31]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[6]), .ZN(SlicesFromChi[85]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[43]), .A2(OutData[24]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[90]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[25]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[24]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[9]), .B(OutData[43]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[31]), .A2(OutData[25]), .ZN(SlicesFromChi[95]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[37]), .A2(OutData[31]), .ZN(SlicesFromChi[100]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[43]), .A2(OutData[37]), .ZN(SlicesFromChi[105]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[49]), .A2(OutData[43]), .ZN(SlicesFromChi[110]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[11]), .ZN(SlicesFromChi[115]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[49]), .A2(OutData[50]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3), .B(FreshRand[14]), .ZN(SlicesFromChi[120]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A1(OutData[50]), .A2(OutData[31]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3), .B(FreshRand[2]), .ZN(SlicesFromChi[125]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A1(OutData[31]), .A2(OutData[62]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3), .B(FreshRand[5]), .ZN(SlicesFromChi[130]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[62]), .A2(OutData[43]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3), .B(FreshRand[8]), .ZN(SlicesFromChi[135]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A1(OutData[43]), .A2(OutData[74]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3), .B(FreshRand[10]), .ZN(SlicesFromChi[140]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[74]), .A2(OutData[0]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U3 ( 
        .A(FreshRand[12]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5), .ZN(SlicesFromChi[145]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A1(OutData[31]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A(OutData[0]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[150]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[56]), .A2(OutData[12]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[1]), .B(OutData[50]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[155]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[68]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[12]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[4]), .B(OutData[56]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[7]), .ZN(SlicesFromChi[160]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[68]), .A2(OutData[24]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[165]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[50]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[24]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[10]), .B(OutData[68]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[56]), .A2(OutData[50]), .ZN(SlicesFromChi[170]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3), .B(FreshRand[2]), .ZN(SlicesFromChi[175]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[56]), .A2(OutData[37]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[5]), .ZN(SlicesFromChi[180]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[37]), .A2(OutData[68]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3), .B(FreshRand[8]), .ZN(SlicesFromChi[185]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[68]), .A2(OutData[49]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[9]), .ZN(SlicesFromChi[190]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[49]), .A2(OutData[0]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(FreshRand[13]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[195]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[56]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(OutData[0]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A1(OutData[62]), .A2(OutData[56]), .ZN(SlicesFromChi[200]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[68]), .A2(OutData[62]), .ZN(SlicesFromChi[205]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A1(OutData[74]), .A2(OutData[68]), .ZN(SlicesFromChi[210]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3), .B(FreshRand[11]), .ZN(SlicesFromChi[215]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[74]), .A2(OutData[25]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3), .B(FreshRand[14]), .ZN(SlicesFromChi[220]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A1(OutData[25]), .A2(OutData[56]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(OutData[15]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7), .ZN(SlicesFromChi[1]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[2]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(OutData[21]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A(OutData[21]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[6]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A1(OutData[8]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(OutData[2]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U3 ( 
        .A(OutData[2]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7), .ZN(SlicesFromChi[11]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A1(OutData[14]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A(OutData[8]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A(OutData[8]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[16]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A1(OutData[15]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(OutData[14]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U3 ( 
        .A(OutData[14]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7), .ZN(SlicesFromChi[21]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U2 ( 
        .A1(OutData[21]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A(OutData[15]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U3 ( 
        .A(FreshRand[15]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5), .ZN(SlicesFromChi[26]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A1(OutData[27]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A(OutData[21]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[18]), .ZN(SlicesFromChi[31]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[27]), .A2(OutData[8]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7), .ZN(SlicesFromChi[36]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U3 ( 
        .A1(OutData[39]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(OutData[8]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A(FreshRand[21]), .B(OutData[27]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[40]), .A2(OutData[39]), .ZN(SlicesFromChi[41]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[46]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[40]), .A2(OutData[21]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(FreshRand[27]), .B(OutData[39]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U3 ( 
        .A(FreshRand[16]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5), .ZN(SlicesFromChi[51]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U2 ( 
        .A1(OutData[52]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A(OutData[21]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3), .B(FreshRand[19]), .ZN(SlicesFromChi[56]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[52]), .A2(OutData[8]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7), .ZN(SlicesFromChi[61]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U3 ( 
        .A1(OutData[64]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U2 ( 
        .A(OutData[8]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A(FreshRand[22]), .B(OutData[52]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[65]), .A2(OutData[64]), .ZN(SlicesFromChi[66]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5), .ZN(SlicesFromChi[71]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A1(OutData[65]), .A2(OutData[21]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A(FreshRand[28]), .B(OutData[64]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[76]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[46]), .A2(OutData[2]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[15]), .B(OutData[40]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[81]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[33]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[2]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[18]), .B(OutData[46]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[21]), .ZN(SlicesFromChi[86]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[33]), .A2(OutData[14]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[91]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[40]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[14]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[24]), .B(OutData[33]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[46]), .A2(OutData[40]), .ZN(SlicesFromChi[96]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[27]), .A2(OutData[46]), .ZN(SlicesFromChi[101]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[33]), .A2(OutData[27]), .ZN(SlicesFromChi[106]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[39]), .A2(OutData[33]), .ZN(SlicesFromChi[111]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[26]), .ZN(SlicesFromChi[116]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[39]), .A2(OutData[65]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3), .B(FreshRand[29]), .ZN(SlicesFromChi[121]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A1(OutData[65]), .A2(OutData[46]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3), .B(FreshRand[17]), .ZN(SlicesFromChi[126]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A1(OutData[46]), .A2(OutData[52]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3), .B(FreshRand[20]), .ZN(SlicesFromChi[131]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[52]), .A2(OutData[33]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3), .B(FreshRand[23]), .ZN(SlicesFromChi[136]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A1(OutData[33]), .A2(OutData[64]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3), .B(FreshRand[25]), .ZN(SlicesFromChi[141]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[64]), .A2(OutData[15]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U3 ( 
        .A(FreshRand[27]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5), .ZN(SlicesFromChi[146]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A1(OutData[46]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A(OutData[15]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[151]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[71]), .A2(OutData[2]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[16]), .B(OutData[65]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[156]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[58]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[2]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[19]), .B(OutData[71]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[22]), .ZN(SlicesFromChi[161]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[58]), .A2(OutData[14]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[166]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[65]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[14]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[25]), .B(OutData[58]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[71]), .A2(OutData[65]), .ZN(SlicesFromChi[171]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3), .B(FreshRand[17]), .ZN(SlicesFromChi[176]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[71]), .A2(OutData[27]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[20]), .ZN(SlicesFromChi[181]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[27]), .A2(OutData[58]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3), .B(FreshRand[23]), .ZN(SlicesFromChi[186]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[58]), .A2(OutData[39]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[24]), .ZN(SlicesFromChi[191]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[39]), .A2(OutData[15]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(FreshRand[28]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[196]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[71]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(OutData[15]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A1(OutData[52]), .A2(OutData[71]), .ZN(SlicesFromChi[201]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[58]), .A2(OutData[52]), .ZN(SlicesFromChi[206]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A1(OutData[64]), .A2(OutData[58]), .ZN(SlicesFromChi[211]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3), .B(FreshRand[26]), .ZN(SlicesFromChi[216]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[64]), .A2(OutData[40]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3), .B(FreshRand[29]), .ZN(SlicesFromChi[221]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A1(OutData[40]), .A2(OutData[71]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(OutData[5]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7), .ZN(SlicesFromChi[2]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[17]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(OutData[11]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A(OutData[11]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[7]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A1(OutData[23]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(OutData[17]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U3 ( 
        .A(OutData[17]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7), .ZN(SlicesFromChi[12]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A1(OutData[4]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A(OutData[23]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A(OutData[23]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[17]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A1(OutData[5]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(OutData[4]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U3 ( 
        .A(OutData[4]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7), .ZN(SlicesFromChi[22]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U2 ( 
        .A1(OutData[11]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A(OutData[5]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U3 ( 
        .A(FreshRand[30]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5), .ZN(SlicesFromChi[27]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A1(OutData[42]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A(OutData[11]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[33]), .ZN(SlicesFromChi[32]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[42]), .A2(OutData[23]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7), .ZN(SlicesFromChi[37]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U3 ( 
        .A1(OutData[29]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(OutData[23]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A(FreshRand[36]), .B(OutData[42]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[30]), .A2(OutData[29]), .ZN(SlicesFromChi[42]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[47]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[30]), .A2(OutData[11]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(FreshRand[42]), .B(OutData[29]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U3 ( 
        .A(FreshRand[31]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5), .ZN(SlicesFromChi[52]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U2 ( 
        .A1(OutData[67]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A(OutData[11]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3), .B(FreshRand[34]), .ZN(SlicesFromChi[57]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[67]), .A2(OutData[23]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7), .ZN(SlicesFromChi[62]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U3 ( 
        .A1(OutData[54]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U2 ( 
        .A(OutData[23]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A(FreshRand[37]), .B(OutData[67]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[55]), .A2(OutData[54]), .ZN(SlicesFromChi[67]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5), .ZN(SlicesFromChi[72]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A1(OutData[55]), .A2(OutData[11]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A(FreshRand[43]), .B(OutData[54]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[77]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[36]), .A2(OutData[17]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[30]), .B(OutData[30]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[82]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[48]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[17]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[33]), .B(OutData[36]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[36]), .ZN(SlicesFromChi[87]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[48]), .A2(OutData[4]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[92]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[30]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[4]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[39]), .B(OutData[48]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[36]), .A2(OutData[30]), .ZN(SlicesFromChi[97]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[42]), .A2(OutData[36]), .ZN(SlicesFromChi[102]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[48]), .A2(OutData[42]), .ZN(SlicesFromChi[107]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[29]), .A2(OutData[48]), .ZN(SlicesFromChi[112]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[41]), .ZN(SlicesFromChi[117]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[29]), .A2(OutData[55]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3), .B(FreshRand[44]), .ZN(SlicesFromChi[122]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A1(OutData[55]), .A2(OutData[36]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3), .B(FreshRand[32]), .ZN(SlicesFromChi[127]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A1(OutData[36]), .A2(OutData[67]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3), .B(FreshRand[35]), .ZN(SlicesFromChi[132]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[67]), .A2(OutData[48]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3), .B(FreshRand[38]), .ZN(SlicesFromChi[137]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A1(OutData[48]), .A2(OutData[54]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3), .B(FreshRand[40]), .ZN(SlicesFromChi[142]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[54]), .A2(OutData[5]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U3 ( 
        .A(FreshRand[42]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5), .ZN(SlicesFromChi[147]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A1(OutData[36]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A(OutData[5]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[152]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[61]), .A2(OutData[17]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[31]), .B(OutData[55]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[157]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[73]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[17]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[34]), .B(OutData[61]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[37]), .ZN(SlicesFromChi[162]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[73]), .A2(OutData[4]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[167]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[55]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[4]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[40]), .B(OutData[73]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[61]), .A2(OutData[55]), .ZN(SlicesFromChi[172]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3), .B(FreshRand[32]), .ZN(SlicesFromChi[177]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[61]), .A2(OutData[42]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[35]), .ZN(SlicesFromChi[182]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[42]), .A2(OutData[73]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3), .B(FreshRand[38]), .ZN(SlicesFromChi[187]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[73]), .A2(OutData[29]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[39]), .ZN(SlicesFromChi[192]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[29]), .A2(OutData[5]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(FreshRand[43]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[197]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[61]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(OutData[5]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A1(OutData[67]), .A2(OutData[61]), .ZN(SlicesFromChi[202]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[73]), .A2(OutData[67]), .ZN(SlicesFromChi[207]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A1(OutData[54]), .A2(OutData[73]), .ZN(SlicesFromChi[212]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3), .B(FreshRand[41]), .ZN(SlicesFromChi[217]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[54]), .A2(OutData[30]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3), .B(FreshRand[44]), .ZN(SlicesFromChi[222]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A1(OutData[30]), .A2(OutData[61]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(OutData[20]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7), .ZN(SlicesFromChi[3]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[7]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(OutData[1]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A(OutData[1]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[8]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A1(OutData[13]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(OutData[7]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U3 ( 
        .A(OutData[7]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7), .ZN(SlicesFromChi[13]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A1(OutData[19]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A(OutData[13]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A(OutData[13]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[18]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A1(OutData[20]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(OutData[19]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U3 ( 
        .A(OutData[19]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7), .ZN(SlicesFromChi[23]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U2 ( 
        .A1(OutData[1]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A(OutData[20]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U3 ( 
        .A(FreshRand[45]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5), .ZN(SlicesFromChi[28]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A1(OutData[32]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A(OutData[1]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[48]), .ZN(SlicesFromChi[33]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[32]), .A2(OutData[13]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7), .ZN(SlicesFromChi[38]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U3 ( 
        .A1(OutData[44]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(OutData[13]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A(FreshRand[51]), .B(OutData[32]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[45]), .A2(OutData[44]), .ZN(SlicesFromChi[43]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[48]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[45]), .A2(OutData[1]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(FreshRand[57]), .B(OutData[44]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U3 ( 
        .A(FreshRand[46]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5), .ZN(SlicesFromChi[53]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U2 ( 
        .A1(OutData[57]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A(OutData[1]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3), .B(FreshRand[49]), .ZN(SlicesFromChi[58]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[57]), .A2(OutData[13]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7), .ZN(SlicesFromChi[63]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U3 ( 
        .A1(OutData[69]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U2 ( 
        .A(OutData[13]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A(FreshRand[52]), .B(OutData[57]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[70]), .A2(OutData[69]), .ZN(SlicesFromChi[68]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5), .ZN(SlicesFromChi[73]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A1(OutData[70]), .A2(OutData[1]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A(FreshRand[58]), .B(OutData[69]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[78]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[26]), .A2(OutData[7]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[45]), .B(OutData[45]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[83]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[38]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[7]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[48]), .B(OutData[26]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[51]), .ZN(SlicesFromChi[88]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[38]), .A2(OutData[19]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[93]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[45]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[19]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[54]), .B(OutData[38]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[26]), .A2(OutData[45]), .ZN(SlicesFromChi[98]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[32]), .A2(OutData[26]), .ZN(SlicesFromChi[103]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[38]), .A2(OutData[32]), .ZN(SlicesFromChi[108]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[44]), .A2(OutData[38]), .ZN(SlicesFromChi[113]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[56]), .ZN(SlicesFromChi[118]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[44]), .A2(OutData[70]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3), .B(FreshRand[59]), .ZN(SlicesFromChi[123]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A1(OutData[70]), .A2(OutData[26]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3), .B(FreshRand[47]), .ZN(SlicesFromChi[128]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A1(OutData[26]), .A2(OutData[57]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3), .B(FreshRand[50]), .ZN(SlicesFromChi[133]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[57]), .A2(OutData[38]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3), .B(FreshRand[53]), .ZN(SlicesFromChi[138]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A1(OutData[38]), .A2(OutData[69]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3), .B(FreshRand[55]), .ZN(SlicesFromChi[143]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[69]), .A2(OutData[20]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U3 ( 
        .A(FreshRand[57]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5), .ZN(SlicesFromChi[148]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A1(OutData[26]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A(OutData[20]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[153]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[51]), .A2(OutData[7]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[46]), .B(OutData[70]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[158]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[63]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[7]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[49]), .B(OutData[51]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[52]), .ZN(SlicesFromChi[163]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[63]), .A2(OutData[19]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[168]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[70]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[19]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[55]), .B(OutData[63]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[51]), .A2(OutData[70]), .ZN(SlicesFromChi[173]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3), .B(FreshRand[47]), .ZN(SlicesFromChi[178]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[51]), .A2(OutData[32]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[50]), .ZN(SlicesFromChi[183]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[32]), .A2(OutData[63]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3), .B(FreshRand[53]), .ZN(SlicesFromChi[188]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[63]), .A2(OutData[44]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[54]), .ZN(SlicesFromChi[193]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[44]), .A2(OutData[20]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(FreshRand[58]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[198]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[51]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(OutData[20]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A1(OutData[57]), .A2(OutData[51]), .ZN(SlicesFromChi[203]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[63]), .A2(OutData[57]), .ZN(SlicesFromChi[208]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A1(OutData[69]), .A2(OutData[63]), .ZN(SlicesFromChi[213]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3), .B(FreshRand[56]), .ZN(SlicesFromChi[218]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[69]), .A2(OutData[45]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3), .B(FreshRand[59]), .ZN(SlicesFromChi[223]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A1(OutData[45]), .A2(OutData[51]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(OutData[10]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7), .ZN(SlicesFromChi[4]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[22]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(OutData[16]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A(OutData[16]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[9]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A1(OutData[3]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(OutData[22]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U3 ( 
        .A(OutData[22]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7), .ZN(SlicesFromChi[14]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A1(OutData[9]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A(OutData[3]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_c_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A(OutData[3]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[19]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A1(OutData[10]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(OutData[9]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U3 ( 
        .A(OutData[9]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7), .ZN(SlicesFromChi[24]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U2 ( 
        .A1(OutData[16]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A(OutData[10]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_0__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U3 ( 
        .A(FreshRand[60]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5), .ZN(SlicesFromChi[29]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A1(OutData[47]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A(OutData[16]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[63]), .ZN(SlicesFromChi[34]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[47]), .A2(OutData[3]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7), .ZN(SlicesFromChi[39]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U3 ( 
        .A1(OutData[34]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(OutData[3]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A(FreshRand[66]), .B(OutData[47]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[35]), .A2(OutData[34]), .ZN(SlicesFromChi[44]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[49]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[35]), .A2(OutData[16]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(FreshRand[72]), .B(OutData[34]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_1__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U3 ( 
        .A(FreshRand[61]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5), .ZN(SlicesFromChi[54]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U2 ( 
        .A1(OutData[72]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A(OutData[16]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_a_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3), .B(FreshRand[64]), .ZN(SlicesFromChi[59]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[72]), .A2(OutData[3]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7), .ZN(SlicesFromChi[64]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U3 ( 
        .A1(OutData[59]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U2 ( 
        .A(OutData[3]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A(FreshRand[67]), .B(OutData[72]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_c_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[60]), .A2(OutData[59]), .ZN(SlicesFromChi[69]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5), .ZN(SlicesFromChi[74]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A1(OutData[60]), .A2(OutData[16]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A(FreshRand[73]), .B(OutData[59]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_0__ComponentFunctionGen1_2__and_xor_inst_e_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[79]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[41]), .A2(OutData[22]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[60]), .B(OutData[35]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[84]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[28]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[22]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[63]), .B(OutData[41]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[66]), .ZN(SlicesFromChi[89]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[28]), .A2(OutData[9]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[94]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[35]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[9]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[69]), .B(OutData[28]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[41]), .A2(OutData[35]), .ZN(SlicesFromChi[99]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[47]), .A2(OutData[41]), .ZN(SlicesFromChi[104]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[28]), .A2(OutData[47]), .ZN(SlicesFromChi[109]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[34]), .A2(OutData[28]), .ZN(SlicesFromChi[114]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[71]), .ZN(SlicesFromChi[119]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[34]), .A2(OutData[60]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3), .B(FreshRand[74]), .ZN(SlicesFromChi[124]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A1(OutData[60]), .A2(OutData[41]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_1__and_xor_inst_e_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3), .B(FreshRand[62]), .ZN(SlicesFromChi[129]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A1(OutData[41]), .A2(OutData[72]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_a_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3), .B(FreshRand[65]), .ZN(SlicesFromChi[134]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[72]), .A2(OutData[28]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3), .B(FreshRand[68]), .ZN(SlicesFromChi[139]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A1(OutData[28]), .A2(OutData[59]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3), .B(FreshRand[70]), .ZN(SlicesFromChi[144]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[59]), .A2(OutData[10]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U3 ( 
        .A(FreshRand[72]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5), .ZN(SlicesFromChi[149]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A1(OutData[41]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A(OutData[10]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_1__ComponentFunctionGen1_2__and_xor_inst_e_n4) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U3 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5), .ZN(SlicesFromChi[154]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U2 ( 
        .A1(OutData[66]), .A2(OutData[22]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n5) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_U1 ( 
        .A(FreshRand[61]), .B(OutData[60]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_a_n6) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7), .ZN(SlicesFromChi[159]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U3 ( 
        .A1(OutData[53]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U2 ( 
        .A(OutData[22]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_U1 ( 
        .A(FreshRand[64]), .B(OutData[66]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_b_n8) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3), .B(FreshRand[67]), .ZN(SlicesFromChi[164]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_U1 ( 
        .A1(OutData[53]), .A2(OutData[9]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U4 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7), .ZN(SlicesFromChi[169]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U3 ( 
        .A1(OutData[60]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n7) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U2 ( 
        .A(OutData[9]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n6) );
  XOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_U1 ( 
        .A(FreshRand[70]), .B(OutData[53]), .Z(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_d_n8) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_0__and_xor_inst_e_U1 ( 
        .A1(OutData[66]), .A2(OutData[60]), .ZN(SlicesFromChi[174]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3), .B(FreshRand[62]), .ZN(SlicesFromChi[179]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_U1 ( 
        .A1(OutData[66]), .A2(OutData[47]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_a_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3), .B(FreshRand[65]), .ZN(SlicesFromChi[184]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_U1 ( 
        .A1(OutData[47]), .A2(OutData[53]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_b_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3), .B(FreshRand[68]), .ZN(SlicesFromChi[189]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_U1 ( 
        .A1(OutData[53]), .A2(OutData[34]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_c_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3), .B(FreshRand[69]), .ZN(SlicesFromChi[194]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_U1 ( 
        .A1(OutData[34]), .A2(OutData[10]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U3 ( 
        .A(FreshRand[73]), .B(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5), .ZN(SlicesFromChi[199]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U2 ( 
        .A1(OutData[66]), .A2(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n5) );
  INV_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_U1 ( 
        .A(OutData[10]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_1__and_xor_inst_e_n4) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_a_U1 ( 
        .A1(OutData[72]), .A2(OutData[66]), .ZN(SlicesFromChi[204]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_b_U1 ( 
        .A1(OutData[53]), .A2(OutData[72]), .ZN(SlicesFromChi[209]) );
  AND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_c_U1 ( 
        .A1(OutData[59]), .A2(OutData[53]), .ZN(SlicesFromChi[214]) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3), .B(FreshRand[71]), .ZN(SlicesFromChi[219]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_U1 ( 
        .A1(OutData[59]), .A2(OutData[35]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_d_n3) );
  XNOR2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_U2 ( 
        .A(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3), .B(FreshRand[74]), .ZN(SlicesFromChi[224]) );
  NAND2_X1 CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_U1 ( 
        .A1(OutData[35]), .A2(OutData[66]), .ZN(
        CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_ComponentFunctionGen1_2__ComponentFunctionGen1_2__and_xor_inst_e_n3) );
  OAI221_X1 KECCAK_CONTROL_U33 ( .B1(KECCAK_CONTROL_n6), .B2(
        KECCAK_CONTROL_n62), .C1(KECCAK_CONTROL_n6), .C2(KECCAK_CONTROL_n61), 
        .A(KECCAK_CONTROL_n60), .ZN(KECCAK_CONTROL_n34) );
  NAND3_X1 KECCAK_CONTROL_U32 ( .A1(KECCAK_CONTROL_n59), .A2(
        KECCAK_CONTROL_n58), .A3(KECCAK_CONTROL_n6), .ZN(KECCAK_CONTROL_n60)
         );
  OAI22_X1 KECCAK_CONTROL_U31 ( .A1(KECCAK_CONTROL_n27), .A2(
        KECCAK_CONTROL_n62), .B1(KECCAK_CONTROL_n57), .B2(KECCAK_CONTROL_n61), 
        .ZN(KECCAK_CONTROL_n35) );
  NAND2_X1 KECCAK_CONTROL_U30 ( .A1(KECCAK_CONTROL_n59), .A2(
        KECCAK_CONTROL_n27), .ZN(KECCAK_CONTROL_n61) );
  OR2_X1 KECCAK_CONTROL_U29 ( .A1(KECCAK_CONTROL_n40), .A2(KECCAK_CONTROL_n31), 
        .ZN(KECCAK_CONTROL_n57) );
  AOI21_X1 KECCAK_CONTROL_U28 ( .B1(KECCAK_CONTROL_n59), .B2(
        KECCAK_CONTROL_n31), .A(KECCAK_CONTROL_n56), .ZN(KECCAK_CONTROL_n62)
         );
  OAI22_X1 KECCAK_CONTROL_U27 ( .A1(KECCAK_CONTROL_n31), .A2(
        KECCAK_CONTROL_n55), .B1(KECCAK_CONTROL_n54), .B2(KECCAK_CONTROL_n40), 
        .ZN(KECCAK_CONTROL_n36) );
  NAND2_X1 KECCAK_CONTROL_U26 ( .A1(KECCAK_CONTROL_n59), .A2(
        KECCAK_CONTROL_n31), .ZN(KECCAK_CONTROL_n54) );
  INV_X1 KECCAK_CONTROL_U25 ( .A(KECCAK_CONTROL_n53), .ZN(KECCAK_CONTROL_n59)
         );
  INV_X1 KECCAK_CONTROL_U24 ( .A(KECCAK_CONTROL_n56), .ZN(KECCAK_CONTROL_n55)
         );
  OAI21_X1 KECCAK_CONTROL_U23 ( .B1(Reset), .B2(
        KECCAK_CONTROL_RoundCountxDP_0_), .A(KECCAK_CONTROL_n52), .ZN(
        KECCAK_CONTROL_n56) );
  AOI22_X1 KECCAK_CONTROL_U22 ( .A1(KECCAK_CONTROL_RoundCountxDP_0_), .A2(
        KECCAK_CONTROL_n52), .B1(KECCAK_CONTROL_n53), .B2(KECCAK_CONTROL_n40), 
        .ZN(KECCAK_CONTROL_n37) );
  OAI22_X1 KECCAK_CONTROL_U21 ( .A1(KECCAK_CONTROL_n32), .A2(
        KECCAK_CONTROL_n52), .B1(KECCAK_CONTROL_n51), .B2(KECCAK_CONTROL_n53), 
        .ZN(KECCAK_CONTROL_n38) );
  NAND2_X1 KECCAK_CONTROL_U20 ( .A1(KECCAK_CONTROL_n42), .A2(
        KECCAK_CONTROL_n52), .ZN(KECCAK_CONTROL_n53) );
  NAND3_X1 KECCAK_CONTROL_U19 ( .A1(KECCAK_CONTROL_n42), .A2(
        KECCAK_CONTROL_n50), .A3(KECCAK_CONTROL_n49), .ZN(KECCAK_CONTROL_n52)
         );
  AOI21_X1 KECCAK_CONTROL_U18 ( .B1(KECCAK_CONTROL_n39), .B2(
        KECCAK_CONTROL_n50), .A(Reset), .ZN(KECCAK_CONTROL_n48) );
  AOI21_X1 KECCAK_CONTROL_U17 ( .B1(KECCAK_CONTROL_n14), .B2(
        KECCAK_CONTROL_n47), .A(Reset), .ZN(KECCAK_CONTROL_n29) );
  INV_X1 KECCAK_CONTROL_U16 ( .A(KECCAK_CONTROL_n46), .ZN(KECCAK_CONTROL_n47)
         );
  AOI221_X1 KECCAK_CONTROL_U15 ( .B1(KECCAK_CONTROL_n26), .B2(
        KECCAK_CONTROL_n50), .C1(KECCAK_CONTROL_n46), .C2(KECCAK_CONTROL_n50), 
        .A(Reset), .ZN(KECCAK_CONTROL_n28) );
  NOR2_X1 KECCAK_CONTROL_U14 ( .A1(KECCAK_CONTROL_n5), .A2(KECCAK_CONTROL_n49), 
        .ZN(KECCAK_CONTROL_n46) );
  NAND3_X1 KECCAK_CONTROL_U13 ( .A1(KECCAK_CONTROL_n41), .A2(
        KECCAK_CONTROL_n15), .A3(KECCAK_CONTROL_n14), .ZN(KECCAK_CONTROL_n49)
         );
  NAND3_X1 KECCAK_CONTROL_U12 ( .A1(KECCAK_CONTROL_n39), .A2(
        KECCAK_CONTROL_n14), .A3(KECCAK_CONTROL_n26), .ZN(KECCAK_CONTROL_n50)
         );
  NOR3_X1 KECCAK_CONTROL_U11 ( .A1(KECCAK_CONTROL_n14), .A2(KECCAK_CONTROL_n39), .A3(KECCAK_CONTROL_n41), .ZN(Ready) );
  AOI21_X1 KECCAK_CONTROL_U10 ( .B1(KECCAK_CONTROL_n51), .B2(
        KECCAK_CONTROL_n45), .A(Reset), .ZN(KECCAK_CONTROL_N32) );
  INV_X1 KECCAK_CONTROL_U9 ( .A(KECCAK_CONTROL_n44), .ZN(KECCAK_CONTROL_n45)
         );
  AOI211_X1 KECCAK_CONTROL_U8 ( .C1(KECCAK_CONTROL_n27), .C2(
        KECCAK_CONTROL_n31), .A(KECCAK_CONTROL_n58), .B(KECCAK_CONTROL_n6), 
        .ZN(KECCAK_CONTROL_n44) );
  XNOR2_X1 KECCAK_CONTROL_U7 ( .A(KECCAK_CONTROL_n43), .B(KECCAK_CONTROL_n32), 
        .ZN(KECCAK_CONTROL_n51) );
  NAND2_X1 KECCAK_CONTROL_U6 ( .A1(KECCAK_CONTROL_RoundCountxDP_3_), .A2(
        KECCAK_CONTROL_n58), .ZN(KECCAK_CONTROL_n43) );
  NOR3_X1 KECCAK_CONTROL_U5 ( .A1(KECCAK_CONTROL_n31), .A2(KECCAK_CONTROL_n27), 
        .A3(KECCAK_CONTROL_n40), .ZN(KECCAK_CONTROL_n58) );
  NOR2_X1 KECCAK_CONTROL_U4 ( .A1(Reset), .A2(KECCAK_CONTROL_n5), .ZN(
        Lastround) );
  INV_X1 KECCAK_CONTROL_U3 ( .A(Reset), .ZN(KECCAK_CONTROL_n42) );
  DFF_X1 KECCAK_CONTROL_CtrlStatexDP_reg_0_ ( .D(KECCAK_CONTROL_n48), .CK(
        Clock), .Q(KECCAK_CONTROL_n15), .QN(KECCAK_CONTROL_n39) );
  DFF_X1 KECCAK_CONTROL_RoundCountxDP_reg_0_ ( .D(KECCAK_CONTROL_n37), .CK(
        Clock), .Q(KECCAK_CONTROL_RoundCountxDP_0_), .QN(KECCAK_CONTROL_n40)
         );
  DFF_X1 KECCAK_CONTROL_RoundCountxDP_reg_1_ ( .D(KECCAK_CONTROL_n36), .CK(
        Clock), .Q(KECCAK_CONTROL_RoundCountxDP_1_), .QN(KECCAK_CONTROL_n31)
         );
  DFF_X1 KECCAK_CONTROL_RoundCountxDP_reg_2_ ( .D(KECCAK_CONTROL_n35), .CK(
        Clock), .Q(KECCAK_CONTROL_RoundCountxDP_2_), .QN(KECCAK_CONTROL_n27)
         );
  DFF_X1 KECCAK_CONTROL_RoundCountxDP_reg_3_ ( .D(KECCAK_CONTROL_n34), .CK(
        Clock), .Q(KECCAK_CONTROL_RoundCountxDP_3_), .QN(KECCAK_CONTROL_n6) );
  DFF_X1 KECCAK_CONTROL_RoundCountxDP_reg_4_ ( .D(KECCAK_CONTROL_n38), .CK(
        Clock), .Q(KECCAK_CONTROL_RoundCountxDP_4_), .QN(KECCAK_CONTROL_n32)
         );
  DFF_X1 KECCAK_CONTROL_CtrlStatexDP_reg_1_ ( .D(KECCAK_CONTROL_n28), .CK(
        Clock), .Q(KECCAK_CONTROL_n41), .QN(KECCAK_CONTROL_n26) );
  DFF_X1 KECCAK_CONTROL_CtrlStatexDP_reg_2_ ( .D(KECCAK_CONTROL_n29), .CK(
        Clock), .Q(), .QN(KECCAK_CONTROL_n14) );
  DFF_X1 KECCAK_CONTROL_RoundCountLastxDP_reg ( .D(KECCAK_CONTROL_N32), .CK(
        Clock), .Q(), .QN(KECCAK_CONTROL_n5) );
  AOI221_X1 KECCAK_CONTROL_RC_GEN_U4 ( .B1(KECCAK_CONTROL_RoundCountxDP_0_), 
        .B2(KECCAK_CONTROL_RC_GEN_n3), .C1(KECCAK_CONTROL_RC_GEN_n2), .C2(
        KECCAK_CONTROL_RC_GEN_n3), .A(KECCAK_CONTROL_RoundCountxDP_4_), .ZN(
        IotaRC_0_) );
  XOR2_X1 KECCAK_CONTROL_RC_GEN_U3 ( .A(KECCAK_CONTROL_RoundCountxDP_1_), .B(
        KECCAK_CONTROL_RoundCountxDP_3_), .Z(KECCAK_CONTROL_RC_GEN_n2) );
  INV_X1 KECCAK_CONTROL_RC_GEN_U2 ( .A(KECCAK_CONTROL_RoundCountxDP_2_), .ZN(
        KECCAK_CONTROL_RC_GEN_n3) );
endmodule

