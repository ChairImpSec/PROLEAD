module circuit ( ClkxCI, RstxBI, PTxDI, KxDI, randomS2, randomS3, randomS4, 
        randomS5, StartxSI, DonexSO, CxDO );
  input [15:0] PTxDI;
  input [15:0] KxDI;
  input [15:0] randomS2;
  input [7:0] randomS3;
  input [15:0] randomS4;
  input [31:0] randomS5;
  output [15:0] CxDO;
  input ClkxCI, RstxBI, StartxSI;
  output DonexSO;
  wire   disableKeyRegsxS, ClkKeyRegxC, StateKEYSCHEDULExS, nextRCONxS,
         showRCONxS, FinishedxS, StateKEYADDITION1o3xS, LastRoundxS,
         doMixColumnsxS, n114, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341,
         aes_ctrl_lsfr_23_cycles_1_n24, aes_ctrl_lsfr_23_cycles_1_n23,
         aes_ctrl_lsfr_23_cycles_1_n22, aes_ctrl_lsfr_23_cycles_1_n21,
         aes_ctrl_lsfr_23_cycles_1_n20, aes_ctrl_lsfr_23_cycles_1_n19,
         aes_ctrl_lsfr_23_cycles_1_n18, aes_ctrl_lsfr_23_cycles_1_n17,
         aes_ctrl_lsfr_23_cycles_1_n16, aes_ctrl_lsfr_23_cycles_1_n15,
         aes_ctrl_lsfr_23_cycles_1_n14, aes_ctrl_lsfr_23_cycles_1_n13,
         aes_ctrl_lsfr_23_cycles_1_n11, aes_ctrl_lsfr_23_cycles_1_n10,
         aes_ctrl_lsfr_23_cycles_1_n8, aes_ctrl_lsfr_23_cycles_1_n7,
         aes_ctrl_lsfr_23_cycles_1_n5, aes_ctrl_lsfr_23_cycles_1_n3,
         aes_ctrl_lsfr_23_cycles_1_n1, aes_ctrl_lsfr_23_cycles_1_n39,
         aes_ctrl_lsfr_23_cycles_1_n38, aes_ctrl_lsfr_23_cycles_1_n37,
         aes_ctrl_lsfr_23_cycles_1_n36, aes_ctrl_lsfr_23_cycles_1_n35,
         aes_ctrl_lsfr_23_cycles_1_n12, aes_ctrl_lsfr_23_cycles_1_n9,
         aes_ctrl_lsfr_23_cycles_1_n6, aes_ctrl_lsfr_23_cycles_1_n4,
         aes_ctrl_lsfr_23_cycles_1_n2, aes_ctrl_lsfr_23_cycles_1_N83,
         aes_ctrl_lsfr_23_cycles_1_N66, aes_ctrl_lsfr_23_cycles_1_N16,
         rcon_1_n45, rcon_1_n44, rcon_1_n43, rcon_1_n42, rcon_1_n41,
         rcon_1_n40, rcon_1_n39, rcon_1_n38, rcon_1_n37, rcon_1_n36,
         rcon_1_n34, rcon_1_n33, rcon_1_n32, rcon_1_n31, rcon_1_n30,
         rcon_1_n29, rcon_1_n28, rcon_1_n16, rcon_1_n15, rcon_1_n14,
         rcon_1_n13, rcon_1_n12, rcon_1_n11, rcon_1_n35, rcon_1_n26,
         rcon_1_n25, rcon_1_n24, rcon_1_n23, rcon_1_n22, rcon_1_n21,
         rcon_1_n20, rcon_1_n19, rcon_1_n18, rcon_1_n17, rcon_1_n9, rcon_1_n4,
         SBOX_s1_linMapOut_0__0_, SBOX_s1_linMapOut_0__1_,
         SBOX_s1_linMapOut_0__3_, SBOX_s1_linMapOut_0__4_,
         SBOX_s1_linMapOut_0__5_, SBOX_s1_linMapOut_0__6_,
         SBOX_s1_linMapOut_0__7_, SBOX_s1_linMapOut_1__0_,
         SBOX_s1_linMapOut_1__1_, SBOX_s1_linMapOut_1__3_,
         SBOX_s1_linMapOut_1__4_, SBOX_s1_linMapOut_1__5_,
         SBOX_s1_linMapOut_1__6_, SBOX_s1_linMapOut_1__7_,
         SBOX_s1_input_mapping_1_n23, SBOX_s1_input_mapping_1_n22,
         SBOX_s1_input_mapping_1_n21, SBOX_s1_input_mapping_1_n20,
         SBOX_s1_input_mapping_1_n19, SBOX_s1_input_mapping_1_n18,
         SBOX_s1_input_mapping_1_n17, SBOX_s1_input_mapping_0_n23,
         SBOX_s1_input_mapping_0_n22, SBOX_s1_input_mapping_0_n21,
         SBOX_s1_input_mapping_0_n20, SBOX_s1_input_mapping_0_n19,
         SBOX_s1_input_mapping_0_n18, SBOX_s1_input_mapping_0_n17, SBOX_s2_n16,
         SBOX_s2_n15, SBOX_s2_n14, SBOX_s2_n13, SBOX_s2_n12, SBOX_s2_n11,
         SBOX_s2_n10, SBOX_s2_n9, SBOX_s2_n8, SBOX_s2_n7, SBOX_s2_n6,
         SBOX_s2_n5, SBOX_s2_n4, SBOX_s2_n3, SBOX_s2_n2, SBOX_s2_n1,
         SBOX_s2_regOut_0__1__0_, SBOX_s2_regOut_0__1__1_,
         SBOX_s2_regOut_0__1__2_, SBOX_s2_regOut_0__1__3_,
         SBOX_s2_regOut_0__2__0_, SBOX_s2_regOut_0__2__1_,
         SBOX_s2_regOut_0__2__2_, SBOX_s2_regOut_0__2__3_,
         SBOX_s2_regOut_1__1__0_, SBOX_s2_regOut_1__1__1_,
         SBOX_s2_regOut_1__1__2_, SBOX_s2_regOut_1__1__3_,
         SBOX_s2_regOut_1__2__0_, SBOX_s2_regOut_1__2__1_,
         SBOX_s2_regOut_1__2__2_, SBOX_s2_regOut_1__2__3_,
         SBOX_s2_gf2_mul_out_0__0__0_, SBOX_s2_gf2_mul_out_0__0__1_,
         SBOX_s2_gf2_mul_out_0__0__2_, SBOX_s2_gf2_mul_out_0__0__3_,
         SBOX_s2_gf2_mul_out_1__1__0_, SBOX_s2_gf2_mul_out_1__1__1_,
         SBOX_s2_gf2_mul_out_1__1__2_, SBOX_s2_gf2_mul_out_1__1__3_,
         SBOX_s2_mul1_1_1_n77, SBOX_s2_mul1_1_1_n76, SBOX_s2_mul1_1_1_n75,
         SBOX_s2_mul1_1_1_n74, SBOX_s2_mul1_1_1_n73, SBOX_s2_mul1_1_1_n72,
         SBOX_s2_mul1_1_1_n71, SBOX_s2_mul1_1_1_n70, SBOX_s2_mul1_1_1_n69,
         SBOX_s2_mul1_1_1_n68, SBOX_s2_mul1_1_1_n67, SBOX_s2_mul1_1_1_n66,
         SBOX_s2_mul1_1_1_n65, SBOX_s2_mul1_1_1_n64, SBOX_s2_mul1_1_1_n63,
         SBOX_s2_mul1_1_1_n62, SBOX_s2_mul1_1_1_n61, SBOX_s2_mul1_1_1_n59,
         SBOX_s2_mul1_1_1_n58, SBOX_s2_mul1_1_1_n57, SBOX_s2_mul1_1_1_n56,
         SBOX_s2_mul1_1_1_n55, SBOX_s2_mul1_1_1_n54, SBOX_s2_mul1_1_1_n53,
         SBOX_s2_mul1_1_0_n77, SBOX_s2_mul1_1_0_n76, SBOX_s2_mul1_1_0_n75,
         SBOX_s2_mul1_1_0_n74, SBOX_s2_mul1_1_0_n73, SBOX_s2_mul1_1_0_n72,
         SBOX_s2_mul1_1_0_n71, SBOX_s2_mul1_1_0_n70, SBOX_s2_mul1_1_0_n69,
         SBOX_s2_mul1_1_0_n68, SBOX_s2_mul1_1_0_n67, SBOX_s2_mul1_1_0_n66,
         SBOX_s2_mul1_1_0_n65, SBOX_s2_mul1_1_0_n64, SBOX_s2_mul1_1_0_n63,
         SBOX_s2_mul1_1_0_n62, SBOX_s2_mul1_1_0_n61, SBOX_s2_mul1_1_0_n60,
         SBOX_s2_mul1_1_0_n59, SBOX_s2_mul1_1_0_n58, SBOX_s2_mul1_1_0_n57,
         SBOX_s2_mul1_1_0_n56, SBOX_s2_mul1_1_0_n54, SBOX_s2_mul1_1_0_n53,
         SBOX_s2_mul1_0_1_n77, SBOX_s2_mul1_0_1_n76, SBOX_s2_mul1_0_1_n75,
         SBOX_s2_mul1_0_1_n74, SBOX_s2_mul1_0_1_n73, SBOX_s2_mul1_0_1_n72,
         SBOX_s2_mul1_0_1_n71, SBOX_s2_mul1_0_1_n70, SBOX_s2_mul1_0_1_n69,
         SBOX_s2_mul1_0_1_n68, SBOX_s2_mul1_0_1_n67, SBOX_s2_mul1_0_1_n66,
         SBOX_s2_mul1_0_1_n65, SBOX_s2_mul1_0_1_n64, SBOX_s2_mul1_0_1_n63,
         SBOX_s2_mul1_0_1_n62, SBOX_s2_mul1_0_1_n61, SBOX_s2_mul1_0_1_n60,
         SBOX_s2_mul1_0_1_n59, SBOX_s2_mul1_0_1_n58, SBOX_s2_mul1_0_1_n57,
         SBOX_s2_mul1_0_1_n56, SBOX_s2_mul1_0_1_n54, SBOX_s2_mul1_0_1_n53,
         SBOX_s2_mul1_0_0_n77, SBOX_s2_mul1_0_0_n76, SBOX_s2_mul1_0_0_n75,
         SBOX_s2_mul1_0_0_n74, SBOX_s2_mul1_0_0_n73, SBOX_s2_mul1_0_0_n72,
         SBOX_s2_mul1_0_0_n71, SBOX_s2_mul1_0_0_n70, SBOX_s2_mul1_0_0_n69,
         SBOX_s2_mul1_0_0_n68, SBOX_s2_mul1_0_0_n67, SBOX_s2_mul1_0_0_n66,
         SBOX_s2_mul1_0_0_n65, SBOX_s2_mul1_0_0_n64, SBOX_s2_mul1_0_0_n63,
         SBOX_s2_mul1_0_0_n62, SBOX_s2_mul1_0_0_n61, SBOX_s2_mul1_0_0_n60,
         SBOX_s2_mul1_0_0_n59, SBOX_s2_mul1_0_0_n58, SBOX_s2_mul1_0_0_n57,
         SBOX_s2_mul1_0_0_n55, SBOX_s2_mul1_0_0_n54, SBOX_s2_mul1_0_0_n53,
         SBOX_s3_n8, SBOX_s3_n7, SBOX_s3_n6, SBOX_s3_n5, SBOX_s3_n4,
         SBOX_s3_n3, SBOX_s3_n2, SBOX_s3_n1, SBOX_s3_regOut_0__3__0_,
         SBOX_s3_regOut_0__3__1_, SBOX_s3_regOut_0__4__0_,
         SBOX_s3_regOut_0__4__1_, SBOX_s3_regOut_1__3__0_,
         SBOX_s3_regOut_1__3__1_, SBOX_s3_regOut_1__4__0_,
         SBOX_s3_regOut_1__4__1_, SBOX_s3_gf2_mul_out_0__0__0_,
         SBOX_s3_gf2_mul_out_0__0__1_, SBOX_s3_gf2_mul_out_1__1__0_,
         SBOX_s3_gf2_mul_out_1__1__1_, SBOX_s3_mul1_1_1_n14,
         SBOX_s3_mul1_1_1_n13, SBOX_s3_mul1_1_1_n12, SBOX_s3_mul1_1_1_n11,
         SBOX_s3_mul1_1_0_n14, SBOX_s3_mul1_1_0_n13, SBOX_s3_mul1_1_0_n12,
         SBOX_s3_mul1_1_0_n11, SBOX_s3_mul1_0_1_n14, SBOX_s3_mul1_0_1_n13,
         SBOX_s3_mul1_0_1_n12, SBOX_s3_mul1_0_1_n11, SBOX_s3_mul1_0_0_n14,
         SBOX_s3_mul1_0_0_n13, SBOX_s3_mul1_0_0_n12, SBOX_s3_mul1_0_0_n11,
         SBOX_s4_n8, SBOX_s4_n7, SBOX_s4_n6, SBOX_s4_n5, SBOX_s4_n4,
         SBOX_s4_n3, SBOX_s4_n2, SBOX_s4_n1, SBOX_s4_regOut_0__1__0_,
         SBOX_s4_regOut_0__1__1_, SBOX_s4_regOut_0__1__2_,
         SBOX_s4_regOut_0__1__3_, SBOX_s4_regOut_0__2__0_,
         SBOX_s4_regOut_0__2__1_, SBOX_s4_regOut_0__2__2_,
         SBOX_s4_regOut_0__2__3_, SBOX_s4_regOut_1__1__0_,
         SBOX_s4_regOut_1__1__1_, SBOX_s4_regOut_1__1__2_,
         SBOX_s4_regOut_1__1__3_, SBOX_s4_regOut_1__2__0_,
         SBOX_s4_regOut_1__2__1_, SBOX_s4_regOut_1__2__2_,
         SBOX_s4_regOut_1__2__3_, SBOX_s4_inv_out_0__0_, SBOX_s4_inv_out_0__1_,
         SBOX_s4_inv_out_1__0_, SBOX_s4_inv_out_1__1_, SBOX_s4_mul1_1_1_n14,
         SBOX_s4_mul1_1_1_n13, SBOX_s4_mul1_1_1_n12, SBOX_s4_mul1_1_1_n11,
         SBOX_s4_mul1_1_0_n14, SBOX_s4_mul1_1_0_n13, SBOX_s4_mul1_1_0_n12,
         SBOX_s4_mul1_1_0_n11, SBOX_s4_mul1_0_1_n14, SBOX_s4_mul1_0_1_n13,
         SBOX_s4_mul1_0_1_n12, SBOX_s4_mul1_0_1_n11, SBOX_s4_mul1_0_0_n14,
         SBOX_s4_mul1_0_0_n13, SBOX_s4_mul1_0_0_n12, SBOX_s4_mul1_0_0_n11,
         SBOX_s4_mul2_1_1_n14, SBOX_s4_mul2_1_1_n13, SBOX_s4_mul2_1_1_n12,
         SBOX_s4_mul2_1_1_n11, SBOX_s4_mul2_1_0_n14, SBOX_s4_mul2_1_0_n13,
         SBOX_s4_mul2_1_0_n12, SBOX_s4_mul2_1_0_n11, SBOX_s4_mul2_0_1_n14,
         SBOX_s4_mul2_0_1_n13, SBOX_s4_mul2_0_1_n12, SBOX_s4_mul2_0_1_n11,
         SBOX_s4_mul2_0_0_n14, SBOX_s4_mul2_0_0_n13, SBOX_s4_mul2_0_0_n12,
         SBOX_s4_mul2_0_0_n11, SBOX_s5_n16, SBOX_s5_n15, SBOX_s5_n14,
         SBOX_s5_n13, SBOX_s5_n12, SBOX_s5_n11, SBOX_s5_n10, SBOX_s5_n9,
         SBOX_s5_n8, SBOX_s5_n7, SBOX_s5_n6, SBOX_s5_n5, SBOX_s5_n4,
         SBOX_s5_n3, SBOX_s5_n2, SBOX_s5_n1, SBOX_s5_mul1_1_1_n76,
         SBOX_s5_mul1_1_1_n75, SBOX_s5_mul1_1_1_n74, SBOX_s5_mul1_1_1_n73,
         SBOX_s5_mul1_1_1_n72, SBOX_s5_mul1_1_1_n71, SBOX_s5_mul1_1_1_n70,
         SBOX_s5_mul1_1_1_n69, SBOX_s5_mul1_1_1_n68, SBOX_s5_mul1_1_1_n67,
         SBOX_s5_mul1_1_1_n66, SBOX_s5_mul1_1_1_n65, SBOX_s5_mul1_1_1_n64,
         SBOX_s5_mul1_1_1_n63, SBOX_s5_mul1_1_1_n62, SBOX_s5_mul1_1_1_n61,
         SBOX_s5_mul1_1_1_n60, SBOX_s5_mul1_1_1_n59, SBOX_s5_mul1_1_1_n58,
         SBOX_s5_mul1_1_1_n57, SBOX_s5_mul1_1_1_n56, SBOX_s5_mul1_1_1_n55,
         SBOX_s5_mul1_1_1_n54, SBOX_s5_mul1_1_1_n53, SBOX_s5_mul1_1_0_n77,
         SBOX_s5_mul1_1_0_n76, SBOX_s5_mul1_1_0_n75, SBOX_s5_mul1_1_0_n74,
         SBOX_s5_mul1_1_0_n73, SBOX_s5_mul1_1_0_n72, SBOX_s5_mul1_1_0_n71,
         SBOX_s5_mul1_1_0_n70, SBOX_s5_mul1_1_0_n69, SBOX_s5_mul1_1_0_n68,
         SBOX_s5_mul1_1_0_n67, SBOX_s5_mul1_1_0_n66, SBOX_s5_mul1_1_0_n65,
         SBOX_s5_mul1_1_0_n64, SBOX_s5_mul1_1_0_n63, SBOX_s5_mul1_1_0_n62,
         SBOX_s5_mul1_1_0_n61, SBOX_s5_mul1_1_0_n60, SBOX_s5_mul1_1_0_n59,
         SBOX_s5_mul1_1_0_n58, SBOX_s5_mul1_1_0_n57, SBOX_s5_mul1_1_0_n56,
         SBOX_s5_mul1_1_0_n54, SBOX_s5_mul1_1_0_n53, SBOX_s5_mul1_0_1_n76,
         SBOX_s5_mul1_0_1_n75, SBOX_s5_mul1_0_1_n74, SBOX_s5_mul1_0_1_n73,
         SBOX_s5_mul1_0_1_n72, SBOX_s5_mul1_0_1_n71, SBOX_s5_mul1_0_1_n70,
         SBOX_s5_mul1_0_1_n69, SBOX_s5_mul1_0_1_n68, SBOX_s5_mul1_0_1_n67,
         SBOX_s5_mul1_0_1_n66, SBOX_s5_mul1_0_1_n65, SBOX_s5_mul1_0_1_n64,
         SBOX_s5_mul1_0_1_n63, SBOX_s5_mul1_0_1_n62, SBOX_s5_mul1_0_1_n61,
         SBOX_s5_mul1_0_1_n60, SBOX_s5_mul1_0_1_n59, SBOX_s5_mul1_0_1_n58,
         SBOX_s5_mul1_0_1_n57, SBOX_s5_mul1_0_1_n56, SBOX_s5_mul1_0_1_n55,
         SBOX_s5_mul1_0_1_n54, SBOX_s5_mul1_0_1_n53, SBOX_s5_mul1_0_0_n76,
         SBOX_s5_mul1_0_0_n75, SBOX_s5_mul1_0_0_n74, SBOX_s5_mul1_0_0_n73,
         SBOX_s5_mul1_0_0_n72, SBOX_s5_mul1_0_0_n71, SBOX_s5_mul1_0_0_n70,
         SBOX_s5_mul1_0_0_n69, SBOX_s5_mul1_0_0_n68, SBOX_s5_mul1_0_0_n67,
         SBOX_s5_mul1_0_0_n66, SBOX_s5_mul1_0_0_n65, SBOX_s5_mul1_0_0_n64,
         SBOX_s5_mul1_0_0_n63, SBOX_s5_mul1_0_0_n62, SBOX_s5_mul1_0_0_n61,
         SBOX_s5_mul1_0_0_n60, SBOX_s5_mul1_0_0_n59, SBOX_s5_mul1_0_0_n58,
         SBOX_s5_mul1_0_0_n57, SBOX_s5_mul1_0_0_n56, SBOX_s5_mul1_0_0_n55,
         SBOX_s5_mul1_0_0_n54, SBOX_s5_mul1_0_0_n53, SBOX_s5_mul2_1_1_n77,
         SBOX_s5_mul2_1_1_n76, SBOX_s5_mul2_1_1_n75, SBOX_s5_mul2_1_1_n74,
         SBOX_s5_mul2_1_1_n73, SBOX_s5_mul2_1_1_n72, SBOX_s5_mul2_1_1_n71,
         SBOX_s5_mul2_1_1_n70, SBOX_s5_mul2_1_1_n69, SBOX_s5_mul2_1_1_n68,
         SBOX_s5_mul2_1_1_n67, SBOX_s5_mul2_1_1_n66, SBOX_s5_mul2_1_1_n65,
         SBOX_s5_mul2_1_1_n64, SBOX_s5_mul2_1_1_n63, SBOX_s5_mul2_1_1_n62,
         SBOX_s5_mul2_1_1_n61, SBOX_s5_mul2_1_1_n60, SBOX_s5_mul2_1_1_n59,
         SBOX_s5_mul2_1_1_n58, SBOX_s5_mul2_1_1_n57, SBOX_s5_mul2_1_1_n56,
         SBOX_s5_mul2_1_1_n55, SBOX_s5_mul2_1_1_n54, SBOX_s5_mul2_1_0_n76,
         SBOX_s5_mul2_1_0_n75, SBOX_s5_mul2_1_0_n74, SBOX_s5_mul2_1_0_n73,
         SBOX_s5_mul2_1_0_n72, SBOX_s5_mul2_1_0_n71, SBOX_s5_mul2_1_0_n70,
         SBOX_s5_mul2_1_0_n69, SBOX_s5_mul2_1_0_n68, SBOX_s5_mul2_1_0_n67,
         SBOX_s5_mul2_1_0_n66, SBOX_s5_mul2_1_0_n65, SBOX_s5_mul2_1_0_n64,
         SBOX_s5_mul2_1_0_n63, SBOX_s5_mul2_1_0_n62, SBOX_s5_mul2_1_0_n61,
         SBOX_s5_mul2_1_0_n60, SBOX_s5_mul2_1_0_n59, SBOX_s5_mul2_1_0_n58,
         SBOX_s5_mul2_1_0_n57, SBOX_s5_mul2_1_0_n56, SBOX_s5_mul2_1_0_n55,
         SBOX_s5_mul2_1_0_n54, SBOX_s5_mul2_1_0_n53, SBOX_s5_mul2_0_1_n76,
         SBOX_s5_mul2_0_1_n75, SBOX_s5_mul2_0_1_n74, SBOX_s5_mul2_0_1_n73,
         SBOX_s5_mul2_0_1_n72, SBOX_s5_mul2_0_1_n71, SBOX_s5_mul2_0_1_n70,
         SBOX_s5_mul2_0_1_n69, SBOX_s5_mul2_0_1_n68, SBOX_s5_mul2_0_1_n67,
         SBOX_s5_mul2_0_1_n66, SBOX_s5_mul2_0_1_n65, SBOX_s5_mul2_0_1_n64,
         SBOX_s5_mul2_0_1_n63, SBOX_s5_mul2_0_1_n62, SBOX_s5_mul2_0_1_n61,
         SBOX_s5_mul2_0_1_n60, SBOX_s5_mul2_0_1_n59, SBOX_s5_mul2_0_1_n58,
         SBOX_s5_mul2_0_1_n57, SBOX_s5_mul2_0_1_n56, SBOX_s5_mul2_0_1_n55,
         SBOX_s5_mul2_0_1_n54, SBOX_s5_mul2_0_1_n53, SBOX_s5_mul2_0_0_n76,
         SBOX_s5_mul2_0_0_n75, SBOX_s5_mul2_0_0_n74, SBOX_s5_mul2_0_0_n73,
         SBOX_s5_mul2_0_0_n72, SBOX_s5_mul2_0_0_n71, SBOX_s5_mul2_0_0_n70,
         SBOX_s5_mul2_0_0_n69, SBOX_s5_mul2_0_0_n68, SBOX_s5_mul2_0_0_n67,
         SBOX_s5_mul2_0_0_n66, SBOX_s5_mul2_0_0_n65, SBOX_s5_mul2_0_0_n64,
         SBOX_s5_mul2_0_0_n63, SBOX_s5_mul2_0_0_n62, SBOX_s5_mul2_0_0_n61,
         SBOX_s5_mul2_0_0_n60, SBOX_s5_mul2_0_0_n59, SBOX_s5_mul2_0_0_n58,
         SBOX_s5_mul2_0_0_n57, SBOX_s5_mul2_0_0_n56, SBOX_s5_mul2_0_0_n55,
         SBOX_s5_mul2_0_0_n54, SBOX_s5_mul2_0_0_n53, SBOX_s6_1_n9,
         SBOX_s6_1_n8, SBOX_s6_1_n7, SBOX_s6_0_n9, SBOX_s6_0_n8, SBOX_s6_0_n7,
         aes_key_regs_1_n4, aes_key_regs_1_K02xDP_0_, aes_key_regs_1_K02xDP_1_,
         aes_key_regs_1_K02xDP_2_, aes_key_regs_1_K02xDP_3_,
         aes_key_regs_1_K02xDP_4_, aes_key_regs_1_K02xDP_5_,
         aes_key_regs_1_K02xDP_6_, aes_key_regs_1_K02xDP_7_,
         aes_key_regs_1_K01xDP_0_, aes_key_regs_1_K01xDP_1_,
         aes_key_regs_1_K01xDP_2_, aes_key_regs_1_K01xDP_3_,
         aes_key_regs_1_K01xDP_4_, aes_key_regs_1_K01xDP_5_,
         aes_key_regs_1_K01xDP_6_, aes_key_regs_1_K01xDP_7_,
         aes_state_regs_1_n112, aes_state_regs_1_n111, aes_state_regs_1_n110,
         aes_state_regs_1_n109, aes_state_regs_1_n108, aes_state_regs_1_n107,
         aes_state_regs_1_n106, aes_state_regs_1_n81, aes_state_regs_1_n80,
         aes_state_regs_1_n79, aes_state_regs_1_n78, aes_state_regs_1_n77,
         aes_state_regs_1_n76, aes_state_regs_1_n75, aes_state_regs_1_n74,
         aes_state_regs_1_n73, aes_state_regs_1_n72, aes_state_regs_1_n71,
         aes_state_regs_1_n70, aes_state_regs_1_n69, aes_state_regs_1_n68,
         aes_state_regs_1_n67, aes_state_regs_1_n66, aes_state_regs_1_n65,
         aes_state_regs_1_n64, aes_state_regs_1_n63, aes_state_regs_1_n56,
         aes_state_regs_1_n46, aes_state_regs_1_n45, aes_state_regs_1_n105,
         aes_state_regs_1_n104, aes_state_regs_1_n103, aes_state_regs_1_n102,
         aes_state_regs_1_n101, aes_state_regs_1_n100, aes_state_regs_1_n99,
         aes_state_regs_1_n98, aes_state_regs_1_n97, aes_state_regs_1_n96,
         aes_state_regs_1_n95, aes_state_regs_1_n94, aes_state_regs_1_n93,
         aes_state_regs_1_n92, aes_state_regs_1_n91, aes_state_regs_1_n90,
         aes_state_regs_1_n89, aes_state_regs_1_n88, aes_state_regs_1_n87,
         aes_state_regs_1_n86, aes_state_regs_1_n85, aes_state_regs_1_n84,
         aes_state_regs_1_n83, aes_state_regs_1_n82, aes_state_regs_1_n62,
         aes_state_regs_1_n61, aes_state_regs_1_n60, aes_state_regs_1_n59,
         aes_state_regs_1_n58, aes_state_regs_1_n57, aes_state_regs_1_n55,
         aes_state_regs_1_n54, aes_state_regs_1_n53, aes_state_regs_1_n52,
         aes_state_regs_1_n51, aes_state_regs_1_n50, aes_state_regs_1_n49,
         aes_state_regs_1_n48, aes_state_regs_1_n47, aes_state_regs_1_n38,
         aes_state_regs_1_n37, aes_state_regs_1_n36, aes_state_regs_1_n35,
         aes_state_regs_1_n34, aes_state_regs_1_n33, aes_state_regs_1_n32,
         aes_state_regs_1_n31, aes_state_regs_1_n30, aes_state_regs_1_n29,
         aes_state_regs_1_n28, aes_state_regs_1_n27, aes_state_regs_1_n26,
         aes_state_regs_1_n25, aes_state_regs_1_n24, aes_state_regs_1_n23,
         aes_state_regs_1_n22, aes_state_regs_1_n21, aes_state_regs_1_n20,
         aes_state_regs_1_n19, aes_state_regs_1_n18, aes_state_regs_1_n17,
         aes_state_regs_1_n16, aes_state_regs_1_n15, aes_state_regs_1_n14,
         aes_state_regs_1_n13, aes_state_regs_1_n12, aes_state_regs_1_n11,
         aes_state_regs_1_n10, aes_state_regs_1_n9, aes_state_regs_1_n8,
         aes_state_regs_1_n7, aes_state_regs_1_n6, aes_state_regs_1_n5,
         aes_state_regs_1_n4, aes_state_regs_1_n3, aes_state_regs_1_n2,
         aes_state_regs_1_n1, aes_state_regs_1_S03xDP_0_,
         aes_state_regs_1_S02xDP_0_, aes_state_regs_1_S02xDP_1_,
         aes_state_regs_1_S02xDP_2_, aes_state_regs_1_S02xDP_3_,
         aes_state_regs_1_S02xDP_4_, aes_state_regs_1_S02xDP_5_,
         aes_state_regs_1_S02xDP_6_, aes_state_regs_1_S02xDP_7_,
         aes_state_regs_1_S31xDP_0_, aes_state_regs_1_S30xDP_0_,
         aes_state_regs_1_S30xDP_1_, aes_state_regs_1_S30xDP_2_,
         aes_state_regs_1_S30xDP_3_, aes_state_regs_1_S30xDP_4_,
         aes_state_regs_1_S30xDP_5_, aes_state_regs_1_S30xDP_6_,
         aes_state_regs_1_S30xDP_7_, aes_state_regs_1_S20xDP_0_,
         aes_state_regs_1_S20xDP_1_, aes_state_regs_1_S20xDP_2_,
         aes_state_regs_1_S20xDP_3_, aes_state_regs_1_S20xDP_4_,
         aes_state_regs_1_S20xDP_5_, aes_state_regs_1_S20xDP_6_,
         aes_state_regs_1_S20xDP_7_, aes_state_regs_1_S23xDP_0_,
         aes_state_regs_1_S23xDP_1_, aes_state_regs_1_S23xDP_2_,
         aes_state_regs_1_S23xDP_3_, aes_state_regs_1_S23xDP_4_,
         aes_state_regs_1_S23xDP_5_, aes_state_regs_1_S23xDP_6_,
         aes_state_regs_1_S23xDP_7_, aes_state_regs_1_S22xDP_0_,
         aes_state_regs_1_S10xDP_0_, aes_state_regs_1_S10xDP_1_,
         aes_state_regs_1_S10xDP_2_, aes_state_regs_1_S10xDP_3_,
         aes_state_regs_1_S10xDP_4_, aes_state_regs_1_S10xDP_5_,
         aes_state_regs_1_S10xDP_6_, aes_state_regs_1_S10xDP_7_,
         aes_state_regs_1_S01xDO_0_, aes_state_regs_1_S01xDO_1_,
         aes_state_regs_1_S01xDO_2_, aes_state_regs_1_S01xDO_3_,
         aes_state_regs_1_S01xDO_4_, aes_state_regs_1_S01xDO_5_,
         aes_state_regs_1_S01xDO_6_, aes_state_regs_1_S01xDO_7_,
         aes_state_regs_1_mix_columns_1_n245,
         aes_state_regs_1_mix_columns_1_n244,
         aes_state_regs_1_mix_columns_1_n243,
         aes_state_regs_1_mix_columns_1_n242,
         aes_state_regs_1_mix_columns_1_n241,
         aes_state_regs_1_mix_columns_1_n240,
         aes_state_regs_1_mix_columns_1_n239,
         aes_state_regs_1_mix_columns_1_n238,
         aes_state_regs_1_mix_columns_1_n237,
         aes_state_regs_1_mix_columns_1_n236,
         aes_state_regs_1_mix_columns_1_n235,
         aes_state_regs_1_mix_columns_1_n234,
         aes_state_regs_1_mix_columns_1_n233,
         aes_state_regs_1_mix_columns_1_n232,
         aes_state_regs_1_mix_columns_1_n231,
         aes_state_regs_1_mix_columns_1_n230,
         aes_state_regs_1_mix_columns_1_n229,
         aes_state_regs_1_mix_columns_1_n228,
         aes_state_regs_1_mix_columns_1_n227,
         aes_state_regs_1_mix_columns_1_n226,
         aes_state_regs_1_mix_columns_1_n225,
         aes_state_regs_1_mix_columns_1_n224,
         aes_state_regs_1_mix_columns_1_n223,
         aes_state_regs_1_mix_columns_1_n222,
         aes_state_regs_1_mix_columns_1_n221,
         aes_state_regs_1_mix_columns_1_n220,
         aes_state_regs_1_mix_columns_1_n219,
         aes_state_regs_1_mix_columns_1_n218,
         aes_state_regs_1_mix_columns_1_n217,
         aes_state_regs_1_mix_columns_1_n216,
         aes_state_regs_1_mix_columns_1_n215,
         aes_state_regs_1_mix_columns_1_n214,
         aes_state_regs_1_mix_columns_1_n213,
         aes_state_regs_1_mix_columns_1_n212,
         aes_state_regs_1_mix_columns_1_n211,
         aes_state_regs_1_mix_columns_1_n210,
         aes_state_regs_1_mix_columns_1_n209,
         aes_state_regs_1_mix_columns_1_n208,
         aes_state_regs_1_mix_columns_1_n207,
         aes_state_regs_1_mix_columns_1_n206,
         aes_state_regs_1_mix_columns_1_n205,
         aes_state_regs_1_mix_columns_1_n204,
         aes_state_regs_1_mix_columns_1_n203,
         aes_state_regs_1_mix_columns_1_n202,
         aes_state_regs_1_mix_columns_1_n201,
         aes_state_regs_1_mix_columns_1_n200,
         aes_state_regs_1_mix_columns_1_n199,
         aes_state_regs_1_mix_columns_1_n198,
         aes_state_regs_1_mix_columns_1_n197,
         aes_state_regs_1_mix_columns_1_n196,
         aes_state_regs_1_mix_columns_1_n195,
         aes_state_regs_1_mix_columns_1_n194,
         aes_state_regs_1_mix_columns_1_n193,
         aes_state_regs_1_mix_columns_1_n192,
         aes_state_regs_1_mix_columns_1_n191,
         aes_state_regs_1_mix_columns_1_n190,
         aes_state_regs_1_mix_columns_1_n189,
         aes_state_regs_1_mix_columns_1_n188,
         aes_state_regs_1_mix_columns_1_n187,
         aes_state_regs_1_mix_columns_1_n186,
         aes_state_regs_1_mix_columns_1_n185,
         aes_state_regs_1_mix_columns_1_n184,
         aes_state_regs_1_mix_columns_1_n183,
         aes_state_regs_1_mix_columns_1_n182,
         aes_state_regs_1_mix_columns_1_n181,
         aes_state_regs_1_mix_columns_1_n180,
         aes_state_regs_1_mix_columns_1_n179,
         aes_state_regs_1_mix_columns_1_n178,
         aes_state_regs_1_mix_columns_1_n177,
         aes_state_regs_1_mix_columns_1_n176,
         aes_state_regs_1_mix_columns_1_n175,
         aes_state_regs_1_mix_columns_1_n174,
         aes_state_regs_1_mix_columns_1_n173,
         aes_state_regs_1_mix_columns_1_n172,
         aes_state_regs_1_mix_columns_1_n171,
         aes_state_regs_1_mix_columns_1_n170,
         aes_state_regs_1_mix_columns_1_n169,
         aes_state_regs_1_mix_columns_1_n168,
         aes_state_regs_1_mix_columns_1_n167,
         aes_state_regs_1_mix_columns_1_n166,
         aes_state_regs_1_mix_columns_1_n165,
         aes_state_regs_1_mix_columns_1_n164,
         aes_state_regs_1_mix_columns_1_n163,
         aes_state_regs_1_mix_columns_1_n162,
         aes_state_regs_1_mix_columns_1_n161,
         aes_state_regs_1_mix_columns_1_n160,
         aes_state_regs_1_mix_columns_1_n159, aes_key_regs_0_n4,
         aes_key_regs_0_K02xDP_0_, aes_key_regs_0_K02xDP_1_,
         aes_key_regs_0_K02xDP_2_, aes_key_regs_0_K02xDP_3_,
         aes_key_regs_0_K02xDP_4_, aes_key_regs_0_K02xDP_5_,
         aes_key_regs_0_K02xDP_6_, aes_key_regs_0_K02xDP_7_,
         aes_key_regs_0_K01xDP_0_, aes_key_regs_0_K01xDP_1_,
         aes_key_regs_0_K01xDP_2_, aes_key_regs_0_K01xDP_3_,
         aes_key_regs_0_K01xDP_4_, aes_key_regs_0_K01xDP_5_,
         aes_key_regs_0_K01xDP_6_, aes_key_regs_0_K01xDP_7_,
         aes_state_regs_0_n202, aes_state_regs_0_n201, aes_state_regs_0_n200,
         aes_state_regs_0_n199, aes_state_regs_0_n198, aes_state_regs_0_n197,
         aes_state_regs_0_n196, aes_state_regs_0_n195, aes_state_regs_0_n194,
         aes_state_regs_0_n193, aes_state_regs_0_n192, aes_state_regs_0_n191,
         aes_state_regs_0_n190, aes_state_regs_0_n189, aes_state_regs_0_n188,
         aes_state_regs_0_n187, aes_state_regs_0_n186, aes_state_regs_0_n185,
         aes_state_regs_0_n184, aes_state_regs_0_n183, aes_state_regs_0_n182,
         aes_state_regs_0_n181, aes_state_regs_0_n180, aes_state_regs_0_n179,
         aes_state_regs_0_n178, aes_state_regs_0_n177, aes_state_regs_0_n176,
         aes_state_regs_0_n175, aes_state_regs_0_n174, aes_state_regs_0_n51,
         aes_state_regs_0_n50, aes_state_regs_0_n49, aes_state_regs_0_n48,
         aes_state_regs_0_n47, aes_state_regs_0_n46, aes_state_regs_0_n45,
         aes_state_regs_0_n44, aes_state_regs_0_n43, aes_state_regs_0_n42,
         aes_state_regs_0_n41, aes_state_regs_0_n40, aes_state_regs_0_n39,
         aes_state_regs_0_n38, aes_state_regs_0_n37, aes_state_regs_0_n36,
         aes_state_regs_0_n35, aes_state_regs_0_n34, aes_state_regs_0_n33,
         aes_state_regs_0_n32, aes_state_regs_0_n31, aes_state_regs_0_n30,
         aes_state_regs_0_n29, aes_state_regs_0_n28, aes_state_regs_0_n173,
         aes_state_regs_0_n172, aes_state_regs_0_n171, aes_state_regs_0_n170,
         aes_state_regs_0_n169, aes_state_regs_0_n168, aes_state_regs_0_n167,
         aes_state_regs_0_n166, aes_state_regs_0_n165, aes_state_regs_0_n164,
         aes_state_regs_0_n163, aes_state_regs_0_n162, aes_state_regs_0_n161,
         aes_state_regs_0_n160, aes_state_regs_0_n159, aes_state_regs_0_n158,
         aes_state_regs_0_n157, aes_state_regs_0_n156, aes_state_regs_0_n155,
         aes_state_regs_0_n154, aes_state_regs_0_n153, aes_state_regs_0_n152,
         aes_state_regs_0_n151, aes_state_regs_0_n150, aes_state_regs_0_n149,
         aes_state_regs_0_n148, aes_state_regs_0_n147, aes_state_regs_0_n146,
         aes_state_regs_0_n145, aes_state_regs_0_n144, aes_state_regs_0_n143,
         aes_state_regs_0_n142, aes_state_regs_0_n141, aes_state_regs_0_n140,
         aes_state_regs_0_n139, aes_state_regs_0_n138, aes_state_regs_0_n137,
         aes_state_regs_0_n136, aes_state_regs_0_n127, aes_state_regs_0_n126,
         aes_state_regs_0_n125, aes_state_regs_0_n124, aes_state_regs_0_n123,
         aes_state_regs_0_n122, aes_state_regs_0_n121, aes_state_regs_0_n109,
         aes_state_regs_0_S03xDP_0_, aes_state_regs_0_S02xDP_0_,
         aes_state_regs_0_S02xDP_1_, aes_state_regs_0_S02xDP_2_,
         aes_state_regs_0_S02xDP_3_, aes_state_regs_0_S02xDP_4_,
         aes_state_regs_0_S02xDP_5_, aes_state_regs_0_S02xDP_6_,
         aes_state_regs_0_S02xDP_7_, aes_state_regs_0_S31xDP_0_,
         aes_state_regs_0_S30xDP_0_, aes_state_regs_0_S30xDP_1_,
         aes_state_regs_0_S30xDP_2_, aes_state_regs_0_S30xDP_3_,
         aes_state_regs_0_S30xDP_4_, aes_state_regs_0_S30xDP_5_,
         aes_state_regs_0_S30xDP_6_, aes_state_regs_0_S30xDP_7_,
         aes_state_regs_0_S20xDP_0_, aes_state_regs_0_S20xDP_1_,
         aes_state_regs_0_S20xDP_2_, aes_state_regs_0_S20xDP_3_,
         aes_state_regs_0_S20xDP_4_, aes_state_regs_0_S20xDP_5_,
         aes_state_regs_0_S20xDP_6_, aes_state_regs_0_S20xDP_7_,
         aes_state_regs_0_S23xDP_0_, aes_state_regs_0_S23xDP_1_,
         aes_state_regs_0_S23xDP_2_, aes_state_regs_0_S23xDP_3_,
         aes_state_regs_0_S23xDP_4_, aes_state_regs_0_S23xDP_5_,
         aes_state_regs_0_S23xDP_6_, aes_state_regs_0_S23xDP_7_,
         aes_state_regs_0_S22xDP_0_, aes_state_regs_0_S10xDP_0_,
         aes_state_regs_0_S10xDP_1_, aes_state_regs_0_S10xDP_2_,
         aes_state_regs_0_S10xDP_3_, aes_state_regs_0_S10xDP_4_,
         aes_state_regs_0_S10xDP_5_, aes_state_regs_0_S10xDP_6_,
         aes_state_regs_0_S10xDP_7_, aes_state_regs_0_S01xDO_0_,
         aes_state_regs_0_S01xDO_1_, aes_state_regs_0_S01xDO_2_,
         aes_state_regs_0_S01xDO_3_, aes_state_regs_0_S01xDO_4_,
         aes_state_regs_0_S01xDO_5_, aes_state_regs_0_S01xDO_6_,
         aes_state_regs_0_S01xDO_7_, aes_state_regs_0_mix_columns_1_n245,
         aes_state_regs_0_mix_columns_1_n244,
         aes_state_regs_0_mix_columns_1_n243,
         aes_state_regs_0_mix_columns_1_n242,
         aes_state_regs_0_mix_columns_1_n241,
         aes_state_regs_0_mix_columns_1_n240,
         aes_state_regs_0_mix_columns_1_n239,
         aes_state_regs_0_mix_columns_1_n238,
         aes_state_regs_0_mix_columns_1_n237,
         aes_state_regs_0_mix_columns_1_n236,
         aes_state_regs_0_mix_columns_1_n235,
         aes_state_regs_0_mix_columns_1_n234,
         aes_state_regs_0_mix_columns_1_n233,
         aes_state_regs_0_mix_columns_1_n232,
         aes_state_regs_0_mix_columns_1_n231,
         aes_state_regs_0_mix_columns_1_n230,
         aes_state_regs_0_mix_columns_1_n229,
         aes_state_regs_0_mix_columns_1_n228,
         aes_state_regs_0_mix_columns_1_n227,
         aes_state_regs_0_mix_columns_1_n226,
         aes_state_regs_0_mix_columns_1_n225,
         aes_state_regs_0_mix_columns_1_n224,
         aes_state_regs_0_mix_columns_1_n223,
         aes_state_regs_0_mix_columns_1_n222,
         aes_state_regs_0_mix_columns_1_n221,
         aes_state_regs_0_mix_columns_1_n220,
         aes_state_regs_0_mix_columns_1_n219,
         aes_state_regs_0_mix_columns_1_n218,
         aes_state_regs_0_mix_columns_1_n217,
         aes_state_regs_0_mix_columns_1_n216,
         aes_state_regs_0_mix_columns_1_n215,
         aes_state_regs_0_mix_columns_1_n214,
         aes_state_regs_0_mix_columns_1_n213,
         aes_state_regs_0_mix_columns_1_n212,
         aes_state_regs_0_mix_columns_1_n211,
         aes_state_regs_0_mix_columns_1_n210,
         aes_state_regs_0_mix_columns_1_n209,
         aes_state_regs_0_mix_columns_1_n208,
         aes_state_regs_0_mix_columns_1_n207,
         aes_state_regs_0_mix_columns_1_n206,
         aes_state_regs_0_mix_columns_1_n205,
         aes_state_regs_0_mix_columns_1_n204,
         aes_state_regs_0_mix_columns_1_n203,
         aes_state_regs_0_mix_columns_1_n202,
         aes_state_regs_0_mix_columns_1_n201,
         aes_state_regs_0_mix_columns_1_n200,
         aes_state_regs_0_mix_columns_1_n199,
         aes_state_regs_0_mix_columns_1_n198,
         aes_state_regs_0_mix_columns_1_n197,
         aes_state_regs_0_mix_columns_1_n196,
         aes_state_regs_0_mix_columns_1_n195,
         aes_state_regs_0_mix_columns_1_n194,
         aes_state_regs_0_mix_columns_1_n193,
         aes_state_regs_0_mix_columns_1_n192,
         aes_state_regs_0_mix_columns_1_n191,
         aes_state_regs_0_mix_columns_1_n190,
         aes_state_regs_0_mix_columns_1_n189,
         aes_state_regs_0_mix_columns_1_n188,
         aes_state_regs_0_mix_columns_1_n187,
         aes_state_regs_0_mix_columns_1_n186,
         aes_state_regs_0_mix_columns_1_n185,
         aes_state_regs_0_mix_columns_1_n184,
         aes_state_regs_0_mix_columns_1_n183,
         aes_state_regs_0_mix_columns_1_n182,
         aes_state_regs_0_mix_columns_1_n181,
         aes_state_regs_0_mix_columns_1_n180,
         aes_state_regs_0_mix_columns_1_n179,
         aes_state_regs_0_mix_columns_1_n178,
         aes_state_regs_0_mix_columns_1_n177,
         aes_state_regs_0_mix_columns_1_n176,
         aes_state_regs_0_mix_columns_1_n175,
         aes_state_regs_0_mix_columns_1_n174,
         aes_state_regs_0_mix_columns_1_n173,
         aes_state_regs_0_mix_columns_1_n172,
         aes_state_regs_0_mix_columns_1_n171,
         aes_state_regs_0_mix_columns_1_n170,
         aes_state_regs_0_mix_columns_1_n169,
         aes_state_regs_0_mix_columns_1_n168,
         aes_state_regs_0_mix_columns_1_n167,
         aes_state_regs_0_mix_columns_1_n166,
         aes_state_regs_0_mix_columns_1_n165,
         aes_state_regs_0_mix_columns_1_n164,
         aes_state_regs_0_mix_columns_1_n163,
         aes_state_regs_0_mix_columns_1_n162,
         aes_state_regs_0_mix_columns_1_n161,
         aes_state_regs_0_mix_columns_1_n160,
         aes_state_regs_0_mix_columns_1_n159;
  wire   [15:0] KeyToSboxOutxD;
  wire   [15:0] KeyInxD;
  wire   [15:0] StateOutxD;
  wire   [15:0] StateInxD;
  wire   [15:0] KeyOutxD;
  wire   [15:0] K03xD;
  wire   [7:0] RCONxD;
  wire   [15:0] SBOX_regOut1;
  wire   [15:0] SBOX_stage6Out;
  wire   [15:0] SBOX_stage5Out;
  wire   [23:0] SBOX_stage4Out;
  wire   [23:0] SBOX_stage3Out;
  wire   [23:0] SBOX_stage2Out;
  wire   [15:0] SBOX_stage1Out;
  wire   [15:0] SBOX_s2_refreshed;
  wire   [7:0] SBOX_s2_xorResult;
  wire   [7:0] SBOX_s2_sqsc_out;
  wire   [5:0] SBOX_s2_sqsc_in;
  wire   [7:0] SBOX_s3_refreshed;
  wire   [3:0] SBOX_s3_xorResult;
  wire   [3:0] SBOX_s3_scale_out;
  wire   [1:0] SBOX_s3_scale_in;
  wire   [15:0] SBOX_s4_refreshed;
  wire   [15:0] SBOX_s4_concat;
  wire   [31:0] SBOX_s5_regOut;
  wire   [31:0] SBOX_s5_refreshed;
  wire   [31:0] SBOX_s5_concat;
  wire   [7:0] aes_key_regs_1_K23xDN;
  wire   [7:0] aes_key_regs_1_K22xDN;
  wire   [7:0] aes_key_regs_1_K21xDN;
  wire   [7:0] aes_key_regs_1_K20xDN;
  wire   [7:0] aes_key_regs_1_K13xDN;
  wire   [7:0] aes_key_regs_1_K12xDN;
  wire   [7:0] aes_key_regs_1_K11xDN;
  wire   [7:0] aes_key_regs_1_K10xDN;
  wire   [7:0] aes_key_regs_1_K02xDN;
  wire   [7:0] aes_key_regs_1_K01xDN;
  wire   [7:0] aes_key_regs_1_K00xDN;
  wire   [7:0] aes_state_regs_1_MixColumnsS3xD;
  wire   [7:0] aes_state_regs_1_MixColumnsS2xD;
  wire   [7:0] aes_state_regs_1_MixColumnsS1xD;
  wire   [7:0] aes_state_regs_1_MixColumnsS0xD;
  wire   [7:0] aes_state_regs_1_S20xDN;
  wire   [7:1] aes_state_regs_1_S21xDP;
  wire   [7:0] aes_state_regs_1_S10xDN;
  wire   [7:0] aes_state_regs_1_S03xDN;
  wire   [7:0] aes_state_regs_1_S02xDN;
  wire   [7:0] aes_state_regs_1_S01xDN;
  wire   [7:0] aes_state_regs_1_S00xDP;
  wire   [7:0] aes_key_regs_0_K23xDN;
  wire   [7:0] aes_key_regs_0_K22xDN;
  wire   [7:0] aes_key_regs_0_K21xDN;
  wire   [7:0] aes_key_regs_0_K20xDN;
  wire   [7:0] aes_key_regs_0_K13xDN;
  wire   [7:0] aes_key_regs_0_K12xDN;
  wire   [7:0] aes_key_regs_0_K11xDN;
  wire   [7:0] aes_key_regs_0_K10xDN;
  wire   [7:0] aes_key_regs_0_K02xDN;
  wire   [7:0] aes_key_regs_0_K01xDN;
  wire   [7:0] aes_key_regs_0_K00xDN;
  wire   [7:0] aes_state_regs_0_MixColumnsS3xD;
  wire   [7:0] aes_state_regs_0_MixColumnsS2xD;
  wire   [7:0] aes_state_regs_0_MixColumnsS1xD;
  wire   [7:0] aes_state_regs_0_MixColumnsS0xD;
  wire   [7:0] aes_state_regs_0_S20xDN;
  wire   [7:1] aes_state_regs_0_S21xDP;
  wire   [7:0] aes_state_regs_0_S10xDN;
  wire   [7:0] aes_state_regs_0_S03xDN;
  wire   [7:0] aes_state_regs_0_S02xDN;
  wire   [7:0] aes_state_regs_0_S01xDN;
  wire   [7:0] aes_state_regs_0_S00xDP;

  DFFS_X1 disableKeyRegsxSP_reg ( .D(disableKeyRegsxS), .CK(ClkxCI), .SN(
        RstxBI), .Q(n226), .QN() );
  OAI22_X1 U296 ( .A1(StateOutxD[13]), .A2(n338), .B1(PTxDI[13]), .B2(n337), 
        .ZN(n325) );
  OAI22_X1 U297 ( .A1(StateOutxD[14]), .A2(n338), .B1(PTxDI[14]), .B2(n337), 
        .ZN(n330) );
  INV_X1 U298 ( .A(n336), .ZN(n338) );
  NAND2_X1 U299 ( .A1(FinishedxS), .A2(n260), .ZN(n337) );
  INV_X1 U300 ( .A(n337), .ZN(n335) );
  NOR2_X1 U301 ( .A1(StateKEYSCHEDULExS), .A2(nextRCONxS), .ZN(n260) );
  OAI22_X1 U302 ( .A1(K03xD[13]), .A2(n334), .B1(StateInxD[13]), .B2(n333), 
        .ZN(n324) );
  AOI22_X1 U303 ( .A1(FinishedxS), .A2(KxDI[14]), .B1(KeyOutxD[14]), .B2(n328), 
        .ZN(n329) );
  OAI22_X1 U304 ( .A1(K03xD[14]), .A2(n334), .B1(StateInxD[14]), .B2(n333), 
        .ZN(n328) );
  INV_X1 U305 ( .A(n332), .ZN(n334) );
  NOR2_X1 U306 ( .A1(FinishedxS), .A2(n255), .ZN(n331) );
  INV_X1 U307 ( .A(StateKEYADDITION1o3xS), .ZN(n255) );
  INV_X1 U308 ( .A(n331), .ZN(n333) );
  OAI21_X1 U309 ( .B1(n270), .B2(KeyInxD[1]), .A(n269), .ZN(CxDO[1]) );
  OAI22_X1 U310 ( .A1(StateOutxD[1]), .A2(n338), .B1(PTxDI[1]), .B2(n337), 
        .ZN(n268) );
  OAI21_X1 U311 ( .B1(n277), .B2(KeyInxD[2]), .A(n276), .ZN(CxDO[2]) );
  AOI22_X1 U312 ( .A1(KeyToSboxOutxD[2]), .A2(n114), .B1(n275), .B2(KeyInxD[2]), .ZN(n276) );
  OAI22_X1 U313 ( .A1(StateOutxD[2]), .A2(n338), .B1(PTxDI[2]), .B2(n337), 
        .ZN(n275) );
  OAI21_X1 U314 ( .B1(n284), .B2(KeyInxD[3]), .A(n283), .ZN(CxDO[3]) );
  AOI22_X1 U315 ( .A1(n336), .A2(StateOutxD[3]), .B1(n335), .B2(PTxDI[3]), 
        .ZN(n284) );
  AOI22_X1 U316 ( .A1(KeyToSboxOutxD[3]), .A2(n114), .B1(n282), .B2(KeyInxD[3]), .ZN(n283) );
  OAI22_X1 U317 ( .A1(StateOutxD[3]), .A2(n338), .B1(PTxDI[3]), .B2(n337), 
        .ZN(n282) );
  OAI21_X1 U318 ( .B1(n291), .B2(KeyInxD[4]), .A(n290), .ZN(CxDO[4]) );
  AOI22_X1 U319 ( .A1(KeyToSboxOutxD[4]), .A2(n114), .B1(n289), .B2(KeyInxD[4]), .ZN(n290) );
  OAI22_X1 U320 ( .A1(StateOutxD[4]), .A2(n338), .B1(PTxDI[4]), .B2(n337), 
        .ZN(n289) );
  OAI21_X1 U321 ( .B1(n298), .B2(KeyInxD[5]), .A(n297), .ZN(CxDO[5]) );
  AOI22_X1 U322 ( .A1(n336), .A2(StateOutxD[5]), .B1(n335), .B2(PTxDI[5]), 
        .ZN(n298) );
  AOI22_X1 U323 ( .A1(KeyToSboxOutxD[5]), .A2(n114), .B1(n296), .B2(KeyInxD[5]), .ZN(n297) );
  OAI22_X1 U324 ( .A1(StateOutxD[5]), .A2(n338), .B1(PTxDI[5]), .B2(n337), 
        .ZN(n296) );
  OAI21_X1 U325 ( .B1(n305), .B2(KeyInxD[6]), .A(n304), .ZN(CxDO[6]) );
  AOI22_X1 U326 ( .A1(KeyToSboxOutxD[6]), .A2(n114), .B1(n303), .B2(KeyInxD[6]), .ZN(n304) );
  OAI22_X1 U327 ( .A1(StateOutxD[6]), .A2(n338), .B1(PTxDI[6]), .B2(n337), 
        .ZN(n303) );
  OAI21_X1 U328 ( .B1(n308), .B2(KeyInxD[7]), .A(n307), .ZN(CxDO[7]) );
  AOI22_X1 U329 ( .A1(KeyToSboxOutxD[7]), .A2(n114), .B1(n306), .B2(KeyInxD[7]), .ZN(n307) );
  OAI22_X1 U330 ( .A1(StateOutxD[7]), .A2(n338), .B1(PTxDI[7]), .B2(n337), 
        .ZN(n306) );
  OAI21_X1 U331 ( .B1(n314), .B2(KeyInxD[9]), .A(n313), .ZN(CxDO[9]) );
  AOI22_X1 U332 ( .A1(n336), .A2(StateOutxD[9]), .B1(n335), .B2(PTxDI[9]), 
        .ZN(n314) );
  AOI22_X1 U333 ( .A1(KeyToSboxOutxD[9]), .A2(n114), .B1(n312), .B2(KeyInxD[9]), .ZN(n313) );
  OAI22_X1 U334 ( .A1(StateOutxD[9]), .A2(n338), .B1(PTxDI[9]), .B2(n337), 
        .ZN(n312) );
  OAI21_X1 U335 ( .B1(n317), .B2(KeyInxD[10]), .A(n316), .ZN(CxDO[10]) );
  AOI22_X1 U336 ( .A1(n336), .A2(StateOutxD[10]), .B1(n335), .B2(PTxDI[10]), 
        .ZN(n317) );
  AOI22_X1 U337 ( .A1(KeyToSboxOutxD[10]), .A2(n114), .B1(n315), .B2(
        KeyInxD[10]), .ZN(n316) );
  OAI22_X1 U338 ( .A1(StateOutxD[10]), .A2(n338), .B1(PTxDI[10]), .B2(n337), 
        .ZN(n315) );
  OAI21_X1 U339 ( .B1(n320), .B2(KeyInxD[11]), .A(n319), .ZN(CxDO[11]) );
  AOI22_X1 U340 ( .A1(n336), .A2(StateOutxD[11]), .B1(n335), .B2(PTxDI[11]), 
        .ZN(n320) );
  AOI22_X1 U341 ( .A1(KeyToSboxOutxD[11]), .A2(n114), .B1(n318), .B2(
        KeyInxD[11]), .ZN(n319) );
  OAI22_X1 U342 ( .A1(StateOutxD[11]), .A2(n338), .B1(PTxDI[11]), .B2(n337), 
        .ZN(n318) );
  OAI21_X1 U343 ( .B1(n323), .B2(KeyInxD[12]), .A(n322), .ZN(CxDO[12]) );
  AOI22_X1 U344 ( .A1(n336), .A2(StateOutxD[12]), .B1(n335), .B2(PTxDI[12]), 
        .ZN(n323) );
  AOI22_X1 U345 ( .A1(KeyToSboxOutxD[12]), .A2(n114), .B1(n321), .B2(
        KeyInxD[12]), .ZN(n322) );
  OAI22_X1 U346 ( .A1(StateOutxD[12]), .A2(n338), .B1(PTxDI[12]), .B2(n337), 
        .ZN(n321) );
  OAI21_X1 U347 ( .B1(n327), .B2(KeyInxD[13]), .A(n326), .ZN(CxDO[13]) );
  AOI22_X1 U348 ( .A1(n336), .A2(StateOutxD[13]), .B1(n335), .B2(PTxDI[13]), 
        .ZN(n327) );
  AOI22_X1 U349 ( .A1(KeyToSboxOutxD[13]), .A2(n114), .B1(n325), .B2(
        KeyInxD[13]), .ZN(n326) );
  OAI21_X1 U350 ( .B1(n341), .B2(KeyInxD[15]), .A(n340), .ZN(CxDO[15]) );
  AOI22_X1 U351 ( .A1(n336), .A2(StateOutxD[15]), .B1(n335), .B2(PTxDI[15]), 
        .ZN(n341) );
  AOI22_X1 U352 ( .A1(KeyToSboxOutxD[15]), .A2(n114), .B1(n339), .B2(
        KeyInxD[15]), .ZN(n340) );
  OAI22_X1 U353 ( .A1(StateOutxD[15]), .A2(n338), .B1(PTxDI[15]), .B2(n337), 
        .ZN(n339) );
  AND2_X1 U354 ( .A1(LastRoundxS), .A2(showRCONxS), .ZN(DonexSO) );
  OAI21_X1 U355 ( .B1(n263), .B2(KeyInxD[0]), .A(n262), .ZN(CxDO[0]) );
  AOI22_X1 U356 ( .A1(KeyToSboxOutxD[0]), .A2(n114), .B1(n261), .B2(KeyInxD[0]), .ZN(n262) );
  OAI22_X1 U357 ( .A1(StateOutxD[0]), .A2(n338), .B1(PTxDI[0]), .B2(n337), 
        .ZN(n261) );
  OAI21_X1 U358 ( .B1(n311), .B2(KeyInxD[8]), .A(n310), .ZN(CxDO[8]) );
  AOI22_X1 U359 ( .A1(n336), .A2(StateOutxD[8]), .B1(n335), .B2(PTxDI[8]), 
        .ZN(n311) );
  AOI22_X1 U360 ( .A1(KeyToSboxOutxD[8]), .A2(n114), .B1(n309), .B2(KeyInxD[8]), .ZN(n310) );
  OAI22_X1 U361 ( .A1(StateOutxD[8]), .A2(n338), .B1(PTxDI[8]), .B2(n337), 
        .ZN(n309) );
  OAI21_X1 U362 ( .B1(n333), .B2(n259), .A(n258), .ZN(KeyInxD[0]) );
  XNOR2_X1 U363 ( .A(StateInxD[0]), .B(n256), .ZN(n259) );
  AOI22_X1 U364 ( .A1(FinishedxS), .A2(KxDI[0]), .B1(n332), .B2(n257), .ZN(
        n258) );
  XOR2_X1 U365 ( .A(KeyOutxD[0]), .B(RCONxD[0]), .Z(n256) );
  XOR2_X1 U366 ( .A(KeyOutxD[0]), .B(K03xD[0]), .Z(n257) );
  OAI21_X1 U367 ( .B1(n333), .B2(n267), .A(n266), .ZN(KeyInxD[1]) );
  XNOR2_X1 U368 ( .A(StateInxD[1]), .B(n264), .ZN(n267) );
  AOI22_X1 U369 ( .A1(FinishedxS), .A2(KxDI[1]), .B1(n332), .B2(n265), .ZN(
        n266) );
  XOR2_X1 U370 ( .A(KeyOutxD[1]), .B(RCONxD[1]), .Z(n264) );
  XOR2_X1 U371 ( .A(KeyOutxD[1]), .B(K03xD[1]), .Z(n265) );
  OAI21_X1 U372 ( .B1(n333), .B2(n274), .A(n273), .ZN(KeyInxD[2]) );
  XNOR2_X1 U373 ( .A(StateInxD[2]), .B(n271), .ZN(n274) );
  AOI22_X1 U374 ( .A1(FinishedxS), .A2(KxDI[2]), .B1(n332), .B2(n272), .ZN(
        n273) );
  XOR2_X1 U375 ( .A(KeyOutxD[2]), .B(RCONxD[2]), .Z(n271) );
  XOR2_X1 U376 ( .A(KeyOutxD[2]), .B(K03xD[2]), .Z(n272) );
  OAI21_X1 U377 ( .B1(n333), .B2(n281), .A(n280), .ZN(KeyInxD[3]) );
  XNOR2_X1 U378 ( .A(StateInxD[3]), .B(n278), .ZN(n281) );
  AOI22_X1 U379 ( .A1(FinishedxS), .A2(KxDI[3]), .B1(n332), .B2(n279), .ZN(
        n280) );
  XOR2_X1 U380 ( .A(KeyOutxD[3]), .B(RCONxD[3]), .Z(n278) );
  XOR2_X1 U381 ( .A(KeyOutxD[3]), .B(K03xD[3]), .Z(n279) );
  OAI21_X1 U382 ( .B1(n333), .B2(n288), .A(n287), .ZN(KeyInxD[4]) );
  XNOR2_X1 U383 ( .A(StateInxD[4]), .B(n285), .ZN(n288) );
  AOI22_X1 U384 ( .A1(FinishedxS), .A2(KxDI[4]), .B1(n332), .B2(n286), .ZN(
        n287) );
  XOR2_X1 U385 ( .A(KeyOutxD[4]), .B(RCONxD[4]), .Z(n285) );
  XOR2_X1 U386 ( .A(KeyOutxD[4]), .B(K03xD[4]), .Z(n286) );
  OAI21_X1 U387 ( .B1(n333), .B2(n295), .A(n294), .ZN(KeyInxD[5]) );
  XNOR2_X1 U388 ( .A(StateInxD[5]), .B(n292), .ZN(n295) );
  AOI22_X1 U389 ( .A1(FinishedxS), .A2(KxDI[5]), .B1(n332), .B2(n293), .ZN(
        n294) );
  XOR2_X1 U390 ( .A(KeyOutxD[5]), .B(RCONxD[5]), .Z(n292) );
  XOR2_X1 U391 ( .A(KeyOutxD[5]), .B(K03xD[5]), .Z(n293) );
  OAI21_X1 U392 ( .B1(n333), .B2(n302), .A(n301), .ZN(KeyInxD[6]) );
  XNOR2_X1 U393 ( .A(StateInxD[6]), .B(n299), .ZN(n302) );
  AOI22_X1 U394 ( .A1(FinishedxS), .A2(KxDI[6]), .B1(n332), .B2(n300), .ZN(
        n301) );
  XOR2_X1 U395 ( .A(KeyOutxD[6]), .B(RCONxD[6]), .Z(n299) );
  XOR2_X1 U396 ( .A(KeyOutxD[6]), .B(K03xD[6]), .Z(n300) );
  XOR2_X1 U397 ( .A(StateInxD[7]), .B(KeyOutxD[7]), .Z(n227) );
  XNOR2_X1 U398 ( .A(RCONxD[7]), .B(n227), .ZN(n228) );
  XOR2_X1 U399 ( .A(KeyOutxD[7]), .B(K03xD[7]), .Z(n229) );
  AOI22_X1 U400 ( .A1(FinishedxS), .A2(KxDI[7]), .B1(n332), .B2(n229), .ZN(
        n230) );
  OAI21_X1 U401 ( .B1(n333), .B2(n228), .A(n230), .ZN(KeyInxD[7]) );
  AOI22_X1 U402 ( .A1(n331), .A2(StateInxD[8]), .B1(n332), .B2(K03xD[8]), .ZN(
        n231) );
  OAI22_X1 U403 ( .A1(n333), .A2(StateInxD[8]), .B1(n334), .B2(K03xD[8]), .ZN(
        n232) );
  AOI22_X1 U404 ( .A1(FinishedxS), .A2(KxDI[8]), .B1(KeyOutxD[8]), .B2(n232), 
        .ZN(n233) );
  OAI21_X1 U405 ( .B1(KeyOutxD[8]), .B2(n231), .A(n233), .ZN(KeyInxD[8]) );
  AOI22_X1 U406 ( .A1(n331), .A2(StateInxD[9]), .B1(n332), .B2(K03xD[9]), .ZN(
        n234) );
  OAI22_X1 U407 ( .A1(n333), .A2(StateInxD[9]), .B1(n334), .B2(K03xD[9]), .ZN(
        n235) );
  AOI22_X1 U408 ( .A1(FinishedxS), .A2(KxDI[9]), .B1(KeyOutxD[9]), .B2(n235), 
        .ZN(n236) );
  OAI21_X1 U409 ( .B1(KeyOutxD[9]), .B2(n234), .A(n236), .ZN(KeyInxD[9]) );
  AOI22_X1 U410 ( .A1(n331), .A2(StateInxD[10]), .B1(n332), .B2(K03xD[10]), 
        .ZN(n237) );
  OAI22_X1 U411 ( .A1(n333), .A2(StateInxD[10]), .B1(n334), .B2(K03xD[10]), 
        .ZN(n238) );
  AOI22_X1 U412 ( .A1(FinishedxS), .A2(KxDI[10]), .B1(KeyOutxD[10]), .B2(n238), 
        .ZN(n239) );
  OAI21_X1 U413 ( .B1(KeyOutxD[10]), .B2(n237), .A(n239), .ZN(KeyInxD[10]) );
  AOI22_X1 U414 ( .A1(n331), .A2(StateInxD[11]), .B1(n332), .B2(K03xD[11]), 
        .ZN(n240) );
  OAI22_X1 U415 ( .A1(n333), .A2(StateInxD[11]), .B1(n334), .B2(K03xD[11]), 
        .ZN(n241) );
  AOI22_X1 U416 ( .A1(FinishedxS), .A2(KxDI[11]), .B1(KeyOutxD[11]), .B2(n241), 
        .ZN(n242) );
  OAI21_X1 U417 ( .B1(KeyOutxD[11]), .B2(n240), .A(n242), .ZN(KeyInxD[11]) );
  AOI22_X1 U418 ( .A1(n331), .A2(StateInxD[12]), .B1(n332), .B2(K03xD[12]), 
        .ZN(n243) );
  OAI22_X1 U419 ( .A1(n333), .A2(StateInxD[12]), .B1(n334), .B2(K03xD[12]), 
        .ZN(n244) );
  AOI22_X1 U420 ( .A1(FinishedxS), .A2(KxDI[12]), .B1(KeyOutxD[12]), .B2(n244), 
        .ZN(n245) );
  OAI21_X1 U421 ( .B1(KeyOutxD[12]), .B2(n243), .A(n245), .ZN(KeyInxD[12]) );
  AOI22_X1 U422 ( .A1(K03xD[13]), .A2(n332), .B1(StateInxD[13]), .B2(n331), 
        .ZN(n246) );
  AOI22_X1 U423 ( .A1(FinishedxS), .A2(KxDI[13]), .B1(KeyOutxD[13]), .B2(n324), 
        .ZN(n247) );
  OAI21_X1 U424 ( .B1(KeyOutxD[13]), .B2(n246), .A(n247), .ZN(KeyInxD[13]) );
  AOI22_X1 U425 ( .A1(StateOutxD[14]), .A2(n336), .B1(PTxDI[14]), .B2(n335), 
        .ZN(n248) );
  AOI22_X1 U426 ( .A1(n114), .A2(KeyToSboxOutxD[14]), .B1(KeyInxD[14]), .B2(
        n330), .ZN(n249) );
  OAI21_X1 U427 ( .B1(KeyInxD[14]), .B2(n248), .A(n249), .ZN(CxDO[14]) );
  AOI22_X1 U428 ( .A1(n331), .A2(StateInxD[15]), .B1(n332), .B2(K03xD[15]), 
        .ZN(n250) );
  OAI22_X1 U429 ( .A1(n333), .A2(StateInxD[15]), .B1(n334), .B2(K03xD[15]), 
        .ZN(n251) );
  AOI22_X1 U430 ( .A1(FinishedxS), .A2(KxDI[15]), .B1(KeyOutxD[15]), .B2(n251), 
        .ZN(n252) );
  OAI21_X1 U431 ( .B1(KeyOutxD[15]), .B2(n250), .A(n252), .ZN(KeyInxD[15]) );
  AOI22_X1 U432 ( .A1(n331), .A2(StateInxD[14]), .B1(K03xD[14]), .B2(n332), 
        .ZN(n253) );
  OAI21_X1 U433 ( .B1(KeyOutxD[14]), .B2(n253), .A(n329), .ZN(KeyInxD[14]) );
  INV_X1 U434 ( .A(ClkxCI), .ZN(n254) );
  NOR2_X4 U435 ( .A1(FinishedxS), .A2(n114), .ZN(n336) );
  INV_X4 U436 ( .A(n260), .ZN(n114) );
  NOR2_X4 U437 ( .A1(FinishedxS), .A2(StateKEYADDITION1o3xS), .ZN(n332) );
  NOR2_X1 U438 ( .A1(n226), .A2(n254), .ZN(ClkKeyRegxC) );
  AOI22_X1 U439 ( .A1(n336), .A2(StateOutxD[0]), .B1(n335), .B2(PTxDI[0]), 
        .ZN(n263) );
  AOI22_X1 U440 ( .A1(n336), .A2(StateOutxD[1]), .B1(n335), .B2(PTxDI[1]), 
        .ZN(n270) );
  AOI22_X1 U441 ( .A1(KeyToSboxOutxD[1]), .A2(n114), .B1(n268), .B2(KeyInxD[1]), .ZN(n269) );
  AOI22_X1 U442 ( .A1(n336), .A2(StateOutxD[2]), .B1(n335), .B2(PTxDI[2]), 
        .ZN(n277) );
  AOI22_X1 U443 ( .A1(n336), .A2(StateOutxD[4]), .B1(n335), .B2(PTxDI[4]), 
        .ZN(n291) );
  AOI22_X1 U444 ( .A1(n336), .A2(StateOutxD[6]), .B1(n335), .B2(PTxDI[6]), 
        .ZN(n305) );
  AOI22_X1 U445 ( .A1(n336), .A2(StateOutxD[7]), .B1(n335), .B2(PTxDI[7]), 
        .ZN(n308) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U31 ( .A1(aes_ctrl_lsfr_23_cycles_1_n23), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n17), .ZN(nextRCONxS) );
  OAI22_X1 aes_ctrl_lsfr_23_cycles_1_U30 ( .A1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n23), .B1(aes_ctrl_lsfr_23_cycles_1_n3), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n24), .ZN(aes_ctrl_lsfr_23_cycles_1_n39)
         );
  AOI221_X1 aes_ctrl_lsfr_23_cycles_1_U29 ( .B1(StartxSI), .B2(
        aes_ctrl_lsfr_23_cycles_1_n22), .C1(aes_ctrl_lsfr_23_cycles_1_n21), 
        .C2(aes_ctrl_lsfr_23_cycles_1_n22), .A(aes_ctrl_lsfr_23_cycles_1_n8), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n3) );
  XNOR2_X1 aes_ctrl_lsfr_23_cycles_1_U28 ( .A(aes_ctrl_lsfr_23_cycles_1_n1), 
        .B(aes_ctrl_lsfr_23_cycles_1_n5), .ZN(aes_ctrl_lsfr_23_cycles_1_n36)
         );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U27 ( .A1(aes_ctrl_lsfr_23_cycles_1_n22), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n19), .ZN(aes_ctrl_lsfr_23_cycles_1_n1)
         );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U26 ( .A1(aes_ctrl_lsfr_23_cycles_1_n18), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n14), .ZN(aes_ctrl_lsfr_23_cycles_1_N16)
         );
  AOI211_X1 aes_ctrl_lsfr_23_cycles_1_U25 ( .C1(aes_ctrl_lsfr_23_cycles_1_n4), 
        .C2(aes_ctrl_lsfr_23_cycles_1_n11), .A(aes_ctrl_lsfr_23_cycles_1_n13), 
        .B(aes_ctrl_lsfr_23_cycles_1_n7), .ZN(aes_ctrl_lsfr_23_cycles_1_N66)
         );
  OAI22_X1 aes_ctrl_lsfr_23_cycles_1_U24 ( .A1(aes_ctrl_lsfr_23_cycles_1_n7), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n15), .B1(aes_ctrl_lsfr_23_cycles_1_n17), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n14), .ZN(aes_ctrl_lsfr_23_cycles_1_N83)
         );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U23 ( .A1(aes_ctrl_lsfr_23_cycles_1_n6), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n17), .ZN(disableKeyRegsxS) );
  AOI22_X1 aes_ctrl_lsfr_23_cycles_1_U22 ( .A1(aes_ctrl_lsfr_23_cycles_1_n20), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n4), .B1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n23), .ZN(aes_ctrl_lsfr_23_cycles_1_n37)
         );
  OAI221_X1 aes_ctrl_lsfr_23_cycles_1_U21 ( .B1(aes_ctrl_lsfr_23_cycles_1_n20), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n4), .C1(aes_ctrl_lsfr_23_cycles_1_n23), 
        .C2(aes_ctrl_lsfr_23_cycles_1_n18), .A(aes_ctrl_lsfr_23_cycles_1_n22), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n35) );
  XNOR2_X1 aes_ctrl_lsfr_23_cycles_1_U20 ( .A(aes_ctrl_lsfr_23_cycles_1_n24), 
        .B(aes_ctrl_lsfr_23_cycles_1_n9), .ZN(aes_ctrl_lsfr_23_cycles_1_n38)
         );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U19 ( .A1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n4), .ZN(aes_ctrl_lsfr_23_cycles_1_n18)
         );
  NAND3_X1 aes_ctrl_lsfr_23_cycles_1_U18 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n9), .A3(aes_ctrl_lsfr_23_cycles_1_n6), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n14) );
  OAI21_X1 aes_ctrl_lsfr_23_cycles_1_U17 ( .B1(aes_ctrl_lsfr_23_cycles_1_n10), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n8), .A(aes_ctrl_lsfr_23_cycles_1_n5), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n11) );
  NOR2_X2 aes_ctrl_lsfr_23_cycles_1_U16 ( .A1(aes_ctrl_lsfr_23_cycles_1_n4), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n11), .ZN(aes_ctrl_lsfr_23_cycles_1_n13)
         );
  INV_X1 aes_ctrl_lsfr_23_cycles_1_U15 ( .A(aes_ctrl_lsfr_23_cycles_1_n13), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n15) );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U14 ( .A1(aes_ctrl_lsfr_23_cycles_1_n4), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n7), .ZN(aes_ctrl_lsfr_23_cycles_1_n17)
         );
  AND2_X1 aes_ctrl_lsfr_23_cycles_1_U13 ( .A1(aes_ctrl_lsfr_23_cycles_1_n8), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n22), .ZN(aes_ctrl_lsfr_23_cycles_1_n24)
         );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U12 ( .A1(aes_ctrl_lsfr_23_cycles_1_n19), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n5), .ZN(aes_ctrl_lsfr_23_cycles_1_n23)
         );
  OR2_X1 aes_ctrl_lsfr_23_cycles_1_U11 ( .A1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n4), .ZN(aes_ctrl_lsfr_23_cycles_1_n22)
         );
  OR3_X1 aes_ctrl_lsfr_23_cycles_1_U10 ( .A1(aes_ctrl_lsfr_23_cycles_1_n18), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n10), .A3(aes_ctrl_lsfr_23_cycles_1_n5), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n21) );
  INV_X1 aes_ctrl_lsfr_23_cycles_1_U9 ( .A(aes_ctrl_lsfr_23_cycles_1_n23), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n20) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U8 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n9), .ZN(aes_ctrl_lsfr_23_cycles_1_n19)
         );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U7 ( .A1(aes_ctrl_lsfr_23_cycles_1_n17), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n16), .ZN(StateKEYSCHEDULExS) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U6 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n21), .ZN(showRCONxS) );
  NOR4_X1 aes_ctrl_lsfr_23_cycles_1_U5 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(LastRoundxS), .A3(aes_ctrl_lsfr_23_cycles_1_n7), .A4(
        aes_ctrl_lsfr_23_cycles_1_n10), .ZN(doMixColumnsxS) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U4 ( .A1(aes_ctrl_lsfr_23_cycles_1_n18), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n16), .ZN(StateKEYADDITION1o3xS) );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U3 ( .A1(aes_ctrl_lsfr_23_cycles_1_n11), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n14), .ZN(aes_ctrl_lsfr_23_cycles_1_n16)
         );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_2_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n36), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n5), .QN(aes_ctrl_lsfr_23_cycles_1_n6) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_1_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n38), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n10), .QN(aes_ctrl_lsfr_23_cycles_1_n9) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_3_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n35), .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(
        aes_ctrl_lsfr_23_cycles_1_n4) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_4_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n37), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n7), .QN(aes_ctrl_lsfr_23_cycles_1_n2) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_0_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n39), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n8), .QN(aes_ctrl_lsfr_23_cycles_1_n12) );
  INV_X1 rcon_1_U37 ( .A(nextRCONxS), .ZN(rcon_1_n39) );
  AOI211_X1 rcon_1_U36 ( .C1(rcon_1_n9), .C2(rcon_1_n28), .A(rcon_1_n43), .B(
        rcon_1_n29), .ZN(rcon_1_n22) );
  OAI22_X1 rcon_1_U35 ( .A1(rcon_1_n38), .A2(rcon_1_n4), .B1(rcon_1_n9), .B2(
        rcon_1_n42), .ZN(rcon_1_n29) );
  INV_X1 rcon_1_U34 ( .A(rcon_1_n44), .ZN(rcon_1_n28) );
  INV_X1 rcon_1_U32 ( .A(rcon_1_n38), .ZN(rcon_1_n16) );
  INV_X1 rcon_1_U31 ( .A(rcon_1_n35), .ZN(rcon_1_n15) );
  OAI211_X1 rcon_1_U30 ( .C1(rcon_1_n38), .C2(rcon_1_n17), .A(rcon_1_n44), .B(
        rcon_1_n14), .ZN(rcon_1_n25) );
  INV_X1 rcon_1_U29 ( .A(rcon_1_n43), .ZN(rcon_1_n14) );
  AOI211_X1 rcon_1_U28 ( .C1(rcon_1_n39), .C2(rcon_1_n34), .A(rcon_1_n43), .B(
        rcon_1_n13), .ZN(rcon_1_n24) );
  AOI22_X1 rcon_1_U27 ( .A1(rcon_1_n37), .A2(rcon_1_n44), .B1(rcon_1_n42), 
        .B2(rcon_1_n17), .ZN(rcon_1_n13) );
  OAI21_X1 rcon_1_U26 ( .B1(rcon_1_n38), .B2(rcon_1_n33), .A(rcon_1_n12), .ZN(
        rcon_1_n21) );
  OAI211_X1 rcon_1_U25 ( .C1(rcon_1_n35), .C2(rcon_1_n4), .A(rcon_1_n38), .B(
        rcon_1_n11), .ZN(rcon_1_n12) );
  OAI21_X1 rcon_1_U24 ( .B1(rcon_1_n35), .B2(rcon_1_n36), .A(rcon_1_n4), .ZN(
        rcon_1_n11) );
  NOR2_X1 rcon_1_U23 ( .A1(rcon_1_n32), .A2(rcon_1_n40), .ZN(RCONxD[7]) );
  OAI22_X1 rcon_1_U22 ( .A1(rcon_1_n26), .A2(rcon_1_n38), .B1(rcon_1_n30), 
        .B2(rcon_1_n41), .ZN(rcon_1_n19) );
  OAI22_X1 rcon_1_U21 ( .A1(rcon_1_n38), .A2(rcon_1_n30), .B1(rcon_1_n33), 
        .B2(rcon_1_n41), .ZN(rcon_1_n20) );
  OAI22_X1 rcon_1_U20 ( .A1(rcon_1_n38), .A2(rcon_1_n31), .B1(rcon_1_n34), 
        .B2(rcon_1_n41), .ZN(rcon_1_n23) );
  NOR2_X1 rcon_1_U19 ( .A1(rcon_1_n26), .A2(rcon_1_n40), .ZN(RCONxD[6]) );
  NOR2_X1 rcon_1_U18 ( .A1(rcon_1_n30), .A2(rcon_1_n40), .ZN(RCONxD[5]) );
  NOR2_X1 rcon_1_U17 ( .A1(rcon_1_n33), .A2(rcon_1_n40), .ZN(RCONxD[4]) );
  AND2_X1 rcon_1_U16 ( .A1(rcon_1_n4), .A2(showRCONxS), .ZN(RCONxD[3]) );
  NOR2_X1 rcon_1_U15 ( .A1(rcon_1_n31), .A2(rcon_1_n40), .ZN(RCONxD[2]) );
  NOR2_X1 rcon_1_U14 ( .A1(rcon_1_n34), .A2(rcon_1_n40), .ZN(RCONxD[1]) );
  NOR2_X1 rcon_1_U13 ( .A1(rcon_1_n17), .A2(rcon_1_n40), .ZN(RCONxD[0]) );
  NAND2_X1 rcon_1_U12 ( .A1(rcon_1_n38), .A2(rcon_1_n45), .ZN(rcon_1_n41) );
  INV_X1 rcon_1_U11 ( .A(rcon_1_n39), .ZN(rcon_1_n38) );
  NOR2_X1 rcon_1_U10 ( .A1(rcon_1_n45), .A2(rcon_1_n39), .ZN(rcon_1_n43) );
  NAND2_X1 rcon_1_U9 ( .A1(rcon_1_n38), .A2(rcon_1_n35), .ZN(rcon_1_n44) );
  NAND2_X1 rcon_1_U8 ( .A1(rcon_1_n38), .A2(rcon_1_n32), .ZN(rcon_1_n42) );
  INV_X2 rcon_1_U7 ( .A(rcon_1_n45), .ZN(FinishedxS) );
  INV_X1 rcon_1_U6 ( .A(showRCONxS), .ZN(rcon_1_n40) );
  NOR2_X1 rcon_1_U5 ( .A1(rcon_1_n30), .A2(rcon_1_n31), .ZN(LastRoundxS) );
  NAND2_X1 rcon_1_U4 ( .A1(rcon_1_n36), .A2(rcon_1_n4), .ZN(rcon_1_n45) );
  OAI33_X1 rcon_1_U3 ( .A1(1'b0), .A2(rcon_1_n38), .A3(rcon_1_n15), .B1(
        rcon_1_n16), .B2(rcon_1_n26), .B3(rcon_1_n4), .ZN(rcon_1_n18) );
  DFFR_X1 rcon_1_RCONxDP_reg_4_ ( .D(rcon_1_n21), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(rcon_1_n33) );
  DFFR_X1 rcon_1_RCONxDP_reg_1_ ( .D(rcon_1_n24), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(rcon_1_n34) );
  DFFR_X1 rcon_1_RCONxDP_reg_0_ ( .D(rcon_1_n25), .CK(ClkxCI), .RN(RstxBI), 
        .Q(rcon_1_n37), .QN(rcon_1_n17) );
  DFFR_X1 rcon_1_RCONxDP_reg_7_ ( .D(rcon_1_n18), .CK(ClkxCI), .RN(RstxBI), 
        .Q(rcon_1_n35), .QN(rcon_1_n32) );
  DFFS_X1 rcon_1_RCONxDP_reg_3_ ( .D(rcon_1_n22), .CK(ClkxCI), .SN(RstxBI), 
        .Q(rcon_1_n4), .QN() );
  DFFS_X1 rcon_1_RCONxDP_reg_2_ ( .D(rcon_1_n23), .CK(ClkxCI), .SN(RstxBI), 
        .Q(rcon_1_n9), .QN(rcon_1_n31) );
  DFFS_X1 rcon_1_RCONxDP_reg_5_ ( .D(rcon_1_n20), .CK(ClkxCI), .SN(RstxBI), 
        .Q(), .QN(rcon_1_n30) );
  DFFS_X1 rcon_1_RCONxDP_reg_6_ ( .D(rcon_1_n19), .CK(ClkxCI), .SN(RstxBI), 
        .Q(rcon_1_n36), .QN(rcon_1_n26) );
  DFF_X1 SBOX_regOut2_reg_0__0_ ( .D(SBOX_regOut1[0]), .CK(ClkxCI), .Q(), .QN(
        StateInxD[0]) );
  DFF_X1 SBOX_regOut1_reg_0__0_ ( .D(SBOX_stage6Out[0]), .CK(ClkxCI), .Q(
        SBOX_regOut1[0]), .QN() );
  DFF_X1 SBOX_regOut2_reg_0__1_ ( .D(SBOX_regOut1[1]), .CK(ClkxCI), .Q(), .QN(
        StateInxD[1]) );
  DFF_X1 SBOX_regOut1_reg_0__1_ ( .D(SBOX_stage6Out[1]), .CK(ClkxCI), .Q(
        SBOX_regOut1[1]), .QN() );
  DFF_X1 SBOX_regOut2_reg_0__2_ ( .D(SBOX_regOut1[2]), .CK(ClkxCI), .Q(
        StateInxD[2]), .QN() );
  DFF_X1 SBOX_regOut1_reg_0__2_ ( .D(SBOX_stage6Out[2]), .CK(ClkxCI), .Q(
        SBOX_regOut1[2]), .QN() );
  DFF_X1 SBOX_regOut2_reg_0__3_ ( .D(SBOX_regOut1[3]), .CK(ClkxCI), .Q(
        StateInxD[3]), .QN() );
  DFF_X1 SBOX_regOut1_reg_0__3_ ( .D(SBOX_stage6Out[3]), .CK(ClkxCI), .Q(
        SBOX_regOut1[3]), .QN() );
  DFF_X1 SBOX_regOut2_reg_0__4_ ( .D(SBOX_regOut1[4]), .CK(ClkxCI), .Q(
        StateInxD[4]), .QN() );
  DFF_X1 SBOX_regOut1_reg_0__4_ ( .D(SBOX_stage6Out[4]), .CK(ClkxCI), .Q(
        SBOX_regOut1[4]), .QN() );
  DFF_X1 SBOX_regOut2_reg_0__5_ ( .D(SBOX_regOut1[5]), .CK(ClkxCI), .Q(), .QN(
        StateInxD[5]) );
  DFF_X1 SBOX_regOut1_reg_0__5_ ( .D(SBOX_stage6Out[5]), .CK(ClkxCI), .Q(
        SBOX_regOut1[5]), .QN() );
  DFF_X1 SBOX_regOut2_reg_0__6_ ( .D(SBOX_regOut1[6]), .CK(ClkxCI), .Q(), .QN(
        StateInxD[6]) );
  DFF_X1 SBOX_regOut1_reg_0__6_ ( .D(SBOX_stage6Out[6]), .CK(ClkxCI), .Q(
        SBOX_regOut1[6]), .QN() );
  DFF_X1 SBOX_regOut2_reg_0__7_ ( .D(SBOX_regOut1[7]), .CK(ClkxCI), .Q(
        StateInxD[7]), .QN() );
  DFF_X1 SBOX_regOut1_reg_0__7_ ( .D(SBOX_stage6Out[7]), .CK(ClkxCI), .Q(
        SBOX_regOut1[7]), .QN() );
  DFF_X1 SBOX_regOut2_reg_1__0_ ( .D(SBOX_regOut1[8]), .CK(ClkxCI), .Q(
        StateInxD[8]), .QN() );
  DFF_X1 SBOX_regOut1_reg_1__0_ ( .D(SBOX_stage6Out[8]), .CK(ClkxCI), .Q(
        SBOX_regOut1[8]), .QN() );
  DFF_X1 SBOX_regOut2_reg_1__1_ ( .D(SBOX_regOut1[9]), .CK(ClkxCI), .Q(
        StateInxD[9]), .QN() );
  DFF_X1 SBOX_regOut1_reg_1__1_ ( .D(SBOX_stage6Out[9]), .CK(ClkxCI), .Q(
        SBOX_regOut1[9]), .QN() );
  DFF_X1 SBOX_regOut2_reg_1__2_ ( .D(SBOX_regOut1[10]), .CK(ClkxCI), .Q(
        StateInxD[10]), .QN() );
  DFF_X1 SBOX_regOut1_reg_1__2_ ( .D(SBOX_stage6Out[10]), .CK(ClkxCI), .Q(
        SBOX_regOut1[10]), .QN() );
  DFF_X1 SBOX_regOut2_reg_1__3_ ( .D(SBOX_regOut1[11]), .CK(ClkxCI), .Q(
        StateInxD[11]), .QN() );
  DFF_X1 SBOX_regOut1_reg_1__3_ ( .D(SBOX_stage6Out[11]), .CK(ClkxCI), .Q(
        SBOX_regOut1[11]), .QN() );
  DFF_X1 SBOX_regOut2_reg_1__4_ ( .D(SBOX_regOut1[12]), .CK(ClkxCI), .Q(
        StateInxD[12]), .QN() );
  DFF_X1 SBOX_regOut1_reg_1__4_ ( .D(SBOX_stage6Out[12]), .CK(ClkxCI), .Q(
        SBOX_regOut1[12]), .QN() );
  DFF_X1 SBOX_regOut2_reg_1__5_ ( .D(SBOX_regOut1[13]), .CK(ClkxCI), .Q(
        StateInxD[13]), .QN() );
  DFF_X1 SBOX_regOut1_reg_1__5_ ( .D(SBOX_stage6Out[13]), .CK(ClkxCI), .Q(
        SBOX_regOut1[13]), .QN() );
  DFF_X1 SBOX_regOut2_reg_1__6_ ( .D(SBOX_regOut1[14]), .CK(ClkxCI), .Q(
        StateInxD[14]), .QN() );
  DFF_X1 SBOX_regOut1_reg_1__6_ ( .D(SBOX_stage6Out[14]), .CK(ClkxCI), .Q(
        SBOX_regOut1[14]), .QN() );
  DFF_X1 SBOX_regOut2_reg_1__7_ ( .D(SBOX_regOut1[15]), .CK(ClkxCI), .Q(
        StateInxD[15]), .QN() );
  DFF_X1 SBOX_regOut1_reg_1__7_ ( .D(SBOX_stage6Out[15]), .CK(ClkxCI), .Q(
        SBOX_regOut1[15]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_0__0_ ( .D(SBOX_s1_linMapOut_0__0_), .CK(ClkxCI), .Q(SBOX_stage1Out[0]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_0__1_ ( .D(SBOX_s1_linMapOut_0__1_), .CK(ClkxCI), .Q(SBOX_stage1Out[1]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_0__2_ ( .D(CxDO[0]), .CK(ClkxCI), .Q(
        SBOX_stage1Out[2]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_0__3_ ( .D(SBOX_s1_linMapOut_0__3_), .CK(ClkxCI), .Q(SBOX_stage1Out[3]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_0__4_ ( .D(SBOX_s1_linMapOut_0__4_), .CK(ClkxCI), .Q(SBOX_stage1Out[4]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_0__5_ ( .D(SBOX_s1_linMapOut_0__5_), .CK(ClkxCI), .Q(SBOX_stage1Out[5]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_0__6_ ( .D(SBOX_s1_linMapOut_0__6_), .CK(ClkxCI), .Q(SBOX_stage1Out[6]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_0__7_ ( .D(SBOX_s1_linMapOut_0__7_), .CK(ClkxCI), .Q(SBOX_stage1Out[7]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_1__0_ ( .D(SBOX_s1_linMapOut_1__0_), .CK(ClkxCI), .Q(SBOX_stage1Out[8]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_1__1_ ( .D(SBOX_s1_linMapOut_1__1_), .CK(ClkxCI), .Q(SBOX_stage1Out[9]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_1__2_ ( .D(CxDO[8]), .CK(ClkxCI), .Q(
        SBOX_stage1Out[10]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_1__3_ ( .D(SBOX_s1_linMapOut_1__3_), .CK(ClkxCI), .Q(SBOX_stage1Out[11]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_1__4_ ( .D(SBOX_s1_linMapOut_1__4_), .CK(ClkxCI), .Q(SBOX_stage1Out[12]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_1__5_ ( .D(SBOX_s1_linMapOut_1__5_), .CK(ClkxCI), .Q(SBOX_stage1Out[13]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_1__6_ ( .D(SBOX_s1_linMapOut_1__6_), .CK(ClkxCI), .Q(SBOX_stage1Out[14]), .QN() );
  DFF_X1 SBOX_s1_stage1Out_reg_1__7_ ( .D(SBOX_s1_linMapOut_1__7_), .CK(ClkxCI), .Q(SBOX_stage1Out[15]), .QN() );
  XNOR2_X1 SBOX_s1_input_mapping_1_U14 ( .A(SBOX_s1_input_mapping_1_n20), .B(
        SBOX_s1_input_mapping_1_n19), .ZN(SBOX_s1_linMapOut_1__3_) );
  XNOR2_X1 SBOX_s1_input_mapping_1_U13 ( .A(SBOX_s1_input_mapping_1_n18), .B(
        CxDO[11]), .ZN(SBOX_s1_input_mapping_1_n19) );
  XNOR2_X1 SBOX_s1_input_mapping_1_U12 ( .A(CxDO[15]), .B(CxDO[12]), .ZN(
        SBOX_s1_input_mapping_1_n18) );
  XNOR2_X1 SBOX_s1_input_mapping_1_U11 ( .A(SBOX_s1_input_mapping_1_n17), .B(
        CxDO[11]), .ZN(SBOX_s1_linMapOut_1__0_) );
  XNOR2_X1 SBOX_s1_input_mapping_1_U10 ( .A(CxDO[14]), .B(
        SBOX_s1_input_mapping_1_n23), .ZN(SBOX_s1_input_mapping_1_n17) );
  XNOR2_X1 SBOX_s1_input_mapping_1_U9 ( .A(SBOX_s1_input_mapping_1_n23), .B(
        SBOX_s1_input_mapping_1_n22), .ZN(SBOX_s1_linMapOut_1__7_) );
  XOR2_X1 SBOX_s1_input_mapping_1_U8 ( .A(CxDO[12]), .B(
        SBOX_s1_linMapOut_1__1_), .Z(SBOX_s1_linMapOut_1__6_) );
  XNOR2_X1 SBOX_s1_input_mapping_1_U7 ( .A(SBOX_s1_input_mapping_1_n21), .B(
        SBOX_s1_input_mapping_1_n20), .ZN(SBOX_s1_linMapOut_1__5_) );
  XNOR2_X1 SBOX_s1_input_mapping_1_U6 ( .A(CxDO[8]), .B(
        SBOX_s1_input_mapping_1_n22), .ZN(SBOX_s1_linMapOut_1__4_) );
  XOR2_X1 SBOX_s1_input_mapping_1_U5 ( .A(CxDO[8]), .B(
        SBOX_s1_input_mapping_1_n21), .Z(SBOX_s1_linMapOut_1__1_) );
  XNOR2_X1 SBOX_s1_input_mapping_1_U4 ( .A(CxDO[10]), .B(
        SBOX_s1_input_mapping_1_n20), .ZN(SBOX_s1_input_mapping_1_n23) );
  XNOR2_X1 SBOX_s1_input_mapping_1_U3 ( .A(CxDO[15]), .B(
        SBOX_s1_input_mapping_1_n21), .ZN(SBOX_s1_input_mapping_1_n22) );
  XNOR2_X1 SBOX_s1_input_mapping_1_U2 ( .A(CxDO[8]), .B(CxDO[9]), .ZN(
        SBOX_s1_input_mapping_1_n20) );
  XOR2_X1 SBOX_s1_input_mapping_1_U1 ( .A(CxDO[14]), .B(CxDO[13]), .Z(
        SBOX_s1_input_mapping_1_n21) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U14 ( .A(SBOX_s1_input_mapping_0_n20), .B(
        SBOX_s1_input_mapping_0_n19), .ZN(SBOX_s1_linMapOut_0__3_) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U13 ( .A(SBOX_s1_input_mapping_0_n18), .B(
        CxDO[3]), .ZN(SBOX_s1_input_mapping_0_n19) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U12 ( .A(CxDO[7]), .B(CxDO[4]), .ZN(
        SBOX_s1_input_mapping_0_n18) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U11 ( .A(SBOX_s1_input_mapping_0_n17), .B(
        CxDO[3]), .ZN(SBOX_s1_linMapOut_0__0_) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U10 ( .A(CxDO[6]), .B(
        SBOX_s1_input_mapping_0_n23), .ZN(SBOX_s1_input_mapping_0_n17) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U9 ( .A(SBOX_s1_input_mapping_0_n23), .B(
        SBOX_s1_input_mapping_0_n22), .ZN(SBOX_s1_linMapOut_0__7_) );
  XOR2_X1 SBOX_s1_input_mapping_0_U8 ( .A(CxDO[4]), .B(SBOX_s1_linMapOut_0__1_), .Z(SBOX_s1_linMapOut_0__6_) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U7 ( .A(SBOX_s1_input_mapping_0_n21), .B(
        SBOX_s1_input_mapping_0_n20), .ZN(SBOX_s1_linMapOut_0__5_) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U6 ( .A(CxDO[0]), .B(
        SBOX_s1_input_mapping_0_n22), .ZN(SBOX_s1_linMapOut_0__4_) );
  XOR2_X1 SBOX_s1_input_mapping_0_U5 ( .A(CxDO[0]), .B(
        SBOX_s1_input_mapping_0_n21), .Z(SBOX_s1_linMapOut_0__1_) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U4 ( .A(CxDO[2]), .B(
        SBOX_s1_input_mapping_0_n20), .ZN(SBOX_s1_input_mapping_0_n23) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U3 ( .A(CxDO[7]), .B(
        SBOX_s1_input_mapping_0_n21), .ZN(SBOX_s1_input_mapping_0_n22) );
  XOR2_X1 SBOX_s1_input_mapping_0_U2 ( .A(CxDO[6]), .B(CxDO[5]), .Z(
        SBOX_s1_input_mapping_0_n21) );
  XNOR2_X1 SBOX_s1_input_mapping_0_U1 ( .A(CxDO[0]), .B(CxDO[1]), .ZN(
        SBOX_s1_input_mapping_0_n20) );
  XOR2_X1 SBOX_s2_U42 ( .A(SBOX_s2_sqsc_out[5]), .B(SBOX_s2_n16), .Z(
        SBOX_s2_refreshed[13]) );
  XNOR2_X1 SBOX_s2_U41 ( .A(SBOX_s2_n14), .B(SBOX_s2_n15), .ZN(SBOX_s2_n16) );
  XNOR2_X1 SBOX_s2_U40 ( .A(SBOX_s2_gf2_mul_out_1__1__1_), .B(randomS2[9]), 
        .ZN(SBOX_s2_n15) );
  XOR2_X1 SBOX_s2_U39 ( .A(randomS2[1]), .B(randomS2[5]), .Z(SBOX_s2_n14) );
  XNOR2_X1 SBOX_s2_U38 ( .A(SBOX_s2_n13), .B(SBOX_s2_sqsc_out[1]), .ZN(
        SBOX_s2_refreshed[1]) );
  XNOR2_X1 SBOX_s2_U37 ( .A(randomS2[1]), .B(SBOX_s2_gf2_mul_out_0__0__1_), 
        .ZN(SBOX_s2_n13) );
  XOR2_X1 SBOX_s2_U36 ( .A(SBOX_stage1Out[11]), .B(SBOX_stage1Out[15]), .Z(
        SBOX_s2_sqsc_in[5]) );
  XOR2_X1 SBOX_s2_U35 ( .A(SBOX_s2_sqsc_out[6]), .B(SBOX_s2_n12), .Z(
        SBOX_s2_refreshed[14]) );
  XNOR2_X1 SBOX_s2_U34 ( .A(SBOX_s2_n10), .B(SBOX_s2_n11), .ZN(SBOX_s2_n12) );
  XNOR2_X1 SBOX_s2_U33 ( .A(SBOX_s2_gf2_mul_out_1__1__2_), .B(randomS2[10]), 
        .ZN(SBOX_s2_n11) );
  XOR2_X1 SBOX_s2_U32 ( .A(randomS2[2]), .B(randomS2[6]), .Z(SBOX_s2_n10) );
  XOR2_X1 SBOX_s2_U31 ( .A(SBOX_stage1Out[3]), .B(SBOX_stage1Out[7]), .Z(
        SBOX_s2_sqsc_in[2]) );
  XNOR2_X1 SBOX_s2_U30 ( .A(SBOX_s2_n9), .B(SBOX_s2_sqsc_out[2]), .ZN(
        SBOX_s2_refreshed[2]) );
  XNOR2_X1 SBOX_s2_U29 ( .A(randomS2[2]), .B(SBOX_s2_gf2_mul_out_0__0__2_), 
        .ZN(SBOX_s2_n9) );
  XOR2_X1 SBOX_s2_U28 ( .A(SBOX_stage1Out[10]), .B(SBOX_stage1Out[14]), .Z(
        SBOX_s2_sqsc_in[4]) );
  XOR2_X1 SBOX_s2_U27 ( .A(SBOX_s2_sqsc_out[7]), .B(SBOX_s2_n8), .Z(
        SBOX_s2_refreshed[15]) );
  XNOR2_X1 SBOX_s2_U26 ( .A(SBOX_s2_n6), .B(SBOX_s2_n7), .ZN(SBOX_s2_n8) );
  XNOR2_X1 SBOX_s2_U25 ( .A(SBOX_s2_gf2_mul_out_1__1__3_), .B(randomS2[11]), 
        .ZN(SBOX_s2_n7) );
  XOR2_X1 SBOX_s2_U24 ( .A(randomS2[3]), .B(randomS2[7]), .Z(SBOX_s2_n6) );
  XOR2_X1 SBOX_s2_U23 ( .A(SBOX_stage1Out[2]), .B(SBOX_stage1Out[6]), .Z(
        SBOX_s2_sqsc_in[1]) );
  XNOR2_X1 SBOX_s2_U22 ( .A(SBOX_s2_n5), .B(SBOX_s2_sqsc_out[3]), .ZN(
        SBOX_s2_refreshed[3]) );
  XNOR2_X1 SBOX_s2_U21 ( .A(randomS2[3]), .B(SBOX_s2_gf2_mul_out_0__0__3_), 
        .ZN(SBOX_s2_n5) );
  XOR2_X1 SBOX_s2_U20 ( .A(SBOX_s2_sqsc_out[4]), .B(SBOX_s2_n4), .Z(
        SBOX_s2_refreshed[12]) );
  XNOR2_X1 SBOX_s2_U19 ( .A(SBOX_s2_n2), .B(SBOX_s2_n3), .ZN(SBOX_s2_n4) );
  XNOR2_X1 SBOX_s2_U18 ( .A(SBOX_s2_gf2_mul_out_1__1__0_), .B(randomS2[8]), 
        .ZN(SBOX_s2_n3) );
  XOR2_X1 SBOX_s2_U17 ( .A(randomS2[0]), .B(randomS2[4]), .Z(SBOX_s2_n2) );
  XOR2_X1 SBOX_s2_U16 ( .A(randomS2[11]), .B(SBOX_s2_xorResult[7]), .Z(
        SBOX_s2_refreshed[11]) );
  XOR2_X1 SBOX_s2_U15 ( .A(randomS2[7]), .B(SBOX_s2_xorResult[3]), .Z(
        SBOX_s2_refreshed[7]) );
  XNOR2_X1 SBOX_s2_U14 ( .A(SBOX_s2_n1), .B(SBOX_s2_sqsc_out[0]), .ZN(
        SBOX_s2_refreshed[0]) );
  XNOR2_X1 SBOX_s2_U13 ( .A(randomS2[0]), .B(SBOX_s2_gf2_mul_out_0__0__0_), 
        .ZN(SBOX_s2_n1) );
  XOR2_X1 SBOX_s2_U12 ( .A(randomS2[10]), .B(SBOX_s2_xorResult[6]), .Z(
        SBOX_s2_refreshed[10]) );
  XOR2_X1 SBOX_s2_U11 ( .A(randomS2[9]), .B(SBOX_s2_xorResult[5]), .Z(
        SBOX_s2_refreshed[9]) );
  XOR2_X1 SBOX_s2_U10 ( .A(randomS2[6]), .B(SBOX_s2_xorResult[2]), .Z(
        SBOX_s2_refreshed[6]) );
  XOR2_X1 SBOX_s2_U9 ( .A(randomS2[5]), .B(SBOX_s2_xorResult[1]), .Z(
        SBOX_s2_refreshed[5]) );
  XOR2_X1 SBOX_s2_U8 ( .A(randomS2[8]), .B(SBOX_s2_xorResult[4]), .Z(
        SBOX_s2_refreshed[8]) );
  XOR2_X1 SBOX_s2_U7 ( .A(randomS2[4]), .B(SBOX_s2_xorResult[0]), .Z(
        SBOX_s2_refreshed[4]) );
  XOR2_X1 SBOX_s2_U6 ( .A(SBOX_stage1Out[8]), .B(SBOX_stage1Out[12]), .Z(
        SBOX_s2_sqsc_out[4]) );
  XOR2_X1 SBOX_s2_U5 ( .A(SBOX_stage1Out[9]), .B(SBOX_stage1Out[13]), .Z(
        SBOX_s2_sqsc_in[3]) );
  XOR2_X1 SBOX_s2_U4 ( .A(SBOX_stage1Out[0]), .B(SBOX_stage1Out[4]), .Z(
        SBOX_s2_sqsc_out[0]) );
  XOR2_X1 SBOX_s2_U3 ( .A(SBOX_stage1Out[1]), .B(SBOX_stage1Out[5]), .Z(
        SBOX_s2_sqsc_in[0]) );
  DFF_X1 SBOX_s2_regOut_reg_0__0__0_ ( .D(SBOX_stage1Out[0]), .CK(ClkxCI), .Q(
        SBOX_stage2Out[0]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__0__1_ ( .D(SBOX_stage1Out[1]), .CK(ClkxCI), .Q(
        SBOX_stage2Out[1]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__0__2_ ( .D(SBOX_stage1Out[2]), .CK(ClkxCI), .Q(
        SBOX_stage2Out[2]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__0__3_ ( .D(SBOX_stage1Out[3]), .CK(ClkxCI), .Q(
        SBOX_stage2Out[3]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__1__0_ ( .D(SBOX_s2_refreshed[0]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_0__1__0_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__1__1_ ( .D(SBOX_s2_refreshed[1]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_0__1__1_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__1__2_ ( .D(SBOX_s2_refreshed[2]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_0__1__2_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__1__3_ ( .D(SBOX_s2_refreshed[3]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_0__1__3_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__2__0_ ( .D(SBOX_s2_refreshed[4]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_0__2__0_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__2__1_ ( .D(SBOX_s2_refreshed[5]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_0__2__1_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__2__2_ ( .D(SBOX_s2_refreshed[6]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_0__2__2_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__2__3_ ( .D(SBOX_s2_refreshed[7]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_0__2__3_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__3__0_ ( .D(SBOX_stage1Out[4]), .CK(ClkxCI), .Q(
        SBOX_stage2Out[8]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__3__1_ ( .D(SBOX_stage1Out[5]), .CK(ClkxCI), .Q(
        SBOX_stage2Out[9]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__3__2_ ( .D(SBOX_stage1Out[6]), .CK(ClkxCI), .Q(
        SBOX_stage2Out[10]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_0__3__3_ ( .D(SBOX_stage1Out[7]), .CK(ClkxCI), .Q(
        SBOX_stage2Out[11]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__0__0_ ( .D(SBOX_stage1Out[8]), .CK(ClkxCI), .Q(
        SBOX_stage2Out[12]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__0__1_ ( .D(SBOX_stage1Out[9]), .CK(ClkxCI), .Q(
        SBOX_stage2Out[13]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__0__2_ ( .D(SBOX_stage1Out[10]), .CK(ClkxCI), 
        .Q(SBOX_stage2Out[14]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__0__3_ ( .D(SBOX_stage1Out[11]), .CK(ClkxCI), 
        .Q(SBOX_stage2Out[15]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__1__0_ ( .D(SBOX_s2_refreshed[8]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_1__1__0_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__1__1_ ( .D(SBOX_s2_refreshed[9]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_1__1__1_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__1__2_ ( .D(SBOX_s2_refreshed[10]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_1__1__2_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__1__3_ ( .D(SBOX_s2_refreshed[11]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_1__1__3_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__2__0_ ( .D(SBOX_s2_refreshed[12]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_1__2__0_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__2__1_ ( .D(SBOX_s2_refreshed[13]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_1__2__1_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__2__2_ ( .D(SBOX_s2_refreshed[14]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_1__2__2_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__2__3_ ( .D(SBOX_s2_refreshed[15]), .CK(ClkxCI), 
        .Q(SBOX_s2_regOut_1__2__3_), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__3__0_ ( .D(SBOX_stage1Out[12]), .CK(ClkxCI), 
        .Q(SBOX_stage2Out[20]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__3__1_ ( .D(SBOX_stage1Out[13]), .CK(ClkxCI), 
        .Q(SBOX_stage2Out[21]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__3__2_ ( .D(SBOX_stage1Out[14]), .CK(ClkxCI), 
        .Q(SBOX_stage2Out[22]), .QN() );
  DFF_X1 SBOX_s2_regOut_reg_1__3__3_ ( .D(SBOX_stage1Out[15]), .CK(ClkxCI), 
        .Q(SBOX_stage2Out[23]), .QN() );
  XOR2_X1 SBOX_s2_sqsc_1_U3 ( .A(SBOX_s2_sqsc_out[4]), .B(SBOX_s2_sqsc_in[3]), 
        .Z(SBOX_s2_sqsc_out[5]) );
  XOR2_X1 SBOX_s2_sqsc_1_U2 ( .A(SBOX_s2_sqsc_in[3]), .B(SBOX_s2_sqsc_in[5]), 
        .Z(SBOX_s2_sqsc_out[6]) );
  XOR2_X1 SBOX_s2_sqsc_1_U1 ( .A(SBOX_s2_sqsc_out[4]), .B(SBOX_s2_sqsc_in[4]), 
        .Z(SBOX_s2_sqsc_out[7]) );
  XOR2_X1 SBOX_s2_sqsc_0_U3 ( .A(SBOX_s2_sqsc_out[0]), .B(SBOX_s2_sqsc_in[0]), 
        .Z(SBOX_s2_sqsc_out[1]) );
  XOR2_X1 SBOX_s2_sqsc_0_U2 ( .A(SBOX_s2_sqsc_in[0]), .B(SBOX_s2_sqsc_in[2]), 
        .Z(SBOX_s2_sqsc_out[2]) );
  XOR2_X1 SBOX_s2_sqsc_0_U1 ( .A(SBOX_s2_sqsc_out[0]), .B(SBOX_s2_sqsc_in[1]), 
        .Z(SBOX_s2_sqsc_out[3]) );
  XNOR2_X1 SBOX_s2_mul1_1_1_U29 ( .A(SBOX_s2_mul1_1_1_n68), .B(
        SBOX_s2_mul1_1_1_n69), .ZN(SBOX_s2_gf2_mul_out_1__1__1_) );
  XOR2_X1 SBOX_s2_mul1_1_1_U28 ( .A(SBOX_s2_mul1_1_1_n77), .B(
        SBOX_s2_mul1_1_1_n74), .Z(SBOX_s2_mul1_1_1_n69) );
  NAND2_X1 SBOX_s2_mul1_1_1_U27 ( .A1(SBOX_stage1Out[9]), .A2(
        SBOX_stage1Out[13]), .ZN(SBOX_s2_mul1_1_1_n68) );
  XNOR2_X1 SBOX_s2_mul1_1_1_U26 ( .A(SBOX_s2_mul1_1_1_n66), .B(
        SBOX_s2_mul1_1_1_n67), .ZN(SBOX_s2_gf2_mul_out_1__1__2_) );
  XOR2_X1 SBOX_s2_mul1_1_1_U25 ( .A(SBOX_s2_mul1_1_1_n76), .B(
        SBOX_s2_mul1_1_1_n75), .Z(SBOX_s2_mul1_1_1_n67) );
  NAND2_X1 SBOX_s2_mul1_1_1_U24 ( .A1(SBOX_stage1Out[10]), .A2(
        SBOX_stage1Out[14]), .ZN(SBOX_s2_mul1_1_1_n66) );
  XNOR2_X1 SBOX_s2_mul1_1_1_U23 ( .A(SBOX_s2_mul1_1_1_n64), .B(
        SBOX_s2_mul1_1_1_n65), .ZN(SBOX_s2_gf2_mul_out_1__1__3_) );
  XOR2_X1 SBOX_s2_mul1_1_1_U22 ( .A(SBOX_s2_mul1_1_1_n77), .B(
        SBOX_s2_mul1_1_1_n76), .Z(SBOX_s2_mul1_1_1_n65) );
  NAND2_X1 SBOX_s2_mul1_1_1_U21 ( .A1(SBOX_stage1Out[11]), .A2(
        SBOX_stage1Out[15]), .ZN(SBOX_s2_mul1_1_1_n64) );
  XNOR2_X1 SBOX_s2_mul1_1_1_U20 ( .A(SBOX_s2_mul1_1_1_n62), .B(
        SBOX_s2_mul1_1_1_n63), .ZN(SBOX_s2_gf2_mul_out_1__1__0_) );
  XOR2_X1 SBOX_s2_mul1_1_1_U19 ( .A(SBOX_s2_mul1_1_1_n74), .B(
        SBOX_s2_mul1_1_1_n75), .Z(SBOX_s2_mul1_1_1_n63) );
  NAND2_X1 SBOX_s2_mul1_1_1_U18 ( .A1(SBOX_stage1Out[8]), .A2(
        SBOX_stage1Out[12]), .ZN(SBOX_s2_mul1_1_1_n62) );
  AOI221_X1 SBOX_s2_mul1_1_1_U17 ( .B1(SBOX_stage1Out[15]), .B2(
        SBOX_stage1Out[14]), .C1(SBOX_stage1Out[10]), .C2(SBOX_stage1Out[11]), 
        .A(SBOX_s2_mul1_1_1_n61), .ZN(SBOX_s2_mul1_1_1_n76) );
  OAI22_X1 SBOX_s2_mul1_1_1_U16 ( .A1(SBOX_stage1Out[15]), .A2(
        SBOX_stage1Out[14]), .B1(SBOX_stage1Out[11]), .B2(SBOX_stage1Out[10]), 
        .ZN(SBOX_s2_mul1_1_1_n61) );
  INV_X1 SBOX_s2_mul1_1_1_U14 ( .A(SBOX_s2_mul1_1_1_n72), .ZN(
        SBOX_s2_mul1_1_1_n59) );
  INV_X1 SBOX_s2_mul1_1_1_U13 ( .A(SBOX_s2_mul1_1_1_n70), .ZN(
        SBOX_s2_mul1_1_1_n58) );
  XNOR2_X1 SBOX_s2_mul1_1_1_U12 ( .A(SBOX_s2_mul1_1_1_n56), .B(
        SBOX_s2_mul1_1_1_n71), .ZN(SBOX_s2_mul1_1_1_n57) );
  NAND2_X1 SBOX_s2_mul1_1_1_U11 ( .A1(SBOX_s2_mul1_1_1_n72), .A2(
        SBOX_s2_mul1_1_1_n73), .ZN(SBOX_s2_mul1_1_1_n56) );
  XNOR2_X1 SBOX_s2_mul1_1_1_U10 ( .A(SBOX_s2_mul1_1_1_n54), .B(
        SBOX_s2_mul1_1_1_n55), .ZN(SBOX_s2_mul1_1_1_n75) );
  NAND2_X1 SBOX_s2_mul1_1_1_U9 ( .A1(SBOX_s2_mul1_1_1_n70), .A2(
        SBOX_s2_mul1_1_1_n72), .ZN(SBOX_s2_mul1_1_1_n55) );
  NOR2_X1 SBOX_s2_mul1_1_1_U8 ( .A1(SBOX_s2_mul1_1_1_n73), .A2(
        SBOX_s2_mul1_1_1_n71), .ZN(SBOX_s2_mul1_1_1_n54) );
  AOI221_X1 SBOX_s2_mul1_1_1_U7 ( .B1(SBOX_stage1Out[13]), .B2(
        SBOX_stage1Out[12]), .C1(SBOX_stage1Out[8]), .C2(SBOX_stage1Out[9]), 
        .A(SBOX_s2_mul1_1_1_n53), .ZN(SBOX_s2_mul1_1_1_n74) );
  OAI22_X1 SBOX_s2_mul1_1_1_U6 ( .A1(SBOX_stage1Out[13]), .A2(
        SBOX_stage1Out[12]), .B1(SBOX_stage1Out[9]), .B2(SBOX_stage1Out[8]), 
        .ZN(SBOX_s2_mul1_1_1_n53) );
  XNOR2_X1 SBOX_s2_mul1_1_1_U5 ( .A(SBOX_stage1Out[12]), .B(SBOX_stage1Out[14]), .ZN(SBOX_s2_mul1_1_1_n71) );
  XOR2_X1 SBOX_s2_mul1_1_1_U4 ( .A(SBOX_stage1Out[13]), .B(SBOX_stage1Out[15]), 
        .Z(SBOX_s2_mul1_1_1_n72) );
  XNOR2_X1 SBOX_s2_mul1_1_1_U3 ( .A(SBOX_stage1Out[8]), .B(SBOX_stage1Out[10]), 
        .ZN(SBOX_s2_mul1_1_1_n73) );
  XOR2_X1 SBOX_s2_mul1_1_1_U2 ( .A(SBOX_stage1Out[9]), .B(SBOX_stage1Out[11]), 
        .Z(SBOX_s2_mul1_1_1_n70) );
  OAI33_X1 SBOX_s2_mul1_1_1_U1 ( .A1(1'b0), .A2(SBOX_s2_mul1_1_1_n57), .A3(
        SBOX_s2_mul1_1_1_n58), .B1(SBOX_s2_mul1_1_1_n70), .B2(
        SBOX_s2_mul1_1_1_n73), .B3(SBOX_s2_mul1_1_1_n59), .ZN(
        SBOX_s2_mul1_1_1_n77) );
  XNOR2_X1 SBOX_s2_mul1_1_0_U29 ( .A(SBOX_s2_mul1_1_0_n67), .B(
        SBOX_s2_mul1_1_0_n68), .ZN(SBOX_s2_xorResult[7]) );
  XOR2_X1 SBOX_s2_mul1_1_0_U28 ( .A(SBOX_s2_mul1_1_0_n77), .B(
        SBOX_s2_mul1_1_0_n76), .Z(SBOX_s2_mul1_1_0_n68) );
  NAND2_X1 SBOX_s2_mul1_1_0_U27 ( .A1(SBOX_stage1Out[3]), .A2(
        SBOX_stage1Out[15]), .ZN(SBOX_s2_mul1_1_0_n67) );
  XNOR2_X1 SBOX_s2_mul1_1_0_U26 ( .A(SBOX_s2_mul1_1_0_n65), .B(
        SBOX_s2_mul1_1_0_n66), .ZN(SBOX_s2_xorResult[6]) );
  XOR2_X1 SBOX_s2_mul1_1_0_U25 ( .A(SBOX_s2_mul1_1_0_n75), .B(
        SBOX_s2_mul1_1_0_n76), .Z(SBOX_s2_mul1_1_0_n66) );
  NAND2_X1 SBOX_s2_mul1_1_0_U24 ( .A1(SBOX_stage1Out[2]), .A2(
        SBOX_stage1Out[14]), .ZN(SBOX_s2_mul1_1_0_n65) );
  XNOR2_X1 SBOX_s2_mul1_1_0_U23 ( .A(SBOX_s2_mul1_1_0_n63), .B(
        SBOX_s2_mul1_1_0_n64), .ZN(SBOX_s2_xorResult[5]) );
  XOR2_X1 SBOX_s2_mul1_1_0_U22 ( .A(SBOX_s2_mul1_1_0_n77), .B(
        SBOX_s2_mul1_1_0_n74), .Z(SBOX_s2_mul1_1_0_n64) );
  NAND2_X1 SBOX_s2_mul1_1_0_U21 ( .A1(SBOX_stage1Out[1]), .A2(
        SBOX_stage1Out[13]), .ZN(SBOX_s2_mul1_1_0_n63) );
  XNOR2_X1 SBOX_s2_mul1_1_0_U20 ( .A(SBOX_s2_mul1_1_0_n61), .B(
        SBOX_s2_mul1_1_0_n62), .ZN(SBOX_s2_xorResult[4]) );
  XOR2_X1 SBOX_s2_mul1_1_0_U19 ( .A(SBOX_s2_mul1_1_0_n74), .B(
        SBOX_s2_mul1_1_0_n75), .Z(SBOX_s2_mul1_1_0_n62) );
  NAND2_X1 SBOX_s2_mul1_1_0_U18 ( .A1(SBOX_stage1Out[0]), .A2(
        SBOX_stage1Out[12]), .ZN(SBOX_s2_mul1_1_0_n61) );
  AOI221_X1 SBOX_s2_mul1_1_0_U17 ( .B1(SBOX_stage1Out[15]), .B2(
        SBOX_stage1Out[14]), .C1(SBOX_stage1Out[2]), .C2(SBOX_stage1Out[3]), 
        .A(SBOX_s2_mul1_1_0_n60), .ZN(SBOX_s2_mul1_1_0_n76) );
  OAI22_X1 SBOX_s2_mul1_1_0_U16 ( .A1(SBOX_stage1Out[15]), .A2(
        SBOX_stage1Out[14]), .B1(SBOX_stage1Out[3]), .B2(SBOX_stage1Out[2]), 
        .ZN(SBOX_s2_mul1_1_0_n60) );
  INV_X1 SBOX_s2_mul1_1_0_U15 ( .A(SBOX_s2_mul1_1_0_n72), .ZN(
        SBOX_s2_mul1_1_0_n59) );
  INV_X1 SBOX_s2_mul1_1_0_U14 ( .A(SBOX_s2_mul1_1_0_n70), .ZN(
        SBOX_s2_mul1_1_0_n58) );
  XNOR2_X1 SBOX_s2_mul1_1_0_U13 ( .A(SBOX_s2_mul1_1_0_n56), .B(
        SBOX_s2_mul1_1_0_n71), .ZN(SBOX_s2_mul1_1_0_n57) );
  NAND2_X1 SBOX_s2_mul1_1_0_U12 ( .A1(SBOX_s2_mul1_1_0_n72), .A2(
        SBOX_s2_mul1_1_0_n73), .ZN(SBOX_s2_mul1_1_0_n56) );
  XNOR2_X1 SBOX_s2_mul1_1_0_U10 ( .A(SBOX_s2_mul1_1_0_n53), .B(
        SBOX_s2_mul1_1_0_n54), .ZN(SBOX_s2_mul1_1_0_n75) );
  NAND2_X1 SBOX_s2_mul1_1_0_U9 ( .A1(SBOX_s2_mul1_1_0_n70), .A2(
        SBOX_s2_mul1_1_0_n72), .ZN(SBOX_s2_mul1_1_0_n54) );
  NOR2_X1 SBOX_s2_mul1_1_0_U8 ( .A1(SBOX_s2_mul1_1_0_n73), .A2(
        SBOX_s2_mul1_1_0_n71), .ZN(SBOX_s2_mul1_1_0_n53) );
  OAI22_X1 SBOX_s2_mul1_1_0_U7 ( .A1(SBOX_stage1Out[0]), .A2(SBOX_stage1Out[1]), .B1(SBOX_stage1Out[13]), .B2(SBOX_stage1Out[12]), .ZN(SBOX_s2_mul1_1_0_n69)
         );
  AOI221_X1 SBOX_s2_mul1_1_0_U6 ( .B1(SBOX_stage1Out[0]), .B2(
        SBOX_stage1Out[1]), .C1(SBOX_stage1Out[12]), .C2(SBOX_stage1Out[13]), 
        .A(SBOX_s2_mul1_1_0_n69), .ZN(SBOX_s2_mul1_1_0_n74) );
  XNOR2_X1 SBOX_s2_mul1_1_0_U5 ( .A(SBOX_stage1Out[12]), .B(SBOX_stage1Out[14]), .ZN(SBOX_s2_mul1_1_0_n71) );
  XOR2_X1 SBOX_s2_mul1_1_0_U4 ( .A(SBOX_stage1Out[13]), .B(SBOX_stage1Out[15]), 
        .Z(SBOX_s2_mul1_1_0_n72) );
  XNOR2_X1 SBOX_s2_mul1_1_0_U3 ( .A(SBOX_stage1Out[0]), .B(SBOX_stage1Out[2]), 
        .ZN(SBOX_s2_mul1_1_0_n73) );
  XOR2_X1 SBOX_s2_mul1_1_0_U2 ( .A(SBOX_stage1Out[1]), .B(SBOX_stage1Out[3]), 
        .Z(SBOX_s2_mul1_1_0_n70) );
  OAI33_X1 SBOX_s2_mul1_1_0_U1 ( .A1(1'b0), .A2(SBOX_s2_mul1_1_0_n57), .A3(
        SBOX_s2_mul1_1_0_n58), .B1(SBOX_s2_mul1_1_0_n70), .B2(
        SBOX_s2_mul1_1_0_n73), .B3(SBOX_s2_mul1_1_0_n59), .ZN(
        SBOX_s2_mul1_1_0_n77) );
  XNOR2_X1 SBOX_s2_mul1_0_1_U29 ( .A(SBOX_s2_mul1_0_1_n67), .B(
        SBOX_s2_mul1_0_1_n68), .ZN(SBOX_s2_xorResult[3]) );
  XOR2_X1 SBOX_s2_mul1_0_1_U28 ( .A(SBOX_s2_mul1_0_1_n77), .B(
        SBOX_s2_mul1_0_1_n76), .Z(SBOX_s2_mul1_0_1_n68) );
  NAND2_X1 SBOX_s2_mul1_0_1_U27 ( .A1(SBOX_stage1Out[11]), .A2(
        SBOX_stage1Out[7]), .ZN(SBOX_s2_mul1_0_1_n67) );
  XNOR2_X1 SBOX_s2_mul1_0_1_U26 ( .A(SBOX_s2_mul1_0_1_n65), .B(
        SBOX_s2_mul1_0_1_n66), .ZN(SBOX_s2_xorResult[2]) );
  XOR2_X1 SBOX_s2_mul1_0_1_U25 ( .A(SBOX_s2_mul1_0_1_n75), .B(
        SBOX_s2_mul1_0_1_n76), .Z(SBOX_s2_mul1_0_1_n66) );
  NAND2_X1 SBOX_s2_mul1_0_1_U24 ( .A1(SBOX_stage1Out[10]), .A2(
        SBOX_stage1Out[6]), .ZN(SBOX_s2_mul1_0_1_n65) );
  XNOR2_X1 SBOX_s2_mul1_0_1_U23 ( .A(SBOX_s2_mul1_0_1_n63), .B(
        SBOX_s2_mul1_0_1_n64), .ZN(SBOX_s2_xorResult[1]) );
  XOR2_X1 SBOX_s2_mul1_0_1_U22 ( .A(SBOX_s2_mul1_0_1_n77), .B(
        SBOX_s2_mul1_0_1_n74), .Z(SBOX_s2_mul1_0_1_n64) );
  NAND2_X1 SBOX_s2_mul1_0_1_U21 ( .A1(SBOX_stage1Out[9]), .A2(
        SBOX_stage1Out[5]), .ZN(SBOX_s2_mul1_0_1_n63) );
  XNOR2_X1 SBOX_s2_mul1_0_1_U20 ( .A(SBOX_s2_mul1_0_1_n61), .B(
        SBOX_s2_mul1_0_1_n62), .ZN(SBOX_s2_xorResult[0]) );
  XOR2_X1 SBOX_s2_mul1_0_1_U19 ( .A(SBOX_s2_mul1_0_1_n74), .B(
        SBOX_s2_mul1_0_1_n75), .Z(SBOX_s2_mul1_0_1_n62) );
  NAND2_X1 SBOX_s2_mul1_0_1_U18 ( .A1(SBOX_stage1Out[8]), .A2(
        SBOX_stage1Out[4]), .ZN(SBOX_s2_mul1_0_1_n61) );
  AOI221_X1 SBOX_s2_mul1_0_1_U17 ( .B1(SBOX_stage1Out[7]), .B2(
        SBOX_stage1Out[6]), .C1(SBOX_stage1Out[10]), .C2(SBOX_stage1Out[11]), 
        .A(SBOX_s2_mul1_0_1_n60), .ZN(SBOX_s2_mul1_0_1_n76) );
  OAI22_X1 SBOX_s2_mul1_0_1_U16 ( .A1(SBOX_stage1Out[7]), .A2(
        SBOX_stage1Out[6]), .B1(SBOX_stage1Out[11]), .B2(SBOX_stage1Out[10]), 
        .ZN(SBOX_s2_mul1_0_1_n60) );
  INV_X1 SBOX_s2_mul1_0_1_U15 ( .A(SBOX_s2_mul1_0_1_n72), .ZN(
        SBOX_s2_mul1_0_1_n59) );
  INV_X1 SBOX_s2_mul1_0_1_U14 ( .A(SBOX_s2_mul1_0_1_n70), .ZN(
        SBOX_s2_mul1_0_1_n58) );
  XNOR2_X1 SBOX_s2_mul1_0_1_U13 ( .A(SBOX_s2_mul1_0_1_n56), .B(
        SBOX_s2_mul1_0_1_n71), .ZN(SBOX_s2_mul1_0_1_n57) );
  NAND2_X1 SBOX_s2_mul1_0_1_U12 ( .A1(SBOX_s2_mul1_0_1_n72), .A2(
        SBOX_s2_mul1_0_1_n73), .ZN(SBOX_s2_mul1_0_1_n56) );
  XNOR2_X1 SBOX_s2_mul1_0_1_U10 ( .A(SBOX_s2_mul1_0_1_n53), .B(
        SBOX_s2_mul1_0_1_n54), .ZN(SBOX_s2_mul1_0_1_n75) );
  NAND2_X1 SBOX_s2_mul1_0_1_U9 ( .A1(SBOX_s2_mul1_0_1_n70), .A2(
        SBOX_s2_mul1_0_1_n72), .ZN(SBOX_s2_mul1_0_1_n54) );
  NOR2_X1 SBOX_s2_mul1_0_1_U8 ( .A1(SBOX_s2_mul1_0_1_n73), .A2(
        SBOX_s2_mul1_0_1_n71), .ZN(SBOX_s2_mul1_0_1_n53) );
  OAI22_X1 SBOX_s2_mul1_0_1_U7 ( .A1(SBOX_stage1Out[8]), .A2(SBOX_stage1Out[9]), .B1(SBOX_stage1Out[5]), .B2(SBOX_stage1Out[4]), .ZN(SBOX_s2_mul1_0_1_n69) );
  AOI221_X1 SBOX_s2_mul1_0_1_U6 ( .B1(SBOX_stage1Out[8]), .B2(
        SBOX_stage1Out[9]), .C1(SBOX_stage1Out[4]), .C2(SBOX_stage1Out[5]), 
        .A(SBOX_s2_mul1_0_1_n69), .ZN(SBOX_s2_mul1_0_1_n74) );
  XNOR2_X1 SBOX_s2_mul1_0_1_U5 ( .A(SBOX_stage1Out[4]), .B(SBOX_stage1Out[6]), 
        .ZN(SBOX_s2_mul1_0_1_n71) );
  XOR2_X1 SBOX_s2_mul1_0_1_U4 ( .A(SBOX_stage1Out[5]), .B(SBOX_stage1Out[7]), 
        .Z(SBOX_s2_mul1_0_1_n72) );
  XNOR2_X1 SBOX_s2_mul1_0_1_U3 ( .A(SBOX_stage1Out[8]), .B(SBOX_stage1Out[10]), 
        .ZN(SBOX_s2_mul1_0_1_n73) );
  XOR2_X1 SBOX_s2_mul1_0_1_U2 ( .A(SBOX_stage1Out[9]), .B(SBOX_stage1Out[11]), 
        .Z(SBOX_s2_mul1_0_1_n70) );
  OAI33_X1 SBOX_s2_mul1_0_1_U1 ( .A1(1'b0), .A2(SBOX_s2_mul1_0_1_n57), .A3(
        SBOX_s2_mul1_0_1_n58), .B1(SBOX_s2_mul1_0_1_n70), .B2(
        SBOX_s2_mul1_0_1_n73), .B3(SBOX_s2_mul1_0_1_n59), .ZN(
        SBOX_s2_mul1_0_1_n77) );
  XNOR2_X1 SBOX_s2_mul1_0_0_U29 ( .A(SBOX_s2_mul1_0_0_n68), .B(
        SBOX_s2_mul1_0_0_n69), .ZN(SBOX_s2_gf2_mul_out_0__0__1_) );
  XOR2_X1 SBOX_s2_mul1_0_0_U28 ( .A(SBOX_s2_mul1_0_0_n77), .B(
        SBOX_s2_mul1_0_0_n74), .Z(SBOX_s2_mul1_0_0_n69) );
  NAND2_X1 SBOX_s2_mul1_0_0_U27 ( .A1(SBOX_stage1Out[1]), .A2(
        SBOX_stage1Out[5]), .ZN(SBOX_s2_mul1_0_0_n68) );
  XNOR2_X1 SBOX_s2_mul1_0_0_U26 ( .A(SBOX_s2_mul1_0_0_n66), .B(
        SBOX_s2_mul1_0_0_n67), .ZN(SBOX_s2_gf2_mul_out_0__0__2_) );
  XOR2_X1 SBOX_s2_mul1_0_0_U25 ( .A(SBOX_s2_mul1_0_0_n75), .B(
        SBOX_s2_mul1_0_0_n76), .Z(SBOX_s2_mul1_0_0_n67) );
  NAND2_X1 SBOX_s2_mul1_0_0_U24 ( .A1(SBOX_stage1Out[2]), .A2(
        SBOX_stage1Out[6]), .ZN(SBOX_s2_mul1_0_0_n66) );
  XNOR2_X1 SBOX_s2_mul1_0_0_U23 ( .A(SBOX_s2_mul1_0_0_n64), .B(
        SBOX_s2_mul1_0_0_n65), .ZN(SBOX_s2_gf2_mul_out_0__0__3_) );
  XOR2_X1 SBOX_s2_mul1_0_0_U22 ( .A(SBOX_s2_mul1_0_0_n77), .B(
        SBOX_s2_mul1_0_0_n76), .Z(SBOX_s2_mul1_0_0_n65) );
  NAND2_X1 SBOX_s2_mul1_0_0_U21 ( .A1(SBOX_stage1Out[3]), .A2(
        SBOX_stage1Out[7]), .ZN(SBOX_s2_mul1_0_0_n64) );
  XNOR2_X1 SBOX_s2_mul1_0_0_U20 ( .A(SBOX_s2_mul1_0_0_n62), .B(
        SBOX_s2_mul1_0_0_n63), .ZN(SBOX_s2_gf2_mul_out_0__0__0_) );
  XOR2_X1 SBOX_s2_mul1_0_0_U19 ( .A(SBOX_s2_mul1_0_0_n74), .B(
        SBOX_s2_mul1_0_0_n75), .Z(SBOX_s2_mul1_0_0_n63) );
  NAND2_X1 SBOX_s2_mul1_0_0_U18 ( .A1(SBOX_stage1Out[0]), .A2(
        SBOX_stage1Out[4]), .ZN(SBOX_s2_mul1_0_0_n62) );
  AOI221_X1 SBOX_s2_mul1_0_0_U17 ( .B1(SBOX_stage1Out[7]), .B2(
        SBOX_stage1Out[6]), .C1(SBOX_stage1Out[2]), .C2(SBOX_stage1Out[3]), 
        .A(SBOX_s2_mul1_0_0_n61), .ZN(SBOX_s2_mul1_0_0_n76) );
  OAI22_X1 SBOX_s2_mul1_0_0_U16 ( .A1(SBOX_stage1Out[7]), .A2(
        SBOX_stage1Out[6]), .B1(SBOX_stage1Out[3]), .B2(SBOX_stage1Out[2]), 
        .ZN(SBOX_s2_mul1_0_0_n61) );
  INV_X1 SBOX_s2_mul1_0_0_U15 ( .A(SBOX_s2_mul1_0_0_n72), .ZN(
        SBOX_s2_mul1_0_0_n60) );
  INV_X1 SBOX_s2_mul1_0_0_U14 ( .A(SBOX_s2_mul1_0_0_n70), .ZN(
        SBOX_s2_mul1_0_0_n59) );
  XNOR2_X1 SBOX_s2_mul1_0_0_U13 ( .A(SBOX_s2_mul1_0_0_n57), .B(
        SBOX_s2_mul1_0_0_n71), .ZN(SBOX_s2_mul1_0_0_n58) );
  NAND2_X1 SBOX_s2_mul1_0_0_U12 ( .A1(SBOX_s2_mul1_0_0_n72), .A2(
        SBOX_s2_mul1_0_0_n73), .ZN(SBOX_s2_mul1_0_0_n57) );
  XNOR2_X1 SBOX_s2_mul1_0_0_U10 ( .A(SBOX_s2_mul1_0_0_n54), .B(
        SBOX_s2_mul1_0_0_n55), .ZN(SBOX_s2_mul1_0_0_n75) );
  NAND2_X1 SBOX_s2_mul1_0_0_U9 ( .A1(SBOX_s2_mul1_0_0_n70), .A2(
        SBOX_s2_mul1_0_0_n72), .ZN(SBOX_s2_mul1_0_0_n55) );
  NOR2_X1 SBOX_s2_mul1_0_0_U8 ( .A1(SBOX_s2_mul1_0_0_n73), .A2(
        SBOX_s2_mul1_0_0_n71), .ZN(SBOX_s2_mul1_0_0_n54) );
  AOI221_X1 SBOX_s2_mul1_0_0_U7 ( .B1(SBOX_stage1Out[5]), .B2(
        SBOX_stage1Out[4]), .C1(SBOX_stage1Out[0]), .C2(SBOX_stage1Out[1]), 
        .A(SBOX_s2_mul1_0_0_n53), .ZN(SBOX_s2_mul1_0_0_n74) );
  OAI22_X1 SBOX_s2_mul1_0_0_U6 ( .A1(SBOX_stage1Out[5]), .A2(SBOX_stage1Out[4]), .B1(SBOX_stage1Out[1]), .B2(SBOX_stage1Out[0]), .ZN(SBOX_s2_mul1_0_0_n53) );
  XNOR2_X1 SBOX_s2_mul1_0_0_U5 ( .A(SBOX_stage1Out[4]), .B(SBOX_stage1Out[6]), 
        .ZN(SBOX_s2_mul1_0_0_n71) );
  XOR2_X1 SBOX_s2_mul1_0_0_U4 ( .A(SBOX_stage1Out[5]), .B(SBOX_stage1Out[7]), 
        .Z(SBOX_s2_mul1_0_0_n72) );
  XNOR2_X1 SBOX_s2_mul1_0_0_U3 ( .A(SBOX_stage1Out[0]), .B(SBOX_stage1Out[2]), 
        .ZN(SBOX_s2_mul1_0_0_n73) );
  XOR2_X1 SBOX_s2_mul1_0_0_U2 ( .A(SBOX_stage1Out[1]), .B(SBOX_stage1Out[3]), 
        .Z(SBOX_s2_mul1_0_0_n70) );
  OAI33_X1 SBOX_s2_mul1_0_0_U1 ( .A1(1'b0), .A2(SBOX_s2_mul1_0_0_n58), .A3(
        SBOX_s2_mul1_0_0_n59), .B1(SBOX_s2_mul1_0_0_n70), .B2(
        SBOX_s2_mul1_0_0_n73), .B3(SBOX_s2_mul1_0_0_n60), .ZN(
        SBOX_s2_mul1_0_0_n77) );
  XOR2_X1 SBOX_s2_compr_0_0_U4 ( .A(SBOX_s2_regOut_0__1__3_), .B(
        SBOX_s2_regOut_0__2__3_), .Z(SBOX_stage2Out[7]) );
  XOR2_X1 SBOX_s2_compr_0_0_U3 ( .A(SBOX_s2_regOut_0__1__2_), .B(
        SBOX_s2_regOut_0__2__2_), .Z(SBOX_stage2Out[6]) );
  XOR2_X1 SBOX_s2_compr_0_0_U2 ( .A(SBOX_s2_regOut_0__1__1_), .B(
        SBOX_s2_regOut_0__2__1_), .Z(SBOX_stage2Out[5]) );
  XOR2_X1 SBOX_s2_compr_0_0_U1 ( .A(SBOX_s2_regOut_0__1__0_), .B(
        SBOX_s2_regOut_0__2__0_), .Z(SBOX_stage2Out[4]) );
  XOR2_X1 SBOX_s2_compr_1_0_U4 ( .A(SBOX_s2_regOut_1__1__3_), .B(
        SBOX_s2_regOut_1__2__3_), .Z(SBOX_stage2Out[19]) );
  XOR2_X1 SBOX_s2_compr_1_0_U3 ( .A(SBOX_s2_regOut_1__1__2_), .B(
        SBOX_s2_regOut_1__2__2_), .Z(SBOX_stage2Out[18]) );
  XOR2_X1 SBOX_s2_compr_1_0_U2 ( .A(SBOX_s2_regOut_1__1__1_), .B(
        SBOX_s2_regOut_1__2__1_), .Z(SBOX_stage2Out[17]) );
  XOR2_X1 SBOX_s2_compr_1_0_U1 ( .A(SBOX_s2_regOut_1__1__0_), .B(
        SBOX_s2_regOut_1__2__0_), .Z(SBOX_stage2Out[16]) );
  XOR2_X1 SBOX_s3_U22 ( .A(SBOX_stage2Out[17]), .B(SBOX_stage2Out[19]), .Z(
        SBOX_s3_scale_out[3]) );
  XOR2_X1 SBOX_s3_U21 ( .A(SBOX_stage2Out[16]), .B(SBOX_stage2Out[18]), .Z(
        SBOX_s3_scale_in[1]) );
  XOR2_X1 SBOX_s3_U20 ( .A(SBOX_s3_scale_out[2]), .B(SBOX_s3_n8), .Z(
        SBOX_s3_refreshed[6]) );
  XNOR2_X1 SBOX_s3_U19 ( .A(SBOX_s3_n6), .B(SBOX_s3_n7), .ZN(SBOX_s3_n8) );
  XNOR2_X1 SBOX_s3_U18 ( .A(SBOX_s3_gf2_mul_out_1__1__0_), .B(randomS3[4]), 
        .ZN(SBOX_s3_n7) );
  XOR2_X1 SBOX_s3_U17 ( .A(randomS3[0]), .B(randomS3[2]), .Z(SBOX_s3_n6) );
  XOR2_X1 SBOX_s3_U16 ( .A(SBOX_stage2Out[4]), .B(SBOX_stage2Out[6]), .Z(
        SBOX_s3_scale_in[0]) );
  XNOR2_X1 SBOX_s3_U15 ( .A(SBOX_s3_n5), .B(SBOX_s3_scale_out[0]), .ZN(
        SBOX_s3_refreshed[0]) );
  XNOR2_X1 SBOX_s3_U14 ( .A(randomS3[0]), .B(SBOX_s3_gf2_mul_out_0__0__0_), 
        .ZN(SBOX_s3_n5) );
  XOR2_X1 SBOX_s3_U13 ( .A(SBOX_s3_scale_out[3]), .B(SBOX_s3_n4), .Z(
        SBOX_s3_refreshed[7]) );
  XNOR2_X1 SBOX_s3_U12 ( .A(SBOX_s3_n2), .B(SBOX_s3_n3), .ZN(SBOX_s3_n4) );
  XNOR2_X1 SBOX_s3_U11 ( .A(SBOX_s3_gf2_mul_out_1__1__1_), .B(randomS3[5]), 
        .ZN(SBOX_s3_n3) );
  XOR2_X1 SBOX_s3_U10 ( .A(randomS3[1]), .B(randomS3[3]), .Z(SBOX_s3_n2) );
  XNOR2_X1 SBOX_s3_U9 ( .A(SBOX_s3_n1), .B(SBOX_s3_scale_out[1]), .ZN(
        SBOX_s3_refreshed[1]) );
  XNOR2_X1 SBOX_s3_U8 ( .A(randomS3[1]), .B(SBOX_s3_gf2_mul_out_0__0__1_), 
        .ZN(SBOX_s3_n1) );
  XOR2_X1 SBOX_s3_U7 ( .A(randomS3[4]), .B(SBOX_s3_xorResult[2]), .Z(
        SBOX_s3_refreshed[4]) );
  XOR2_X1 SBOX_s3_U6 ( .A(randomS3[2]), .B(SBOX_s3_xorResult[0]), .Z(
        SBOX_s3_refreshed[2]) );
  XOR2_X1 SBOX_s3_U5 ( .A(randomS3[5]), .B(SBOX_s3_xorResult[3]), .Z(
        SBOX_s3_refreshed[5]) );
  XOR2_X1 SBOX_s3_U4 ( .A(randomS3[3]), .B(SBOX_s3_xorResult[1]), .Z(
        SBOX_s3_refreshed[3]) );
  XOR2_X1 SBOX_s3_U3 ( .A(SBOX_stage2Out[5]), .B(SBOX_stage2Out[7]), .Z(
        SBOX_s3_scale_out[1]) );
  DFF_X1 SBOX_s3_regOut_reg_0__0__0_ ( .D(SBOX_stage2Out[0]), .CK(ClkxCI), .Q(
        SBOX_stage3Out[0]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__0__1_ ( .D(SBOX_stage2Out[1]), .CK(ClkxCI), .Q(
        SBOX_stage3Out[1]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__1__0_ ( .D(SBOX_stage2Out[2]), .CK(ClkxCI), .Q(
        SBOX_stage3Out[2]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__1__1_ ( .D(SBOX_stage2Out[3]), .CK(ClkxCI), .Q(
        SBOX_stage3Out[3]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__2__0_ ( .D(SBOX_stage2Out[4]), .CK(ClkxCI), .Q(
        SBOX_stage3Out[4]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__2__1_ ( .D(SBOX_stage2Out[5]), .CK(ClkxCI), .Q(
        SBOX_stage3Out[5]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__3__0_ ( .D(SBOX_s3_refreshed[0]), .CK(ClkxCI), 
        .Q(SBOX_s3_regOut_0__3__0_), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__3__1_ ( .D(SBOX_s3_refreshed[1]), .CK(ClkxCI), 
        .Q(SBOX_s3_regOut_0__3__1_), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__4__0_ ( .D(SBOX_s3_refreshed[2]), .CK(ClkxCI), 
        .Q(SBOX_s3_regOut_0__4__0_), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__4__1_ ( .D(SBOX_s3_refreshed[3]), .CK(ClkxCI), 
        .Q(SBOX_s3_regOut_0__4__1_), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__5__0_ ( .D(SBOX_stage2Out[6]), .CK(ClkxCI), .Q(
        SBOX_stage3Out[6]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__5__1_ ( .D(SBOX_stage2Out[7]), .CK(ClkxCI), .Q(
        SBOX_stage3Out[7]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__6__0_ ( .D(SBOX_stage2Out[8]), .CK(ClkxCI), .Q(
        SBOX_stage3Out[8]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__6__1_ ( .D(SBOX_stage2Out[9]), .CK(ClkxCI), .Q(
        SBOX_stage3Out[9]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__7__0_ ( .D(SBOX_stage2Out[10]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[10]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_0__7__1_ ( .D(SBOX_stage2Out[11]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[11]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__0__0_ ( .D(SBOX_stage2Out[12]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[12]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__0__1_ ( .D(SBOX_stage2Out[13]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[13]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__1__0_ ( .D(SBOX_stage2Out[14]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[14]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__1__1_ ( .D(SBOX_stage2Out[15]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[15]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__2__0_ ( .D(SBOX_stage2Out[16]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[16]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__2__1_ ( .D(SBOX_stage2Out[17]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[17]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__3__0_ ( .D(SBOX_s3_refreshed[4]), .CK(ClkxCI), 
        .Q(SBOX_s3_regOut_1__3__0_), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__3__1_ ( .D(SBOX_s3_refreshed[5]), .CK(ClkxCI), 
        .Q(SBOX_s3_regOut_1__3__1_), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__4__0_ ( .D(SBOX_s3_refreshed[6]), .CK(ClkxCI), 
        .Q(SBOX_s3_regOut_1__4__0_), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__4__1_ ( .D(SBOX_s3_refreshed[7]), .CK(ClkxCI), 
        .Q(SBOX_s3_regOut_1__4__1_), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__5__0_ ( .D(SBOX_stage2Out[18]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[18]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__5__1_ ( .D(SBOX_stage2Out[19]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[19]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__6__0_ ( .D(SBOX_stage2Out[20]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[20]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__6__1_ ( .D(SBOX_stage2Out[21]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[21]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__7__0_ ( .D(SBOX_stage2Out[22]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[22]), .QN() );
  DFF_X1 SBOX_s3_regOut_reg_1__7__1_ ( .D(SBOX_stage2Out[23]), .CK(ClkxCI), 
        .Q(SBOX_stage3Out[23]), .QN() );
  XOR2_X1 SBOX_s3_sqsc_1_U1 ( .A(SBOX_s3_scale_in[1]), .B(SBOX_s3_scale_out[3]), .Z(SBOX_s3_scale_out[2]) );
  XOR2_X1 SBOX_s3_sqsc_0_U1 ( .A(SBOX_s3_scale_in[0]), .B(SBOX_s3_scale_out[1]), .Z(SBOX_s3_scale_out[0]) );
  XNOR2_X1 SBOX_s3_mul1_1_1_U6 ( .A(SBOX_s3_mul1_1_1_n13), .B(
        SBOX_s3_mul1_1_1_n14), .ZN(SBOX_s3_gf2_mul_out_1__1__0_) );
  NAND2_X1 SBOX_s3_mul1_1_1_U5 ( .A1(SBOX_stage2Out[18]), .A2(
        SBOX_stage2Out[16]), .ZN(SBOX_s3_mul1_1_1_n13) );
  XNOR2_X1 SBOX_s3_mul1_1_1_U4 ( .A(SBOX_s3_mul1_1_1_n12), .B(
        SBOX_s3_mul1_1_1_n14), .ZN(SBOX_s3_gf2_mul_out_1__1__1_) );
  NAND2_X1 SBOX_s3_mul1_1_1_U3 ( .A1(SBOX_stage2Out[19]), .A2(
        SBOX_stage2Out[17]), .ZN(SBOX_s3_mul1_1_1_n12) );
  AOI221_X1 SBOX_s3_mul1_1_1_U2 ( .B1(SBOX_stage2Out[18]), .B2(
        SBOX_stage2Out[19]), .C1(SBOX_stage2Out[16]), .C2(SBOX_stage2Out[17]), 
        .A(SBOX_s3_mul1_1_1_n11), .ZN(SBOX_s3_mul1_1_1_n14) );
  OAI22_X1 SBOX_s3_mul1_1_1_U1 ( .A1(SBOX_stage2Out[18]), .A2(
        SBOX_stage2Out[19]), .B1(SBOX_stage2Out[17]), .B2(SBOX_stage2Out[16]), 
        .ZN(SBOX_s3_mul1_1_1_n11) );
  AOI221_X1 SBOX_s3_mul1_1_0_U6 ( .B1(SBOX_stage2Out[4]), .B2(
        SBOX_stage2Out[5]), .C1(SBOX_stage2Out[19]), .C2(SBOX_stage2Out[18]), 
        .A(SBOX_s3_mul1_1_0_n13), .ZN(SBOX_s3_mul1_1_0_n14) );
  OAI22_X1 SBOX_s3_mul1_1_0_U5 ( .A1(SBOX_stage2Out[4]), .A2(SBOX_stage2Out[5]), .B1(SBOX_stage2Out[18]), .B2(SBOX_stage2Out[19]), .ZN(SBOX_s3_mul1_1_0_n13)
         );
  XNOR2_X1 SBOX_s3_mul1_1_0_U4 ( .A(SBOX_s3_mul1_1_0_n12), .B(
        SBOX_s3_mul1_1_0_n14), .ZN(SBOX_s3_xorResult[2]) );
  NAND2_X1 SBOX_s3_mul1_1_0_U3 ( .A1(SBOX_stage2Out[18]), .A2(
        SBOX_stage2Out[4]), .ZN(SBOX_s3_mul1_1_0_n12) );
  XNOR2_X1 SBOX_s3_mul1_1_0_U2 ( .A(SBOX_s3_mul1_1_0_n11), .B(
        SBOX_s3_mul1_1_0_n14), .ZN(SBOX_s3_xorResult[3]) );
  NAND2_X1 SBOX_s3_mul1_1_0_U1 ( .A1(SBOX_stage2Out[19]), .A2(
        SBOX_stage2Out[5]), .ZN(SBOX_s3_mul1_1_0_n11) );
  AOI221_X1 SBOX_s3_mul1_0_1_U6 ( .B1(SBOX_stage2Out[16]), .B2(
        SBOX_stage2Out[17]), .C1(SBOX_stage2Out[7]), .C2(SBOX_stage2Out[6]), 
        .A(SBOX_s3_mul1_0_1_n13), .ZN(SBOX_s3_mul1_0_1_n14) );
  OAI22_X1 SBOX_s3_mul1_0_1_U5 ( .A1(SBOX_stage2Out[16]), .A2(
        SBOX_stage2Out[17]), .B1(SBOX_stage2Out[6]), .B2(SBOX_stage2Out[7]), 
        .ZN(SBOX_s3_mul1_0_1_n13) );
  XNOR2_X1 SBOX_s3_mul1_0_1_U4 ( .A(SBOX_s3_mul1_0_1_n12), .B(
        SBOX_s3_mul1_0_1_n14), .ZN(SBOX_s3_xorResult[0]) );
  NAND2_X1 SBOX_s3_mul1_0_1_U3 ( .A1(SBOX_stage2Out[6]), .A2(
        SBOX_stage2Out[16]), .ZN(SBOX_s3_mul1_0_1_n12) );
  XNOR2_X1 SBOX_s3_mul1_0_1_U2 ( .A(SBOX_s3_mul1_0_1_n11), .B(
        SBOX_s3_mul1_0_1_n14), .ZN(SBOX_s3_xorResult[1]) );
  NAND2_X1 SBOX_s3_mul1_0_1_U1 ( .A1(SBOX_stage2Out[7]), .A2(
        SBOX_stage2Out[17]), .ZN(SBOX_s3_mul1_0_1_n11) );
  XNOR2_X1 SBOX_s3_mul1_0_0_U6 ( .A(SBOX_s3_mul1_0_0_n13), .B(
        SBOX_s3_mul1_0_0_n14), .ZN(SBOX_s3_gf2_mul_out_0__0__0_) );
  NAND2_X1 SBOX_s3_mul1_0_0_U5 ( .A1(SBOX_stage2Out[6]), .A2(SBOX_stage2Out[4]), .ZN(SBOX_s3_mul1_0_0_n13) );
  XNOR2_X1 SBOX_s3_mul1_0_0_U4 ( .A(SBOX_s3_mul1_0_0_n12), .B(
        SBOX_s3_mul1_0_0_n14), .ZN(SBOX_s3_gf2_mul_out_0__0__1_) );
  NAND2_X1 SBOX_s3_mul1_0_0_U3 ( .A1(SBOX_stage2Out[7]), .A2(SBOX_stage2Out[5]), .ZN(SBOX_s3_mul1_0_0_n12) );
  AOI221_X1 SBOX_s3_mul1_0_0_U2 ( .B1(SBOX_stage2Out[6]), .B2(
        SBOX_stage2Out[7]), .C1(SBOX_stage2Out[4]), .C2(SBOX_stage2Out[5]), 
        .A(SBOX_s3_mul1_0_0_n11), .ZN(SBOX_s3_mul1_0_0_n14) );
  OAI22_X1 SBOX_s3_mul1_0_0_U1 ( .A1(SBOX_stage2Out[6]), .A2(SBOX_stage2Out[7]), .B1(SBOX_stage2Out[5]), .B2(SBOX_stage2Out[4]), .ZN(SBOX_s3_mul1_0_0_n11) );
  XOR2_X2 SBOX_s3_compr_0_0_U2 ( .A(SBOX_s3_regOut_0__3__0_), .B(
        SBOX_s3_regOut_0__4__0_), .Z(SBOX_s4_inv_out_0__1_) );
  XOR2_X2 SBOX_s3_compr_0_0_U1 ( .A(SBOX_s3_regOut_0__3__1_), .B(
        SBOX_s3_regOut_0__4__1_), .Z(SBOX_s4_inv_out_0__0_) );
  XOR2_X2 SBOX_s3_compr_1_0_U2 ( .A(SBOX_s3_regOut_1__3__0_), .B(
        SBOX_s3_regOut_1__4__0_), .Z(SBOX_s4_inv_out_1__1_) );
  XOR2_X2 SBOX_s3_compr_1_0_U1 ( .A(SBOX_s3_regOut_1__3__1_), .B(
        SBOX_s3_regOut_1__4__1_), .Z(SBOX_s4_inv_out_1__0_) );
  XOR2_X1 SBOX_s4_U26 ( .A(randomS4[4]), .B(SBOX_s4_concat[4]), .Z(
        SBOX_s4_refreshed[4]) );
  XOR2_X1 SBOX_s4_U25 ( .A(randomS4[2]), .B(SBOX_s4_concat[2]), .Z(
        SBOX_s4_refreshed[2]) );
  XNOR2_X1 SBOX_s4_U24 ( .A(SBOX_s4_n7), .B(SBOX_s4_n8), .ZN(
        SBOX_s4_refreshed[15]) );
  XNOR2_X1 SBOX_s4_U23 ( .A(randomS4[3]), .B(randomS4[7]), .ZN(SBOX_s4_n8) );
  XOR2_X1 SBOX_s4_U22 ( .A(randomS4[11]), .B(SBOX_s4_concat[15]), .Z(
        SBOX_s4_n7) );
  XOR2_X1 SBOX_s4_U21 ( .A(randomS4[9]), .B(SBOX_s4_concat[9]), .Z(
        SBOX_s4_refreshed[9]) );
  XNOR2_X1 SBOX_s4_U20 ( .A(SBOX_s4_n5), .B(SBOX_s4_n6), .ZN(
        SBOX_s4_refreshed[14]) );
  XNOR2_X1 SBOX_s4_U19 ( .A(randomS4[2]), .B(randomS4[6]), .ZN(SBOX_s4_n6) );
  XOR2_X1 SBOX_s4_U18 ( .A(randomS4[10]), .B(SBOX_s4_concat[14]), .Z(
        SBOX_s4_n5) );
  XOR2_X1 SBOX_s4_U17 ( .A(randomS4[8]), .B(SBOX_s4_concat[8]), .Z(
        SBOX_s4_refreshed[8]) );
  XNOR2_X1 SBOX_s4_U16 ( .A(SBOX_s4_n3), .B(SBOX_s4_n4), .ZN(
        SBOX_s4_refreshed[13]) );
  XNOR2_X1 SBOX_s4_U15 ( .A(randomS4[1]), .B(randomS4[5]), .ZN(SBOX_s4_n4) );
  XOR2_X1 SBOX_s4_U14 ( .A(randomS4[9]), .B(SBOX_s4_concat[13]), .Z(SBOX_s4_n3) );
  XOR2_X1 SBOX_s4_U13 ( .A(randomS4[11]), .B(SBOX_s4_concat[11]), .Z(
        SBOX_s4_refreshed[11]) );
  XNOR2_X1 SBOX_s4_U12 ( .A(SBOX_s4_n1), .B(SBOX_s4_n2), .ZN(
        SBOX_s4_refreshed[12]) );
  XNOR2_X1 SBOX_s4_U11 ( .A(randomS4[0]), .B(randomS4[4]), .ZN(SBOX_s4_n2) );
  XOR2_X1 SBOX_s4_U10 ( .A(randomS4[8]), .B(SBOX_s4_concat[12]), .Z(SBOX_s4_n1) );
  XOR2_X1 SBOX_s4_U9 ( .A(randomS4[10]), .B(SBOX_s4_concat[10]), .Z(
        SBOX_s4_refreshed[10]) );
  XOR2_X1 SBOX_s4_U8 ( .A(randomS4[7]), .B(SBOX_s4_concat[7]), .Z(
        SBOX_s4_refreshed[7]) );
  XOR2_X1 SBOX_s4_U7 ( .A(randomS4[1]), .B(SBOX_s4_concat[1]), .Z(
        SBOX_s4_refreshed[1]) );
  XOR2_X1 SBOX_s4_U6 ( .A(randomS4[6]), .B(SBOX_s4_concat[6]), .Z(
        SBOX_s4_refreshed[6]) );
  XOR2_X1 SBOX_s4_U5 ( .A(randomS4[0]), .B(SBOX_s4_concat[0]), .Z(
        SBOX_s4_refreshed[0]) );
  XOR2_X1 SBOX_s4_U4 ( .A(randomS4[5]), .B(SBOX_s4_concat[5]), .Z(
        SBOX_s4_refreshed[5]) );
  XOR2_X1 SBOX_s4_U3 ( .A(randomS4[3]), .B(SBOX_s4_concat[3]), .Z(
        SBOX_s4_refreshed[3]) );
  DFF_X1 SBOX_s4_regOut_reg_0__0__0_ ( .D(SBOX_stage3Out[0]), .CK(ClkxCI), .Q(
        SBOX_stage4Out[0]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__0__1_ ( .D(SBOX_stage3Out[1]), .CK(ClkxCI), .Q(
        SBOX_stage4Out[1]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__0__2_ ( .D(SBOX_stage3Out[2]), .CK(ClkxCI), .Q(
        SBOX_stage4Out[2]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__0__3_ ( .D(SBOX_stage3Out[3]), .CK(ClkxCI), .Q(
        SBOX_stage4Out[3]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__1__0_ ( .D(SBOX_s4_refreshed[0]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_0__1__0_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__1__1_ ( .D(SBOX_s4_refreshed[1]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_0__1__1_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__1__2_ ( .D(SBOX_s4_refreshed[2]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_0__1__2_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__1__3_ ( .D(SBOX_s4_refreshed[3]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_0__1__3_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__2__0_ ( .D(SBOX_s4_refreshed[4]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_0__2__0_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__2__1_ ( .D(SBOX_s4_refreshed[5]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_0__2__1_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__2__2_ ( .D(SBOX_s4_refreshed[6]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_0__2__2_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__2__3_ ( .D(SBOX_s4_refreshed[7]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_0__2__3_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__3__0_ ( .D(SBOX_stage3Out[8]), .CK(ClkxCI), .Q(
        SBOX_stage4Out[8]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__3__1_ ( .D(SBOX_stage3Out[9]), .CK(ClkxCI), .Q(
        SBOX_stage4Out[9]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__3__2_ ( .D(SBOX_stage3Out[10]), .CK(ClkxCI), 
        .Q(SBOX_stage4Out[10]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_0__3__3_ ( .D(SBOX_stage3Out[11]), .CK(ClkxCI), 
        .Q(SBOX_stage4Out[11]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__0__0_ ( .D(SBOX_stage3Out[12]), .CK(ClkxCI), 
        .Q(SBOX_stage4Out[12]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__0__1_ ( .D(SBOX_stage3Out[13]), .CK(ClkxCI), 
        .Q(SBOX_stage4Out[13]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__0__2_ ( .D(SBOX_stage3Out[14]), .CK(ClkxCI), 
        .Q(SBOX_stage4Out[14]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__0__3_ ( .D(SBOX_stage3Out[15]), .CK(ClkxCI), 
        .Q(SBOX_stage4Out[15]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__1__0_ ( .D(SBOX_s4_refreshed[8]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_1__1__0_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__1__1_ ( .D(SBOX_s4_refreshed[9]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_1__1__1_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__1__2_ ( .D(SBOX_s4_refreshed[10]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_1__1__2_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__1__3_ ( .D(SBOX_s4_refreshed[11]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_1__1__3_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__2__0_ ( .D(SBOX_s4_refreshed[12]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_1__2__0_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__2__1_ ( .D(SBOX_s4_refreshed[13]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_1__2__1_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__2__2_ ( .D(SBOX_s4_refreshed[14]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_1__2__2_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__2__3_ ( .D(SBOX_s4_refreshed[15]), .CK(ClkxCI), 
        .Q(SBOX_s4_regOut_1__2__3_), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__3__0_ ( .D(SBOX_stage3Out[20]), .CK(ClkxCI), 
        .Q(SBOX_stage4Out[20]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__3__1_ ( .D(SBOX_stage3Out[21]), .CK(ClkxCI), 
        .Q(SBOX_stage4Out[21]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__3__2_ ( .D(SBOX_stage3Out[22]), .CK(ClkxCI), 
        .Q(SBOX_stage4Out[22]), .QN() );
  DFF_X1 SBOX_s4_regOut_reg_1__3__3_ ( .D(SBOX_stage3Out[23]), .CK(ClkxCI), 
        .Q(SBOX_stage4Out[23]), .QN() );
  OAI22_X1 SBOX_s4_mul1_1_1_U6 ( .A1(SBOX_s4_inv_out_1__0_), .A2(
        SBOX_s4_inv_out_1__1_), .B1(SBOX_stage3Out[18]), .B2(
        SBOX_stage3Out[19]), .ZN(SBOX_s4_mul1_1_1_n13) );
  AOI221_X1 SBOX_s4_mul1_1_1_U5 ( .B1(SBOX_s4_inv_out_1__0_), .B2(
        SBOX_s4_inv_out_1__1_), .C1(SBOX_stage3Out[19]), .C2(
        SBOX_stage3Out[18]), .A(SBOX_s4_mul1_1_1_n13), .ZN(
        SBOX_s4_mul1_1_1_n14) );
  XNOR2_X1 SBOX_s4_mul1_1_1_U4 ( .A(SBOX_s4_mul1_1_1_n12), .B(
        SBOX_s4_mul1_1_1_n14), .ZN(SBOX_s4_concat[13]) );
  NAND2_X1 SBOX_s4_mul1_1_1_U3 ( .A1(SBOX_stage3Out[19]), .A2(
        SBOX_s4_inv_out_1__1_), .ZN(SBOX_s4_mul1_1_1_n12) );
  XNOR2_X1 SBOX_s4_mul1_1_1_U2 ( .A(SBOX_s4_mul1_1_1_n11), .B(
        SBOX_s4_mul1_1_1_n14), .ZN(SBOX_s4_concat[12]) );
  NAND2_X1 SBOX_s4_mul1_1_1_U1 ( .A1(SBOX_stage3Out[18]), .A2(
        SBOX_s4_inv_out_1__0_), .ZN(SBOX_s4_mul1_1_1_n11) );
  AOI221_X1 SBOX_s4_mul1_1_0_U6 ( .B1(SBOX_s4_inv_out_0__0_), .B2(
        SBOX_s4_inv_out_0__1_), .C1(SBOX_stage3Out[19]), .C2(
        SBOX_stage3Out[18]), .A(SBOX_s4_mul1_1_0_n13), .ZN(
        SBOX_s4_mul1_1_0_n14) );
  OAI22_X1 SBOX_s4_mul1_1_0_U5 ( .A1(SBOX_s4_inv_out_0__0_), .A2(
        SBOX_s4_inv_out_0__1_), .B1(SBOX_stage3Out[18]), .B2(
        SBOX_stage3Out[19]), .ZN(SBOX_s4_mul1_1_0_n13) );
  XNOR2_X1 SBOX_s4_mul1_1_0_U4 ( .A(SBOX_s4_mul1_1_0_n12), .B(
        SBOX_s4_mul1_1_0_n14), .ZN(SBOX_s4_concat[9]) );
  NAND2_X1 SBOX_s4_mul1_1_0_U3 ( .A1(SBOX_stage3Out[19]), .A2(
        SBOX_s4_inv_out_0__1_), .ZN(SBOX_s4_mul1_1_0_n12) );
  XNOR2_X1 SBOX_s4_mul1_1_0_U2 ( .A(SBOX_s4_mul1_1_0_n11), .B(
        SBOX_s4_mul1_1_0_n14), .ZN(SBOX_s4_concat[8]) );
  NAND2_X1 SBOX_s4_mul1_1_0_U1 ( .A1(SBOX_stage3Out[18]), .A2(
        SBOX_s4_inv_out_0__0_), .ZN(SBOX_s4_mul1_1_0_n11) );
  AOI221_X1 SBOX_s4_mul1_0_1_U6 ( .B1(SBOX_s4_inv_out_1__0_), .B2(
        SBOX_s4_inv_out_1__1_), .C1(SBOX_stage3Out[7]), .C2(SBOX_stage3Out[6]), 
        .A(SBOX_s4_mul1_0_1_n12), .ZN(SBOX_s4_mul1_0_1_n14) );
  XNOR2_X1 SBOX_s4_mul1_0_1_U5 ( .A(SBOX_s4_mul1_0_1_n11), .B(
        SBOX_s4_mul1_0_1_n14), .ZN(SBOX_s4_concat[5]) );
  NAND2_X1 SBOX_s4_mul1_0_1_U4 ( .A1(SBOX_stage3Out[7]), .A2(
        SBOX_s4_inv_out_1__1_), .ZN(SBOX_s4_mul1_0_1_n11) );
  NAND2_X1 SBOX_s4_mul1_0_1_U3 ( .A1(SBOX_s4_inv_out_1__0_), .A2(
        SBOX_stage3Out[6]), .ZN(SBOX_s4_mul1_0_1_n13) );
  XNOR2_X1 SBOX_s4_mul1_0_1_U2 ( .A(SBOX_s4_mul1_0_1_n14), .B(
        SBOX_s4_mul1_0_1_n13), .ZN(SBOX_s4_concat[4]) );
  OAI22_X1 SBOX_s4_mul1_0_1_U1 ( .A1(SBOX_s4_inv_out_1__0_), .A2(
        SBOX_s4_inv_out_1__1_), .B1(SBOX_stage3Out[6]), .B2(SBOX_stage3Out[7]), 
        .ZN(SBOX_s4_mul1_0_1_n12) );
  AOI221_X1 SBOX_s4_mul1_0_0_U6 ( .B1(SBOX_s4_inv_out_0__0_), .B2(
        SBOX_s4_inv_out_0__1_), .C1(SBOX_stage3Out[7]), .C2(SBOX_stage3Out[6]), 
        .A(SBOX_s4_mul1_0_0_n13), .ZN(SBOX_s4_mul1_0_0_n14) );
  XNOR2_X1 SBOX_s4_mul1_0_0_U5 ( .A(SBOX_s4_mul1_0_0_n12), .B(
        SBOX_s4_mul1_0_0_n14), .ZN(SBOX_s4_concat[1]) );
  NAND2_X1 SBOX_s4_mul1_0_0_U4 ( .A1(SBOX_stage3Out[7]), .A2(
        SBOX_s4_inv_out_0__1_), .ZN(SBOX_s4_mul1_0_0_n12) );
  XNOR2_X1 SBOX_s4_mul1_0_0_U3 ( .A(SBOX_s4_mul1_0_0_n11), .B(
        SBOX_s4_mul1_0_0_n14), .ZN(SBOX_s4_concat[0]) );
  NAND2_X1 SBOX_s4_mul1_0_0_U2 ( .A1(SBOX_stage3Out[6]), .A2(
        SBOX_s4_inv_out_0__0_), .ZN(SBOX_s4_mul1_0_0_n11) );
  OAI22_X1 SBOX_s4_mul1_0_0_U1 ( .A1(SBOX_s4_inv_out_0__0_), .A2(
        SBOX_s4_inv_out_0__1_), .B1(SBOX_stage3Out[6]), .B2(SBOX_stage3Out[7]), 
        .ZN(SBOX_s4_mul1_0_0_n13) );
  OAI22_X1 SBOX_s4_mul2_1_1_U6 ( .A1(SBOX_s4_inv_out_1__0_), .A2(
        SBOX_s4_inv_out_1__1_), .B1(SBOX_stage3Out[16]), .B2(
        SBOX_stage3Out[17]), .ZN(SBOX_s4_mul2_1_1_n13) );
  AOI221_X1 SBOX_s4_mul2_1_1_U5 ( .B1(SBOX_s4_inv_out_1__0_), .B2(
        SBOX_s4_inv_out_1__1_), .C1(SBOX_stage3Out[17]), .C2(
        SBOX_stage3Out[16]), .A(SBOX_s4_mul2_1_1_n13), .ZN(
        SBOX_s4_mul2_1_1_n14) );
  XNOR2_X1 SBOX_s4_mul2_1_1_U4 ( .A(SBOX_s4_mul2_1_1_n12), .B(
        SBOX_s4_mul2_1_1_n14), .ZN(SBOX_s4_concat[15]) );
  NAND2_X1 SBOX_s4_mul2_1_1_U3 ( .A1(SBOX_stage3Out[17]), .A2(
        SBOX_s4_inv_out_1__1_), .ZN(SBOX_s4_mul2_1_1_n12) );
  XNOR2_X1 SBOX_s4_mul2_1_1_U2 ( .A(SBOX_s4_mul2_1_1_n11), .B(
        SBOX_s4_mul2_1_1_n14), .ZN(SBOX_s4_concat[14]) );
  NAND2_X1 SBOX_s4_mul2_1_1_U1 ( .A1(SBOX_stage3Out[16]), .A2(
        SBOX_s4_inv_out_1__0_), .ZN(SBOX_s4_mul2_1_1_n11) );
  OAI22_X1 SBOX_s4_mul2_1_0_U6 ( .A1(SBOX_s4_inv_out_0__0_), .A2(
        SBOX_s4_inv_out_0__1_), .B1(SBOX_stage3Out[16]), .B2(
        SBOX_stage3Out[17]), .ZN(SBOX_s4_mul2_1_0_n13) );
  AOI221_X1 SBOX_s4_mul2_1_0_U5 ( .B1(SBOX_s4_inv_out_0__0_), .B2(
        SBOX_s4_inv_out_0__1_), .C1(SBOX_stage3Out[17]), .C2(
        SBOX_stage3Out[16]), .A(SBOX_s4_mul2_1_0_n13), .ZN(
        SBOX_s4_mul2_1_0_n14) );
  XNOR2_X1 SBOX_s4_mul2_1_0_U4 ( .A(SBOX_s4_mul2_1_0_n12), .B(
        SBOX_s4_mul2_1_0_n14), .ZN(SBOX_s4_concat[11]) );
  NAND2_X1 SBOX_s4_mul2_1_0_U3 ( .A1(SBOX_stage3Out[17]), .A2(
        SBOX_s4_inv_out_0__1_), .ZN(SBOX_s4_mul2_1_0_n12) );
  XNOR2_X1 SBOX_s4_mul2_1_0_U2 ( .A(SBOX_s4_mul2_1_0_n11), .B(
        SBOX_s4_mul2_1_0_n14), .ZN(SBOX_s4_concat[10]) );
  NAND2_X1 SBOX_s4_mul2_1_0_U1 ( .A1(SBOX_stage3Out[16]), .A2(
        SBOX_s4_inv_out_0__0_), .ZN(SBOX_s4_mul2_1_0_n11) );
  AOI221_X1 SBOX_s4_mul2_0_1_U6 ( .B1(SBOX_s4_inv_out_1__0_), .B2(
        SBOX_s4_inv_out_1__1_), .C1(SBOX_stage3Out[5]), .C2(SBOX_stage3Out[4]), 
        .A(SBOX_s4_mul2_0_1_n13), .ZN(SBOX_s4_mul2_0_1_n14) );
  XNOR2_X1 SBOX_s4_mul2_0_1_U5 ( .A(SBOX_s4_mul2_0_1_n12), .B(
        SBOX_s4_mul2_0_1_n14), .ZN(SBOX_s4_concat[7]) );
  NAND2_X1 SBOX_s4_mul2_0_1_U4 ( .A1(SBOX_stage3Out[5]), .A2(
        SBOX_s4_inv_out_1__1_), .ZN(SBOX_s4_mul2_0_1_n12) );
  XNOR2_X1 SBOX_s4_mul2_0_1_U3 ( .A(SBOX_s4_mul2_0_1_n11), .B(
        SBOX_s4_mul2_0_1_n14), .ZN(SBOX_s4_concat[6]) );
  NAND2_X1 SBOX_s4_mul2_0_1_U2 ( .A1(SBOX_stage3Out[4]), .A2(
        SBOX_s4_inv_out_1__0_), .ZN(SBOX_s4_mul2_0_1_n11) );
  OAI22_X1 SBOX_s4_mul2_0_1_U1 ( .A1(SBOX_s4_inv_out_1__0_), .A2(
        SBOX_s4_inv_out_1__1_), .B1(SBOX_stage3Out[4]), .B2(SBOX_stage3Out[5]), 
        .ZN(SBOX_s4_mul2_0_1_n13) );
  AOI221_X1 SBOX_s4_mul2_0_0_U6 ( .B1(SBOX_s4_inv_out_0__0_), .B2(
        SBOX_s4_inv_out_0__1_), .C1(SBOX_stage3Out[5]), .C2(SBOX_stage3Out[4]), 
        .A(SBOX_s4_mul2_0_0_n12), .ZN(SBOX_s4_mul2_0_0_n14) );
  XNOR2_X1 SBOX_s4_mul2_0_0_U5 ( .A(SBOX_s4_mul2_0_0_n11), .B(
        SBOX_s4_mul2_0_0_n14), .ZN(SBOX_s4_concat[3]) );
  NAND2_X1 SBOX_s4_mul2_0_0_U4 ( .A1(SBOX_stage3Out[5]), .A2(
        SBOX_s4_inv_out_0__1_), .ZN(SBOX_s4_mul2_0_0_n11) );
  NAND2_X1 SBOX_s4_mul2_0_0_U3 ( .A1(SBOX_s4_inv_out_0__0_), .A2(
        SBOX_stage3Out[4]), .ZN(SBOX_s4_mul2_0_0_n13) );
  XNOR2_X1 SBOX_s4_mul2_0_0_U2 ( .A(SBOX_s4_mul2_0_0_n14), .B(
        SBOX_s4_mul2_0_0_n13), .ZN(SBOX_s4_concat[2]) );
  OAI22_X1 SBOX_s4_mul2_0_0_U1 ( .A1(SBOX_s4_inv_out_0__0_), .A2(
        SBOX_s4_inv_out_0__1_), .B1(SBOX_stage3Out[4]), .B2(SBOX_stage3Out[5]), 
        .ZN(SBOX_s4_mul2_0_0_n12) );
  XOR2_X2 SBOX_s4_compr_0_0_U4 ( .A(SBOX_s4_regOut_0__1__2_), .B(
        SBOX_s4_regOut_0__2__2_), .Z(SBOX_stage4Out[6]) );
  XOR2_X2 SBOX_s4_compr_0_0_U3 ( .A(SBOX_s4_regOut_0__1__1_), .B(
        SBOX_s4_regOut_0__2__1_), .Z(SBOX_stage4Out[5]) );
  XOR2_X2 SBOX_s4_compr_0_0_U2 ( .A(SBOX_s4_regOut_0__1__3_), .B(
        SBOX_s4_regOut_0__2__3_), .Z(SBOX_stage4Out[7]) );
  XOR2_X2 SBOX_s4_compr_0_0_U1 ( .A(SBOX_s4_regOut_0__1__0_), .B(
        SBOX_s4_regOut_0__2__0_), .Z(SBOX_stage4Out[4]) );
  XOR2_X2 SBOX_s4_compr_1_0_U4 ( .A(SBOX_s4_regOut_1__1__2_), .B(
        SBOX_s4_regOut_1__2__2_), .Z(SBOX_stage4Out[18]) );
  XOR2_X2 SBOX_s4_compr_1_0_U3 ( .A(SBOX_s4_regOut_1__1__1_), .B(
        SBOX_s4_regOut_1__2__1_), .Z(SBOX_stage4Out[17]) );
  XOR2_X2 SBOX_s4_compr_1_0_U2 ( .A(SBOX_s4_regOut_1__1__3_), .B(
        SBOX_s4_regOut_1__2__3_), .Z(SBOX_stage4Out[19]) );
  XOR2_X2 SBOX_s4_compr_1_0_U1 ( .A(SBOX_s4_regOut_1__1__0_), .B(
        SBOX_s4_regOut_1__2__0_), .Z(SBOX_stage4Out[16]) );
  XNOR2_X1 SBOX_s5_U50 ( .A(SBOX_s5_n15), .B(SBOX_s5_n16), .ZN(
        SBOX_s5_refreshed[31]) );
  XNOR2_X1 SBOX_s5_U49 ( .A(randomS5[7]), .B(randomS5[15]), .ZN(SBOX_s5_n16)
         );
  XOR2_X1 SBOX_s5_U48 ( .A(randomS5[23]), .B(SBOX_s5_concat[31]), .Z(
        SBOX_s5_n15) );
  XOR2_X1 SBOX_s5_U47 ( .A(randomS5[19]), .B(SBOX_s5_concat[19]), .Z(
        SBOX_s5_refreshed[19]) );
  XNOR2_X1 SBOX_s5_U46 ( .A(SBOX_s5_n13), .B(SBOX_s5_n14), .ZN(
        SBOX_s5_refreshed[30]) );
  XNOR2_X1 SBOX_s5_U45 ( .A(randomS5[6]), .B(randomS5[14]), .ZN(SBOX_s5_n14)
         );
  XOR2_X1 SBOX_s5_U44 ( .A(randomS5[22]), .B(SBOX_s5_concat[30]), .Z(
        SBOX_s5_n13) );
  XNOR2_X1 SBOX_s5_U43 ( .A(SBOX_s5_n11), .B(SBOX_s5_n12), .ZN(
        SBOX_s5_refreshed[29]) );
  XNOR2_X1 SBOX_s5_U42 ( .A(randomS5[5]), .B(randomS5[13]), .ZN(SBOX_s5_n12)
         );
  XOR2_X1 SBOX_s5_U41 ( .A(randomS5[21]), .B(SBOX_s5_concat[29]), .Z(
        SBOX_s5_n11) );
  XOR2_X1 SBOX_s5_U40 ( .A(randomS5[17]), .B(SBOX_s5_concat[17]), .Z(
        SBOX_s5_refreshed[17]) );
  XOR2_X1 SBOX_s5_U39 ( .A(randomS5[7]), .B(SBOX_s5_concat[7]), .Z(
        SBOX_s5_refreshed[7]) );
  XNOR2_X1 SBOX_s5_U38 ( .A(SBOX_s5_n9), .B(SBOX_s5_n10), .ZN(
        SBOX_s5_refreshed[28]) );
  XNOR2_X1 SBOX_s5_U37 ( .A(randomS5[4]), .B(randomS5[12]), .ZN(SBOX_s5_n10)
         );
  XOR2_X1 SBOX_s5_U36 ( .A(randomS5[20]), .B(SBOX_s5_concat[28]), .Z(
        SBOX_s5_n9) );
  XNOR2_X1 SBOX_s5_U35 ( .A(SBOX_s5_n7), .B(SBOX_s5_n8), .ZN(
        SBOX_s5_refreshed[27]) );
  XNOR2_X1 SBOX_s5_U34 ( .A(randomS5[3]), .B(randomS5[11]), .ZN(SBOX_s5_n8) );
  XOR2_X1 SBOX_s5_U33 ( .A(randomS5[19]), .B(SBOX_s5_concat[27]), .Z(
        SBOX_s5_n7) );
  XOR2_X1 SBOX_s5_U32 ( .A(randomS5[16]), .B(SBOX_s5_concat[16]), .Z(
        SBOX_s5_refreshed[16]) );
  XOR2_X1 SBOX_s5_U31 ( .A(randomS5[15]), .B(SBOX_s5_concat[15]), .Z(
        SBOX_s5_refreshed[15]) );
  XNOR2_X1 SBOX_s5_U30 ( .A(SBOX_s5_n5), .B(SBOX_s5_n6), .ZN(
        SBOX_s5_refreshed[26]) );
  XNOR2_X1 SBOX_s5_U29 ( .A(randomS5[2]), .B(randomS5[10]), .ZN(SBOX_s5_n6) );
  XOR2_X1 SBOX_s5_U28 ( .A(randomS5[18]), .B(SBOX_s5_concat[26]), .Z(
        SBOX_s5_n5) );
  XOR2_X1 SBOX_s5_U27 ( .A(randomS5[20]), .B(SBOX_s5_concat[20]), .Z(
        SBOX_s5_refreshed[20]) );
  XOR2_X1 SBOX_s5_U26 ( .A(randomS5[14]), .B(SBOX_s5_concat[14]), .Z(
        SBOX_s5_refreshed[14]) );
  XOR2_X1 SBOX_s5_U25 ( .A(randomS5[13]), .B(SBOX_s5_concat[13]), .Z(
        SBOX_s5_refreshed[13]) );
  XNOR2_X1 SBOX_s5_U24 ( .A(SBOX_s5_n3), .B(SBOX_s5_n4), .ZN(
        SBOX_s5_refreshed[25]) );
  XNOR2_X1 SBOX_s5_U23 ( .A(randomS5[1]), .B(randomS5[9]), .ZN(SBOX_s5_n4) );
  XOR2_X1 SBOX_s5_U22 ( .A(randomS5[17]), .B(SBOX_s5_concat[25]), .Z(
        SBOX_s5_n3) );
  XOR2_X1 SBOX_s5_U21 ( .A(randomS5[23]), .B(SBOX_s5_concat[23]), .Z(
        SBOX_s5_refreshed[23]) );
  XOR2_X1 SBOX_s5_U20 ( .A(randomS5[18]), .B(SBOX_s5_concat[18]), .Z(
        SBOX_s5_refreshed[18]) );
  XOR2_X1 SBOX_s5_U19 ( .A(randomS5[12]), .B(SBOX_s5_concat[12]), .Z(
        SBOX_s5_refreshed[12]) );
  XNOR2_X1 SBOX_s5_U18 ( .A(SBOX_s5_n1), .B(SBOX_s5_n2), .ZN(
        SBOX_s5_refreshed[24]) );
  XNOR2_X1 SBOX_s5_U17 ( .A(randomS5[0]), .B(randomS5[8]), .ZN(SBOX_s5_n2) );
  XOR2_X1 SBOX_s5_U16 ( .A(randomS5[16]), .B(SBOX_s5_concat[24]), .Z(
        SBOX_s5_n1) );
  XOR2_X1 SBOX_s5_U15 ( .A(randomS5[22]), .B(SBOX_s5_concat[22]), .Z(
        SBOX_s5_refreshed[22]) );
  XOR2_X1 SBOX_s5_U14 ( .A(randomS5[5]), .B(SBOX_s5_concat[5]), .Z(
        SBOX_s5_refreshed[5]) );
  XOR2_X1 SBOX_s5_U13 ( .A(randomS5[3]), .B(SBOX_s5_concat[3]), .Z(
        SBOX_s5_refreshed[3]) );
  XOR2_X1 SBOX_s5_U12 ( .A(randomS5[10]), .B(SBOX_s5_concat[10]), .Z(
        SBOX_s5_refreshed[10]) );
  XOR2_X1 SBOX_s5_U11 ( .A(randomS5[6]), .B(SBOX_s5_concat[6]), .Z(
        SBOX_s5_refreshed[6]) );
  XOR2_X1 SBOX_s5_U10 ( .A(randomS5[1]), .B(SBOX_s5_concat[1]), .Z(
        SBOX_s5_refreshed[1]) );
  XOR2_X1 SBOX_s5_U9 ( .A(randomS5[21]), .B(SBOX_s5_concat[21]), .Z(
        SBOX_s5_refreshed[21]) );
  XOR2_X1 SBOX_s5_U8 ( .A(randomS5[11]), .B(SBOX_s5_concat[11]), .Z(
        SBOX_s5_refreshed[11]) );
  XOR2_X1 SBOX_s5_U7 ( .A(randomS5[0]), .B(SBOX_s5_concat[0]), .Z(
        SBOX_s5_refreshed[0]) );
  XOR2_X1 SBOX_s5_U6 ( .A(randomS5[9]), .B(SBOX_s5_concat[9]), .Z(
        SBOX_s5_refreshed[9]) );
  XOR2_X1 SBOX_s5_U5 ( .A(randomS5[4]), .B(SBOX_s5_concat[4]), .Z(
        SBOX_s5_refreshed[4]) );
  XOR2_X1 SBOX_s5_U4 ( .A(randomS5[2]), .B(SBOX_s5_concat[2]), .Z(
        SBOX_s5_refreshed[2]) );
  XOR2_X1 SBOX_s5_U3 ( .A(randomS5[8]), .B(SBOX_s5_concat[8]), .Z(
        SBOX_s5_refreshed[8]) );
  DFF_X1 SBOX_s5_regOut_reg_0__0__0_ ( .D(SBOX_s5_refreshed[0]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[0]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__0__1_ ( .D(SBOX_s5_refreshed[1]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[1]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__0__2_ ( .D(SBOX_s5_refreshed[2]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[2]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__0__3_ ( .D(SBOX_s5_refreshed[3]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[3]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__0__4_ ( .D(SBOX_s5_refreshed[4]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[4]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__0__5_ ( .D(SBOX_s5_refreshed[5]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[5]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__0__6_ ( .D(SBOX_s5_refreshed[6]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[6]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__0__7_ ( .D(SBOX_s5_refreshed[7]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[7]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__1__0_ ( .D(SBOX_s5_refreshed[8]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[8]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__1__1_ ( .D(SBOX_s5_refreshed[9]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[9]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__1__2_ ( .D(SBOX_s5_refreshed[10]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[10]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__1__3_ ( .D(SBOX_s5_refreshed[11]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[11]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__1__4_ ( .D(SBOX_s5_refreshed[12]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[12]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__1__5_ ( .D(SBOX_s5_refreshed[13]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[13]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__1__6_ ( .D(SBOX_s5_refreshed[14]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[14]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_0__1__7_ ( .D(SBOX_s5_refreshed[15]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[15]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__0__0_ ( .D(SBOX_s5_refreshed[16]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[16]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__0__1_ ( .D(SBOX_s5_refreshed[17]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[17]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__0__2_ ( .D(SBOX_s5_refreshed[18]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[18]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__0__3_ ( .D(SBOX_s5_refreshed[19]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[19]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__0__4_ ( .D(SBOX_s5_refreshed[20]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[20]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__0__5_ ( .D(SBOX_s5_refreshed[21]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[21]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__0__6_ ( .D(SBOX_s5_refreshed[22]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[22]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__0__7_ ( .D(SBOX_s5_refreshed[23]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[23]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__1__0_ ( .D(SBOX_s5_refreshed[24]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[24]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__1__1_ ( .D(SBOX_s5_refreshed[25]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[25]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__1__2_ ( .D(SBOX_s5_refreshed[26]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[26]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__1__3_ ( .D(SBOX_s5_refreshed[27]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[27]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__1__4_ ( .D(SBOX_s5_refreshed[28]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[28]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__1__5_ ( .D(SBOX_s5_refreshed[29]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[29]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__1__6_ ( .D(SBOX_s5_refreshed[30]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[30]), .QN() );
  DFF_X1 SBOX_s5_regOut_reg_1__1__7_ ( .D(SBOX_s5_refreshed[31]), .CK(ClkxCI), 
        .Q(SBOX_s5_regOut[31]), .QN() );
  AOI221_X1 SBOX_s5_mul1_1_1_U28 ( .B1(SBOX_stage4Out[18]), .B2(
        SBOX_stage4Out[19]), .C1(SBOX_stage4Out[22]), .C2(SBOX_stage4Out[23]), 
        .A(SBOX_s5_mul1_1_1_n73), .ZN(SBOX_s5_mul1_1_1_n75) );
  OAI22_X1 SBOX_s5_mul1_1_1_U27 ( .A1(SBOX_stage4Out[18]), .A2(
        SBOX_stage4Out[19]), .B1(SBOX_stage4Out[23]), .B2(SBOX_stage4Out[22]), 
        .ZN(SBOX_s5_mul1_1_1_n73) );
  XNOR2_X1 SBOX_s5_mul1_1_1_U26 ( .A(SBOX_s5_mul1_1_1_n63), .B(
        SBOX_s5_mul1_1_1_n62), .ZN(SBOX_s5_mul1_1_1_n74) );
  XOR2_X1 SBOX_s5_mul1_1_1_U25 ( .A(SBOX_stage4Out[17]), .B(SBOX_stage4Out[19]), .Z(SBOX_s5_mul1_1_1_n64) );
  XNOR2_X1 SBOX_s5_mul1_1_1_U24 ( .A(SBOX_stage4Out[16]), .B(
        SBOX_stage4Out[18]), .ZN(SBOX_s5_mul1_1_1_n69) );
  AOI221_X1 SBOX_s5_mul1_1_1_U23 ( .B1(SBOX_stage4Out[16]), .B2(
        SBOX_stage4Out[17]), .C1(SBOX_stage4Out[20]), .C2(SBOX_stage4Out[21]), 
        .A(SBOX_s5_mul1_1_1_n61), .ZN(SBOX_s5_mul1_1_1_n72) );
  OAI22_X1 SBOX_s5_mul1_1_1_U22 ( .A1(SBOX_stage4Out[16]), .A2(
        SBOX_stage4Out[17]), .B1(SBOX_stage4Out[21]), .B2(SBOX_stage4Out[20]), 
        .ZN(SBOX_s5_mul1_1_1_n61) );
  XNOR2_X1 SBOX_s5_mul1_1_1_U21 ( .A(SBOX_s5_mul1_1_1_n59), .B(
        SBOX_s5_mul1_1_1_n60), .ZN(SBOX_s5_concat[27]) );
  XOR2_X1 SBOX_s5_mul1_1_1_U20 ( .A(SBOX_s5_mul1_1_1_n76), .B(
        SBOX_s5_mul1_1_1_n75), .Z(SBOX_s5_mul1_1_1_n60) );
  NAND2_X1 SBOX_s5_mul1_1_1_U19 ( .A1(SBOX_stage4Out[19]), .A2(
        SBOX_stage4Out[23]), .ZN(SBOX_s5_mul1_1_1_n59) );
  XNOR2_X1 SBOX_s5_mul1_1_1_U18 ( .A(SBOX_s5_mul1_1_1_n57), .B(
        SBOX_s5_mul1_1_1_n58), .ZN(SBOX_s5_concat[26]) );
  XOR2_X1 SBOX_s5_mul1_1_1_U17 ( .A(SBOX_s5_mul1_1_1_n74), .B(
        SBOX_s5_mul1_1_1_n75), .Z(SBOX_s5_mul1_1_1_n58) );
  NAND2_X1 SBOX_s5_mul1_1_1_U16 ( .A1(SBOX_stage4Out[18]), .A2(
        SBOX_stage4Out[22]), .ZN(SBOX_s5_mul1_1_1_n57) );
  XNOR2_X1 SBOX_s5_mul1_1_1_U15 ( .A(SBOX_s5_mul1_1_1_n55), .B(
        SBOX_s5_mul1_1_1_n56), .ZN(SBOX_s5_concat[25]) );
  XOR2_X1 SBOX_s5_mul1_1_1_U14 ( .A(SBOX_s5_mul1_1_1_n76), .B(
        SBOX_s5_mul1_1_1_n72), .Z(SBOX_s5_mul1_1_1_n56) );
  NAND2_X1 SBOX_s5_mul1_1_1_U13 ( .A1(SBOX_stage4Out[17]), .A2(
        SBOX_stage4Out[21]), .ZN(SBOX_s5_mul1_1_1_n55) );
  XNOR2_X1 SBOX_s5_mul1_1_1_U12 ( .A(SBOX_s5_mul1_1_1_n53), .B(
        SBOX_s5_mul1_1_1_n54), .ZN(SBOX_s5_concat[24]) );
  XOR2_X1 SBOX_s5_mul1_1_1_U11 ( .A(SBOX_s5_mul1_1_1_n72), .B(
        SBOX_s5_mul1_1_1_n74), .Z(SBOX_s5_mul1_1_1_n54) );
  NAND2_X1 SBOX_s5_mul1_1_1_U10 ( .A1(SBOX_stage4Out[16]), .A2(
        SBOX_stage4Out[20]), .ZN(SBOX_s5_mul1_1_1_n53) );
  NAND2_X1 SBOX_s5_mul1_1_1_U9 ( .A1(SBOX_s5_mul1_1_1_n67), .A2(
        SBOX_s5_mul1_1_1_n69), .ZN(SBOX_s5_mul1_1_1_n65) );
  INV_X1 SBOX_s5_mul1_1_1_U8 ( .A(SBOX_s5_mul1_1_1_n64), .ZN(
        SBOX_s5_mul1_1_1_n71) );
  NAND2_X1 SBOX_s5_mul1_1_1_U7 ( .A1(SBOX_s5_mul1_1_1_n67), .A2(
        SBOX_s5_mul1_1_1_n71), .ZN(SBOX_s5_mul1_1_1_n68) );
  XNOR2_X1 SBOX_s5_mul1_1_1_U6 ( .A(SBOX_s5_mul1_1_1_n66), .B(
        SBOX_s5_mul1_1_1_n65), .ZN(SBOX_s5_mul1_1_1_n70) );
  OAI22_X1 SBOX_s5_mul1_1_1_U5 ( .A1(SBOX_s5_mul1_1_1_n71), .A2(
        SBOX_s5_mul1_1_1_n70), .B1(SBOX_s5_mul1_1_1_n69), .B2(
        SBOX_s5_mul1_1_1_n68), .ZN(SBOX_s5_mul1_1_1_n76) );
  NAND2_X1 SBOX_s5_mul1_1_1_U4 ( .A1(SBOX_s5_mul1_1_1_n67), .A2(
        SBOX_s5_mul1_1_1_n64), .ZN(SBOX_s5_mul1_1_1_n62) );
  NOR2_X1 SBOX_s5_mul1_1_1_U3 ( .A1(SBOX_s5_mul1_1_1_n69), .A2(
        SBOX_s5_mul1_1_1_n66), .ZN(SBOX_s5_mul1_1_1_n63) );
  XNOR2_X1 SBOX_s5_mul1_1_1_U2 ( .A(SBOX_stage4Out[20]), .B(SBOX_stage4Out[22]), .ZN(SBOX_s5_mul1_1_1_n66) );
  XOR2_X1 SBOX_s5_mul1_1_1_U1 ( .A(SBOX_stage4Out[21]), .B(SBOX_stage4Out[23]), 
        .Z(SBOX_s5_mul1_1_1_n67) );
  AOI221_X1 SBOX_s5_mul1_1_0_U29 ( .B1(SBOX_stage4Out[6]), .B2(
        SBOX_stage4Out[7]), .C1(SBOX_stage4Out[22]), .C2(SBOX_stage4Out[23]), 
        .A(SBOX_s5_mul1_1_0_n74), .ZN(SBOX_s5_mul1_1_0_n76) );
  OAI22_X1 SBOX_s5_mul1_1_0_U28 ( .A1(SBOX_stage4Out[6]), .A2(
        SBOX_stage4Out[7]), .B1(SBOX_stage4Out[23]), .B2(SBOX_stage4Out[22]), 
        .ZN(SBOX_s5_mul1_1_0_n74) );
  XOR2_X1 SBOX_s5_mul1_1_0_U27 ( .A(SBOX_stage4Out[5]), .B(SBOX_stage4Out[7]), 
        .Z(SBOX_s5_mul1_1_0_n69) );
  XNOR2_X1 SBOX_s5_mul1_1_0_U26 ( .A(SBOX_stage4Out[4]), .B(SBOX_stage4Out[6]), 
        .ZN(SBOX_s5_mul1_1_0_n72) );
  AOI221_X1 SBOX_s5_mul1_1_0_U25 ( .B1(SBOX_stage4Out[4]), .B2(
        SBOX_stage4Out[5]), .C1(SBOX_stage4Out[20]), .C2(SBOX_stage4Out[21]), 
        .A(SBOX_s5_mul1_1_0_n68), .ZN(SBOX_s5_mul1_1_0_n73) );
  OAI22_X1 SBOX_s5_mul1_1_0_U24 ( .A1(SBOX_stage4Out[4]), .A2(
        SBOX_stage4Out[5]), .B1(SBOX_stage4Out[21]), .B2(SBOX_stage4Out[20]), 
        .ZN(SBOX_s5_mul1_1_0_n68) );
  XNOR2_X1 SBOX_s5_mul1_1_0_U23 ( .A(SBOX_s5_mul1_1_0_n66), .B(
        SBOX_s5_mul1_1_0_n67), .ZN(SBOX_s5_concat[19]) );
  XOR2_X1 SBOX_s5_mul1_1_0_U22 ( .A(SBOX_s5_mul1_1_0_n77), .B(
        SBOX_s5_mul1_1_0_n76), .Z(SBOX_s5_mul1_1_0_n67) );
  NAND2_X1 SBOX_s5_mul1_1_0_U21 ( .A1(SBOX_stage4Out[7]), .A2(
        SBOX_stage4Out[23]), .ZN(SBOX_s5_mul1_1_0_n66) );
  XNOR2_X1 SBOX_s5_mul1_1_0_U20 ( .A(SBOX_s5_mul1_1_0_n64), .B(
        SBOX_s5_mul1_1_0_n65), .ZN(SBOX_s5_concat[17]) );
  XOR2_X1 SBOX_s5_mul1_1_0_U19 ( .A(SBOX_s5_mul1_1_0_n77), .B(
        SBOX_s5_mul1_1_0_n73), .Z(SBOX_s5_mul1_1_0_n65) );
  NAND2_X1 SBOX_s5_mul1_1_0_U18 ( .A1(SBOX_stage4Out[5]), .A2(
        SBOX_stage4Out[21]), .ZN(SBOX_s5_mul1_1_0_n64) );
  XNOR2_X1 SBOX_s5_mul1_1_0_U17 ( .A(SBOX_s5_mul1_1_0_n62), .B(
        SBOX_s5_mul1_1_0_n63), .ZN(SBOX_s5_concat[16]) );
  XOR2_X1 SBOX_s5_mul1_1_0_U16 ( .A(SBOX_s5_mul1_1_0_n75), .B(
        SBOX_s5_mul1_1_0_n73), .Z(SBOX_s5_mul1_1_0_n63) );
  NAND2_X1 SBOX_s5_mul1_1_0_U15 ( .A1(SBOX_stage4Out[4]), .A2(
        SBOX_stage4Out[20]), .ZN(SBOX_s5_mul1_1_0_n62) );
  XNOR2_X1 SBOX_s5_mul1_1_0_U14 ( .A(SBOX_s5_mul1_1_0_n60), .B(
        SBOX_s5_mul1_1_0_n61), .ZN(SBOX_s5_concat[18]) );
  XOR2_X1 SBOX_s5_mul1_1_0_U13 ( .A(SBOX_s5_mul1_1_0_n76), .B(
        SBOX_s5_mul1_1_0_n75), .Z(SBOX_s5_mul1_1_0_n61) );
  NAND2_X1 SBOX_s5_mul1_1_0_U12 ( .A1(SBOX_stage4Out[6]), .A2(
        SBOX_stage4Out[22]), .ZN(SBOX_s5_mul1_1_0_n60) );
  INV_X1 SBOX_s5_mul1_1_0_U11 ( .A(SBOX_s5_mul1_1_0_n71), .ZN(
        SBOX_s5_mul1_1_0_n59) );
  INV_X1 SBOX_s5_mul1_1_0_U10 ( .A(SBOX_s5_mul1_1_0_n69), .ZN(
        SBOX_s5_mul1_1_0_n58) );
  XNOR2_X1 SBOX_s5_mul1_1_0_U9 ( .A(SBOX_s5_mul1_1_0_n56), .B(
        SBOX_s5_mul1_1_0_n70), .ZN(SBOX_s5_mul1_1_0_n57) );
  NAND2_X1 SBOX_s5_mul1_1_0_U8 ( .A1(SBOX_s5_mul1_1_0_n71), .A2(
        SBOX_s5_mul1_1_0_n72), .ZN(SBOX_s5_mul1_1_0_n56) );
  XNOR2_X1 SBOX_s5_mul1_1_0_U6 ( .A(SBOX_s5_mul1_1_0_n53), .B(
        SBOX_s5_mul1_1_0_n54), .ZN(SBOX_s5_mul1_1_0_n75) );
  NAND2_X1 SBOX_s5_mul1_1_0_U5 ( .A1(SBOX_s5_mul1_1_0_n69), .A2(
        SBOX_s5_mul1_1_0_n71), .ZN(SBOX_s5_mul1_1_0_n54) );
  NOR2_X1 SBOX_s5_mul1_1_0_U4 ( .A1(SBOX_s5_mul1_1_0_n72), .A2(
        SBOX_s5_mul1_1_0_n70), .ZN(SBOX_s5_mul1_1_0_n53) );
  XNOR2_X1 SBOX_s5_mul1_1_0_U3 ( .A(SBOX_stage4Out[20]), .B(SBOX_stage4Out[22]), .ZN(SBOX_s5_mul1_1_0_n70) );
  XOR2_X1 SBOX_s5_mul1_1_0_U2 ( .A(SBOX_stage4Out[21]), .B(SBOX_stage4Out[23]), 
        .Z(SBOX_s5_mul1_1_0_n71) );
  OAI33_X1 SBOX_s5_mul1_1_0_U1 ( .A1(1'b0), .A2(SBOX_s5_mul1_1_0_n57), .A3(
        SBOX_s5_mul1_1_0_n58), .B1(SBOX_s5_mul1_1_0_n69), .B2(
        SBOX_s5_mul1_1_0_n72), .B3(SBOX_s5_mul1_1_0_n59), .ZN(
        SBOX_s5_mul1_1_0_n77) );
  AOI221_X1 SBOX_s5_mul1_0_1_U28 ( .B1(SBOX_stage4Out[18]), .B2(
        SBOX_stage4Out[19]), .C1(SBOX_stage4Out[10]), .C2(SBOX_stage4Out[11]), 
        .A(SBOX_s5_mul1_0_1_n73), .ZN(SBOX_s5_mul1_0_1_n75) );
  OAI22_X1 SBOX_s5_mul1_0_1_U27 ( .A1(SBOX_stage4Out[18]), .A2(
        SBOX_stage4Out[19]), .B1(SBOX_stage4Out[11]), .B2(SBOX_stage4Out[10]), 
        .ZN(SBOX_s5_mul1_0_1_n73) );
  XNOR2_X1 SBOX_s5_mul1_0_1_U26 ( .A(SBOX_s5_mul1_0_1_n63), .B(
        SBOX_s5_mul1_0_1_n62), .ZN(SBOX_s5_mul1_0_1_n74) );
  XOR2_X1 SBOX_s5_mul1_0_1_U25 ( .A(SBOX_stage4Out[17]), .B(SBOX_stage4Out[19]), .Z(SBOX_s5_mul1_0_1_n64) );
  XNOR2_X1 SBOX_s5_mul1_0_1_U24 ( .A(SBOX_stage4Out[16]), .B(
        SBOX_stage4Out[18]), .ZN(SBOX_s5_mul1_0_1_n69) );
  AOI221_X1 SBOX_s5_mul1_0_1_U23 ( .B1(SBOX_stage4Out[16]), .B2(
        SBOX_stage4Out[17]), .C1(SBOX_stage4Out[8]), .C2(SBOX_stage4Out[9]), 
        .A(SBOX_s5_mul1_0_1_n61), .ZN(SBOX_s5_mul1_0_1_n72) );
  OAI22_X1 SBOX_s5_mul1_0_1_U22 ( .A1(SBOX_stage4Out[16]), .A2(
        SBOX_stage4Out[17]), .B1(SBOX_stage4Out[9]), .B2(SBOX_stage4Out[8]), 
        .ZN(SBOX_s5_mul1_0_1_n61) );
  XNOR2_X1 SBOX_s5_mul1_0_1_U21 ( .A(SBOX_s5_mul1_0_1_n59), .B(
        SBOX_s5_mul1_0_1_n60), .ZN(SBOX_s5_concat[10]) );
  XOR2_X1 SBOX_s5_mul1_0_1_U20 ( .A(SBOX_s5_mul1_0_1_n74), .B(
        SBOX_s5_mul1_0_1_n75), .Z(SBOX_s5_mul1_0_1_n60) );
  NAND2_X1 SBOX_s5_mul1_0_1_U19 ( .A1(SBOX_stage4Out[18]), .A2(
        SBOX_stage4Out[10]), .ZN(SBOX_s5_mul1_0_1_n59) );
  XNOR2_X1 SBOX_s5_mul1_0_1_U18 ( .A(SBOX_s5_mul1_0_1_n57), .B(
        SBOX_s5_mul1_0_1_n58), .ZN(SBOX_s5_concat[11]) );
  XOR2_X1 SBOX_s5_mul1_0_1_U17 ( .A(SBOX_s5_mul1_0_1_n76), .B(
        SBOX_s5_mul1_0_1_n75), .Z(SBOX_s5_mul1_0_1_n58) );
  NAND2_X1 SBOX_s5_mul1_0_1_U16 ( .A1(SBOX_stage4Out[19]), .A2(
        SBOX_stage4Out[11]), .ZN(SBOX_s5_mul1_0_1_n57) );
  XNOR2_X1 SBOX_s5_mul1_0_1_U15 ( .A(SBOX_s5_mul1_0_1_n55), .B(
        SBOX_s5_mul1_0_1_n56), .ZN(SBOX_s5_concat[9]) );
  XOR2_X1 SBOX_s5_mul1_0_1_U14 ( .A(SBOX_s5_mul1_0_1_n76), .B(
        SBOX_s5_mul1_0_1_n72), .Z(SBOX_s5_mul1_0_1_n56) );
  NAND2_X1 SBOX_s5_mul1_0_1_U13 ( .A1(SBOX_stage4Out[17]), .A2(
        SBOX_stage4Out[9]), .ZN(SBOX_s5_mul1_0_1_n55) );
  XNOR2_X1 SBOX_s5_mul1_0_1_U12 ( .A(SBOX_s5_mul1_0_1_n53), .B(
        SBOX_s5_mul1_0_1_n54), .ZN(SBOX_s5_concat[8]) );
  XOR2_X1 SBOX_s5_mul1_0_1_U11 ( .A(SBOX_s5_mul1_0_1_n72), .B(
        SBOX_s5_mul1_0_1_n74), .Z(SBOX_s5_mul1_0_1_n54) );
  NAND2_X1 SBOX_s5_mul1_0_1_U10 ( .A1(SBOX_stage4Out[16]), .A2(
        SBOX_stage4Out[8]), .ZN(SBOX_s5_mul1_0_1_n53) );
  NAND2_X1 SBOX_s5_mul1_0_1_U9 ( .A1(SBOX_s5_mul1_0_1_n67), .A2(
        SBOX_s5_mul1_0_1_n69), .ZN(SBOX_s5_mul1_0_1_n65) );
  INV_X1 SBOX_s5_mul1_0_1_U8 ( .A(SBOX_s5_mul1_0_1_n64), .ZN(
        SBOX_s5_mul1_0_1_n71) );
  NAND2_X1 SBOX_s5_mul1_0_1_U7 ( .A1(SBOX_s5_mul1_0_1_n67), .A2(
        SBOX_s5_mul1_0_1_n71), .ZN(SBOX_s5_mul1_0_1_n68) );
  XNOR2_X1 SBOX_s5_mul1_0_1_U6 ( .A(SBOX_s5_mul1_0_1_n66), .B(
        SBOX_s5_mul1_0_1_n65), .ZN(SBOX_s5_mul1_0_1_n70) );
  OAI22_X1 SBOX_s5_mul1_0_1_U5 ( .A1(SBOX_s5_mul1_0_1_n71), .A2(
        SBOX_s5_mul1_0_1_n70), .B1(SBOX_s5_mul1_0_1_n69), .B2(
        SBOX_s5_mul1_0_1_n68), .ZN(SBOX_s5_mul1_0_1_n76) );
  NAND2_X1 SBOX_s5_mul1_0_1_U4 ( .A1(SBOX_s5_mul1_0_1_n67), .A2(
        SBOX_s5_mul1_0_1_n64), .ZN(SBOX_s5_mul1_0_1_n62) );
  NOR2_X1 SBOX_s5_mul1_0_1_U3 ( .A1(SBOX_s5_mul1_0_1_n69), .A2(
        SBOX_s5_mul1_0_1_n66), .ZN(SBOX_s5_mul1_0_1_n63) );
  XNOR2_X1 SBOX_s5_mul1_0_1_U2 ( .A(SBOX_stage4Out[8]), .B(SBOX_stage4Out[10]), 
        .ZN(SBOX_s5_mul1_0_1_n66) );
  XOR2_X1 SBOX_s5_mul1_0_1_U1 ( .A(SBOX_stage4Out[9]), .B(SBOX_stage4Out[11]), 
        .Z(SBOX_s5_mul1_0_1_n67) );
  AOI221_X1 SBOX_s5_mul1_0_0_U28 ( .B1(SBOX_stage4Out[6]), .B2(
        SBOX_stage4Out[7]), .C1(SBOX_stage4Out[10]), .C2(SBOX_stage4Out[11]), 
        .A(SBOX_s5_mul1_0_0_n73), .ZN(SBOX_s5_mul1_0_0_n75) );
  OAI22_X1 SBOX_s5_mul1_0_0_U27 ( .A1(SBOX_stage4Out[6]), .A2(
        SBOX_stage4Out[7]), .B1(SBOX_stage4Out[11]), .B2(SBOX_stage4Out[10]), 
        .ZN(SBOX_s5_mul1_0_0_n73) );
  XNOR2_X1 SBOX_s5_mul1_0_0_U26 ( .A(SBOX_s5_mul1_0_0_n63), .B(
        SBOX_s5_mul1_0_0_n62), .ZN(SBOX_s5_mul1_0_0_n74) );
  XOR2_X1 SBOX_s5_mul1_0_0_U25 ( .A(SBOX_stage4Out[5]), .B(SBOX_stage4Out[7]), 
        .Z(SBOX_s5_mul1_0_0_n64) );
  XNOR2_X1 SBOX_s5_mul1_0_0_U24 ( .A(SBOX_stage4Out[4]), .B(SBOX_stage4Out[6]), 
        .ZN(SBOX_s5_mul1_0_0_n69) );
  AOI221_X1 SBOX_s5_mul1_0_0_U23 ( .B1(SBOX_stage4Out[4]), .B2(
        SBOX_stage4Out[5]), .C1(SBOX_stage4Out[8]), .C2(SBOX_stage4Out[9]), 
        .A(SBOX_s5_mul1_0_0_n61), .ZN(SBOX_s5_mul1_0_0_n72) );
  OAI22_X1 SBOX_s5_mul1_0_0_U22 ( .A1(SBOX_stage4Out[4]), .A2(
        SBOX_stage4Out[5]), .B1(SBOX_stage4Out[9]), .B2(SBOX_stage4Out[8]), 
        .ZN(SBOX_s5_mul1_0_0_n61) );
  XNOR2_X1 SBOX_s5_mul1_0_0_U21 ( .A(SBOX_s5_mul1_0_0_n59), .B(
        SBOX_s5_mul1_0_0_n60), .ZN(SBOX_s5_concat[3]) );
  XOR2_X1 SBOX_s5_mul1_0_0_U20 ( .A(SBOX_s5_mul1_0_0_n76), .B(
        SBOX_s5_mul1_0_0_n75), .Z(SBOX_s5_mul1_0_0_n60) );
  NAND2_X1 SBOX_s5_mul1_0_0_U19 ( .A1(SBOX_stage4Out[7]), .A2(
        SBOX_stage4Out[11]), .ZN(SBOX_s5_mul1_0_0_n59) );
  XNOR2_X1 SBOX_s5_mul1_0_0_U18 ( .A(SBOX_s5_mul1_0_0_n57), .B(
        SBOX_s5_mul1_0_0_n58), .ZN(SBOX_s5_concat[1]) );
  XOR2_X1 SBOX_s5_mul1_0_0_U17 ( .A(SBOX_s5_mul1_0_0_n76), .B(
        SBOX_s5_mul1_0_0_n72), .Z(SBOX_s5_mul1_0_0_n58) );
  NAND2_X1 SBOX_s5_mul1_0_0_U16 ( .A1(SBOX_stage4Out[5]), .A2(
        SBOX_stage4Out[9]), .ZN(SBOX_s5_mul1_0_0_n57) );
  XNOR2_X1 SBOX_s5_mul1_0_0_U15 ( .A(SBOX_s5_mul1_0_0_n55), .B(
        SBOX_s5_mul1_0_0_n56), .ZN(SBOX_s5_concat[0]) );
  XOR2_X1 SBOX_s5_mul1_0_0_U14 ( .A(SBOX_s5_mul1_0_0_n74), .B(
        SBOX_s5_mul1_0_0_n72), .Z(SBOX_s5_mul1_0_0_n56) );
  NAND2_X1 SBOX_s5_mul1_0_0_U13 ( .A1(SBOX_stage4Out[4]), .A2(
        SBOX_stage4Out[8]), .ZN(SBOX_s5_mul1_0_0_n55) );
  XNOR2_X1 SBOX_s5_mul1_0_0_U12 ( .A(SBOX_s5_mul1_0_0_n53), .B(
        SBOX_s5_mul1_0_0_n54), .ZN(SBOX_s5_concat[2]) );
  XOR2_X1 SBOX_s5_mul1_0_0_U11 ( .A(SBOX_s5_mul1_0_0_n75), .B(
        SBOX_s5_mul1_0_0_n74), .Z(SBOX_s5_mul1_0_0_n54) );
  NAND2_X1 SBOX_s5_mul1_0_0_U10 ( .A1(SBOX_stage4Out[6]), .A2(
        SBOX_stage4Out[10]), .ZN(SBOX_s5_mul1_0_0_n53) );
  NAND2_X1 SBOX_s5_mul1_0_0_U9 ( .A1(SBOX_s5_mul1_0_0_n67), .A2(
        SBOX_s5_mul1_0_0_n69), .ZN(SBOX_s5_mul1_0_0_n65) );
  INV_X1 SBOX_s5_mul1_0_0_U8 ( .A(SBOX_s5_mul1_0_0_n64), .ZN(
        SBOX_s5_mul1_0_0_n71) );
  NAND2_X1 SBOX_s5_mul1_0_0_U7 ( .A1(SBOX_s5_mul1_0_0_n67), .A2(
        SBOX_s5_mul1_0_0_n71), .ZN(SBOX_s5_mul1_0_0_n68) );
  XNOR2_X1 SBOX_s5_mul1_0_0_U6 ( .A(SBOX_s5_mul1_0_0_n66), .B(
        SBOX_s5_mul1_0_0_n65), .ZN(SBOX_s5_mul1_0_0_n70) );
  OAI22_X1 SBOX_s5_mul1_0_0_U5 ( .A1(SBOX_s5_mul1_0_0_n71), .A2(
        SBOX_s5_mul1_0_0_n70), .B1(SBOX_s5_mul1_0_0_n69), .B2(
        SBOX_s5_mul1_0_0_n68), .ZN(SBOX_s5_mul1_0_0_n76) );
  NAND2_X1 SBOX_s5_mul1_0_0_U4 ( .A1(SBOX_s5_mul1_0_0_n67), .A2(
        SBOX_s5_mul1_0_0_n64), .ZN(SBOX_s5_mul1_0_0_n62) );
  NOR2_X1 SBOX_s5_mul1_0_0_U3 ( .A1(SBOX_s5_mul1_0_0_n69), .A2(
        SBOX_s5_mul1_0_0_n66), .ZN(SBOX_s5_mul1_0_0_n63) );
  XNOR2_X1 SBOX_s5_mul1_0_0_U2 ( .A(SBOX_stage4Out[8]), .B(SBOX_stage4Out[10]), 
        .ZN(SBOX_s5_mul1_0_0_n66) );
  XOR2_X1 SBOX_s5_mul1_0_0_U1 ( .A(SBOX_stage4Out[9]), .B(SBOX_stage4Out[11]), 
        .Z(SBOX_s5_mul1_0_0_n67) );
  AOI221_X1 SBOX_s5_mul2_1_1_U29 ( .B1(SBOX_stage4Out[14]), .B2(
        SBOX_stage4Out[15]), .C1(SBOX_stage4Out[18]), .C2(SBOX_stage4Out[19]), 
        .A(SBOX_s5_mul2_1_1_n74), .ZN(SBOX_s5_mul2_1_1_n76) );
  OAI22_X1 SBOX_s5_mul2_1_1_U28 ( .A1(SBOX_stage4Out[14]), .A2(
        SBOX_stage4Out[15]), .B1(SBOX_stage4Out[19]), .B2(SBOX_stage4Out[18]), 
        .ZN(SBOX_s5_mul2_1_1_n74) );
  XNOR2_X1 SBOX_s5_mul2_1_1_U27 ( .A(SBOX_s5_mul2_1_1_n68), .B(
        SBOX_s5_mul2_1_1_n67), .ZN(SBOX_s5_mul2_1_1_n75) );
  XOR2_X1 SBOX_s5_mul2_1_1_U26 ( .A(SBOX_stage4Out[17]), .B(SBOX_stage4Out[19]), .Z(SBOX_s5_mul2_1_1_n71) );
  XNOR2_X1 SBOX_s5_mul2_1_1_U25 ( .A(SBOX_stage4Out[16]), .B(
        SBOX_stage4Out[18]), .ZN(SBOX_s5_mul2_1_1_n70) );
  AOI221_X1 SBOX_s5_mul2_1_1_U24 ( .B1(SBOX_stage4Out[12]), .B2(
        SBOX_stage4Out[13]), .C1(SBOX_stage4Out[16]), .C2(SBOX_stage4Out[17]), 
        .A(SBOX_s5_mul2_1_1_n66), .ZN(SBOX_s5_mul2_1_1_n73) );
  OAI22_X1 SBOX_s5_mul2_1_1_U23 ( .A1(SBOX_stage4Out[12]), .A2(
        SBOX_stage4Out[13]), .B1(SBOX_stage4Out[17]), .B2(SBOX_stage4Out[16]), 
        .ZN(SBOX_s5_mul2_1_1_n66) );
  XNOR2_X1 SBOX_s5_mul2_1_1_U22 ( .A(SBOX_s5_mul2_1_1_n64), .B(
        SBOX_s5_mul2_1_1_n65), .ZN(SBOX_s5_concat[31]) );
  XOR2_X1 SBOX_s5_mul2_1_1_U21 ( .A(SBOX_s5_mul2_1_1_n77), .B(
        SBOX_s5_mul2_1_1_n76), .Z(SBOX_s5_mul2_1_1_n65) );
  NAND2_X1 SBOX_s5_mul2_1_1_U20 ( .A1(SBOX_stage4Out[15]), .A2(
        SBOX_stage4Out[19]), .ZN(SBOX_s5_mul2_1_1_n64) );
  XNOR2_X1 SBOX_s5_mul2_1_1_U19 ( .A(SBOX_s5_mul2_1_1_n62), .B(
        SBOX_s5_mul2_1_1_n63), .ZN(SBOX_s5_concat[30]) );
  XOR2_X1 SBOX_s5_mul2_1_1_U18 ( .A(SBOX_s5_mul2_1_1_n75), .B(
        SBOX_s5_mul2_1_1_n76), .Z(SBOX_s5_mul2_1_1_n63) );
  NAND2_X1 SBOX_s5_mul2_1_1_U17 ( .A1(SBOX_stage4Out[14]), .A2(
        SBOX_stage4Out[18]), .ZN(SBOX_s5_mul2_1_1_n62) );
  XNOR2_X1 SBOX_s5_mul2_1_1_U16 ( .A(SBOX_s5_mul2_1_1_n60), .B(
        SBOX_s5_mul2_1_1_n61), .ZN(SBOX_s5_concat[29]) );
  XOR2_X1 SBOX_s5_mul2_1_1_U15 ( .A(SBOX_s5_mul2_1_1_n77), .B(
        SBOX_s5_mul2_1_1_n73), .Z(SBOX_s5_mul2_1_1_n61) );
  NAND2_X1 SBOX_s5_mul2_1_1_U14 ( .A1(SBOX_stage4Out[13]), .A2(
        SBOX_stage4Out[17]), .ZN(SBOX_s5_mul2_1_1_n60) );
  XNOR2_X1 SBOX_s5_mul2_1_1_U13 ( .A(SBOX_s5_mul2_1_1_n58), .B(
        SBOX_s5_mul2_1_1_n59), .ZN(SBOX_s5_concat[28]) );
  XOR2_X1 SBOX_s5_mul2_1_1_U12 ( .A(SBOX_s5_mul2_1_1_n73), .B(
        SBOX_s5_mul2_1_1_n75), .Z(SBOX_s5_mul2_1_1_n59) );
  NAND2_X1 SBOX_s5_mul2_1_1_U11 ( .A1(SBOX_stage4Out[12]), .A2(
        SBOX_stage4Out[16]), .ZN(SBOX_s5_mul2_1_1_n58) );
  INV_X1 SBOX_s5_mul2_1_1_U10 ( .A(SBOX_s5_mul2_1_1_n71), .ZN(
        SBOX_s5_mul2_1_1_n57) );
  INV_X1 SBOX_s5_mul2_1_1_U9 ( .A(SBOX_s5_mul2_1_1_n69), .ZN(
        SBOX_s5_mul2_1_1_n56) );
  XNOR2_X1 SBOX_s5_mul2_1_1_U8 ( .A(SBOX_s5_mul2_1_1_n54), .B(
        SBOX_s5_mul2_1_1_n70), .ZN(SBOX_s5_mul2_1_1_n55) );
  NAND2_X1 SBOX_s5_mul2_1_1_U7 ( .A1(SBOX_s5_mul2_1_1_n71), .A2(
        SBOX_s5_mul2_1_1_n72), .ZN(SBOX_s5_mul2_1_1_n54) );
  NAND2_X1 SBOX_s5_mul2_1_1_U5 ( .A1(SBOX_s5_mul2_1_1_n71), .A2(
        SBOX_s5_mul2_1_1_n69), .ZN(SBOX_s5_mul2_1_1_n67) );
  NOR2_X1 SBOX_s5_mul2_1_1_U4 ( .A1(SBOX_s5_mul2_1_1_n72), .A2(
        SBOX_s5_mul2_1_1_n70), .ZN(SBOX_s5_mul2_1_1_n68) );
  XNOR2_X1 SBOX_s5_mul2_1_1_U3 ( .A(SBOX_stage4Out[12]), .B(SBOX_stage4Out[14]), .ZN(SBOX_s5_mul2_1_1_n72) );
  XOR2_X1 SBOX_s5_mul2_1_1_U2 ( .A(SBOX_stage4Out[13]), .B(SBOX_stage4Out[15]), 
        .Z(SBOX_s5_mul2_1_1_n69) );
  OAI33_X1 SBOX_s5_mul2_1_1_U1 ( .A1(1'b0), .A2(SBOX_s5_mul2_1_1_n55), .A3(
        SBOX_s5_mul2_1_1_n56), .B1(SBOX_s5_mul2_1_1_n69), .B2(
        SBOX_s5_mul2_1_1_n72), .B3(SBOX_s5_mul2_1_1_n57), .ZN(
        SBOX_s5_mul2_1_1_n77) );
  AOI221_X1 SBOX_s5_mul2_1_0_U28 ( .B1(SBOX_stage4Out[2]), .B2(
        SBOX_stage4Out[3]), .C1(SBOX_stage4Out[18]), .C2(SBOX_stage4Out[19]), 
        .A(SBOX_s5_mul2_1_0_n73), .ZN(SBOX_s5_mul2_1_0_n75) );
  OAI22_X1 SBOX_s5_mul2_1_0_U27 ( .A1(SBOX_stage4Out[2]), .A2(
        SBOX_stage4Out[3]), .B1(SBOX_stage4Out[19]), .B2(SBOX_stage4Out[18]), 
        .ZN(SBOX_s5_mul2_1_0_n73) );
  XNOR2_X1 SBOX_s5_mul2_1_0_U26 ( .A(SBOX_s5_mul2_1_0_n63), .B(
        SBOX_s5_mul2_1_0_n62), .ZN(SBOX_s5_mul2_1_0_n74) );
  XOR2_X1 SBOX_s5_mul2_1_0_U25 ( .A(SBOX_stage4Out[17]), .B(SBOX_stage4Out[19]), .Z(SBOX_s5_mul2_1_0_n67) );
  XNOR2_X1 SBOX_s5_mul2_1_0_U24 ( .A(SBOX_stage4Out[16]), .B(
        SBOX_stage4Out[18]), .ZN(SBOX_s5_mul2_1_0_n66) );
  AOI221_X1 SBOX_s5_mul2_1_0_U23 ( .B1(SBOX_stage4Out[0]), .B2(
        SBOX_stage4Out[1]), .C1(SBOX_stage4Out[16]), .C2(SBOX_stage4Out[17]), 
        .A(SBOX_s5_mul2_1_0_n61), .ZN(SBOX_s5_mul2_1_0_n72) );
  OAI22_X1 SBOX_s5_mul2_1_0_U22 ( .A1(SBOX_stage4Out[0]), .A2(
        SBOX_stage4Out[1]), .B1(SBOX_stage4Out[17]), .B2(SBOX_stage4Out[16]), 
        .ZN(SBOX_s5_mul2_1_0_n61) );
  XNOR2_X1 SBOX_s5_mul2_1_0_U21 ( .A(SBOX_s5_mul2_1_0_n59), .B(
        SBOX_s5_mul2_1_0_n60), .ZN(SBOX_s5_concat[20]) );
  XOR2_X1 SBOX_s5_mul2_1_0_U20 ( .A(SBOX_s5_mul2_1_0_n74), .B(
        SBOX_s5_mul2_1_0_n72), .Z(SBOX_s5_mul2_1_0_n60) );
  NAND2_X1 SBOX_s5_mul2_1_0_U19 ( .A1(SBOX_stage4Out[0]), .A2(
        SBOX_stage4Out[16]), .ZN(SBOX_s5_mul2_1_0_n59) );
  XNOR2_X1 SBOX_s5_mul2_1_0_U18 ( .A(SBOX_s5_mul2_1_0_n57), .B(
        SBOX_s5_mul2_1_0_n58), .ZN(SBOX_s5_concat[23]) );
  XOR2_X1 SBOX_s5_mul2_1_0_U17 ( .A(SBOX_s5_mul2_1_0_n76), .B(
        SBOX_s5_mul2_1_0_n75), .Z(SBOX_s5_mul2_1_0_n58) );
  NAND2_X1 SBOX_s5_mul2_1_0_U16 ( .A1(SBOX_stage4Out[3]), .A2(
        SBOX_stage4Out[19]), .ZN(SBOX_s5_mul2_1_0_n57) );
  XNOR2_X1 SBOX_s5_mul2_1_0_U15 ( .A(SBOX_s5_mul2_1_0_n55), .B(
        SBOX_s5_mul2_1_0_n56), .ZN(SBOX_s5_concat[22]) );
  XOR2_X1 SBOX_s5_mul2_1_0_U14 ( .A(SBOX_s5_mul2_1_0_n75), .B(
        SBOX_s5_mul2_1_0_n74), .Z(SBOX_s5_mul2_1_0_n56) );
  NAND2_X1 SBOX_s5_mul2_1_0_U13 ( .A1(SBOX_stage4Out[2]), .A2(
        SBOX_stage4Out[18]), .ZN(SBOX_s5_mul2_1_0_n55) );
  XNOR2_X1 SBOX_s5_mul2_1_0_U12 ( .A(SBOX_s5_mul2_1_0_n53), .B(
        SBOX_s5_mul2_1_0_n54), .ZN(SBOX_s5_concat[21]) );
  XOR2_X1 SBOX_s5_mul2_1_0_U11 ( .A(SBOX_s5_mul2_1_0_n76), .B(
        SBOX_s5_mul2_1_0_n72), .Z(SBOX_s5_mul2_1_0_n54) );
  NAND2_X1 SBOX_s5_mul2_1_0_U10 ( .A1(SBOX_stage4Out[1]), .A2(
        SBOX_stage4Out[17]), .ZN(SBOX_s5_mul2_1_0_n53) );
  NAND2_X1 SBOX_s5_mul2_1_0_U9 ( .A1(SBOX_s5_mul2_1_0_n67), .A2(
        SBOX_s5_mul2_1_0_n69), .ZN(SBOX_s5_mul2_1_0_n65) );
  INV_X1 SBOX_s5_mul2_1_0_U8 ( .A(SBOX_s5_mul2_1_0_n64), .ZN(
        SBOX_s5_mul2_1_0_n71) );
  XNOR2_X1 SBOX_s5_mul2_1_0_U7 ( .A(SBOX_s5_mul2_1_0_n66), .B(
        SBOX_s5_mul2_1_0_n65), .ZN(SBOX_s5_mul2_1_0_n70) );
  NAND2_X1 SBOX_s5_mul2_1_0_U6 ( .A1(SBOX_s5_mul2_1_0_n67), .A2(
        SBOX_s5_mul2_1_0_n71), .ZN(SBOX_s5_mul2_1_0_n68) );
  OAI22_X1 SBOX_s5_mul2_1_0_U5 ( .A1(SBOX_s5_mul2_1_0_n71), .A2(
        SBOX_s5_mul2_1_0_n70), .B1(SBOX_s5_mul2_1_0_n69), .B2(
        SBOX_s5_mul2_1_0_n68), .ZN(SBOX_s5_mul2_1_0_n76) );
  NAND2_X1 SBOX_s5_mul2_1_0_U4 ( .A1(SBOX_s5_mul2_1_0_n67), .A2(
        SBOX_s5_mul2_1_0_n64), .ZN(SBOX_s5_mul2_1_0_n62) );
  NOR2_X1 SBOX_s5_mul2_1_0_U3 ( .A1(SBOX_s5_mul2_1_0_n69), .A2(
        SBOX_s5_mul2_1_0_n66), .ZN(SBOX_s5_mul2_1_0_n63) );
  XNOR2_X1 SBOX_s5_mul2_1_0_U2 ( .A(SBOX_stage4Out[0]), .B(SBOX_stage4Out[2]), 
        .ZN(SBOX_s5_mul2_1_0_n69) );
  XOR2_X1 SBOX_s5_mul2_1_0_U1 ( .A(SBOX_stage4Out[1]), .B(SBOX_stage4Out[3]), 
        .Z(SBOX_s5_mul2_1_0_n64) );
  AOI221_X1 SBOX_s5_mul2_0_1_U28 ( .B1(SBOX_stage4Out[14]), .B2(
        SBOX_stage4Out[15]), .C1(SBOX_stage4Out[6]), .C2(SBOX_stage4Out[7]), 
        .A(SBOX_s5_mul2_0_1_n73), .ZN(SBOX_s5_mul2_0_1_n75) );
  OAI22_X1 SBOX_s5_mul2_0_1_U27 ( .A1(SBOX_stage4Out[14]), .A2(
        SBOX_stage4Out[15]), .B1(SBOX_stage4Out[7]), .B2(SBOX_stage4Out[6]), 
        .ZN(SBOX_s5_mul2_0_1_n73) );
  XNOR2_X1 SBOX_s5_mul2_0_1_U26 ( .A(SBOX_s5_mul2_0_1_n63), .B(
        SBOX_s5_mul2_0_1_n62), .ZN(SBOX_s5_mul2_0_1_n74) );
  XOR2_X1 SBOX_s5_mul2_0_1_U25 ( .A(SBOX_stage4Out[5]), .B(SBOX_stage4Out[7]), 
        .Z(SBOX_s5_mul2_0_1_n67) );
  XNOR2_X1 SBOX_s5_mul2_0_1_U24 ( .A(SBOX_stage4Out[4]), .B(SBOX_stage4Out[6]), 
        .ZN(SBOX_s5_mul2_0_1_n66) );
  AOI221_X1 SBOX_s5_mul2_0_1_U23 ( .B1(SBOX_stage4Out[12]), .B2(
        SBOX_stage4Out[13]), .C1(SBOX_stage4Out[4]), .C2(SBOX_stage4Out[5]), 
        .A(SBOX_s5_mul2_0_1_n61), .ZN(SBOX_s5_mul2_0_1_n72) );
  OAI22_X1 SBOX_s5_mul2_0_1_U22 ( .A1(SBOX_stage4Out[12]), .A2(
        SBOX_stage4Out[13]), .B1(SBOX_stage4Out[5]), .B2(SBOX_stage4Out[4]), 
        .ZN(SBOX_s5_mul2_0_1_n61) );
  XNOR2_X1 SBOX_s5_mul2_0_1_U21 ( .A(SBOX_s5_mul2_0_1_n59), .B(
        SBOX_s5_mul2_0_1_n60), .ZN(SBOX_s5_concat[15]) );
  XOR2_X1 SBOX_s5_mul2_0_1_U20 ( .A(SBOX_s5_mul2_0_1_n76), .B(
        SBOX_s5_mul2_0_1_n75), .Z(SBOX_s5_mul2_0_1_n60) );
  NAND2_X1 SBOX_s5_mul2_0_1_U19 ( .A1(SBOX_stage4Out[15]), .A2(
        SBOX_stage4Out[7]), .ZN(SBOX_s5_mul2_0_1_n59) );
  XNOR2_X1 SBOX_s5_mul2_0_1_U18 ( .A(SBOX_s5_mul2_0_1_n57), .B(
        SBOX_s5_mul2_0_1_n58), .ZN(SBOX_s5_concat[14]) );
  XOR2_X1 SBOX_s5_mul2_0_1_U17 ( .A(SBOX_s5_mul2_0_1_n74), .B(
        SBOX_s5_mul2_0_1_n75), .Z(SBOX_s5_mul2_0_1_n58) );
  NAND2_X1 SBOX_s5_mul2_0_1_U16 ( .A1(SBOX_stage4Out[14]), .A2(
        SBOX_stage4Out[6]), .ZN(SBOX_s5_mul2_0_1_n57) );
  XNOR2_X1 SBOX_s5_mul2_0_1_U15 ( .A(SBOX_s5_mul2_0_1_n55), .B(
        SBOX_s5_mul2_0_1_n56), .ZN(SBOX_s5_concat[13]) );
  XOR2_X1 SBOX_s5_mul2_0_1_U14 ( .A(SBOX_s5_mul2_0_1_n76), .B(
        SBOX_s5_mul2_0_1_n72), .Z(SBOX_s5_mul2_0_1_n56) );
  NAND2_X1 SBOX_s5_mul2_0_1_U13 ( .A1(SBOX_stage4Out[13]), .A2(
        SBOX_stage4Out[5]), .ZN(SBOX_s5_mul2_0_1_n55) );
  XNOR2_X1 SBOX_s5_mul2_0_1_U12 ( .A(SBOX_s5_mul2_0_1_n53), .B(
        SBOX_s5_mul2_0_1_n54), .ZN(SBOX_s5_concat[12]) );
  XOR2_X1 SBOX_s5_mul2_0_1_U11 ( .A(SBOX_s5_mul2_0_1_n72), .B(
        SBOX_s5_mul2_0_1_n74), .Z(SBOX_s5_mul2_0_1_n54) );
  NAND2_X1 SBOX_s5_mul2_0_1_U10 ( .A1(SBOX_stage4Out[12]), .A2(
        SBOX_stage4Out[4]), .ZN(SBOX_s5_mul2_0_1_n53) );
  NAND2_X1 SBOX_s5_mul2_0_1_U9 ( .A1(SBOX_s5_mul2_0_1_n67), .A2(
        SBOX_s5_mul2_0_1_n69), .ZN(SBOX_s5_mul2_0_1_n65) );
  INV_X1 SBOX_s5_mul2_0_1_U8 ( .A(SBOX_s5_mul2_0_1_n64), .ZN(
        SBOX_s5_mul2_0_1_n71) );
  XNOR2_X1 SBOX_s5_mul2_0_1_U7 ( .A(SBOX_s5_mul2_0_1_n66), .B(
        SBOX_s5_mul2_0_1_n65), .ZN(SBOX_s5_mul2_0_1_n70) );
  NAND2_X1 SBOX_s5_mul2_0_1_U6 ( .A1(SBOX_s5_mul2_0_1_n67), .A2(
        SBOX_s5_mul2_0_1_n71), .ZN(SBOX_s5_mul2_0_1_n68) );
  OAI22_X1 SBOX_s5_mul2_0_1_U5 ( .A1(SBOX_s5_mul2_0_1_n71), .A2(
        SBOX_s5_mul2_0_1_n70), .B1(SBOX_s5_mul2_0_1_n69), .B2(
        SBOX_s5_mul2_0_1_n68), .ZN(SBOX_s5_mul2_0_1_n76) );
  NAND2_X1 SBOX_s5_mul2_0_1_U4 ( .A1(SBOX_s5_mul2_0_1_n67), .A2(
        SBOX_s5_mul2_0_1_n64), .ZN(SBOX_s5_mul2_0_1_n62) );
  NOR2_X1 SBOX_s5_mul2_0_1_U3 ( .A1(SBOX_s5_mul2_0_1_n69), .A2(
        SBOX_s5_mul2_0_1_n66), .ZN(SBOX_s5_mul2_0_1_n63) );
  XNOR2_X1 SBOX_s5_mul2_0_1_U2 ( .A(SBOX_stage4Out[12]), .B(SBOX_stage4Out[14]), .ZN(SBOX_s5_mul2_0_1_n69) );
  XOR2_X1 SBOX_s5_mul2_0_1_U1 ( .A(SBOX_stage4Out[13]), .B(SBOX_stage4Out[15]), 
        .Z(SBOX_s5_mul2_0_1_n64) );
  AOI221_X1 SBOX_s5_mul2_0_0_U28 ( .B1(SBOX_stage4Out[2]), .B2(
        SBOX_stage4Out[3]), .C1(SBOX_stage4Out[6]), .C2(SBOX_stage4Out[7]), 
        .A(SBOX_s5_mul2_0_0_n73), .ZN(SBOX_s5_mul2_0_0_n75) );
  OAI22_X1 SBOX_s5_mul2_0_0_U27 ( .A1(SBOX_stage4Out[2]), .A2(
        SBOX_stage4Out[3]), .B1(SBOX_stage4Out[7]), .B2(SBOX_stage4Out[6]), 
        .ZN(SBOX_s5_mul2_0_0_n73) );
  XNOR2_X1 SBOX_s5_mul2_0_0_U26 ( .A(SBOX_s5_mul2_0_0_n63), .B(
        SBOX_s5_mul2_0_0_n62), .ZN(SBOX_s5_mul2_0_0_n74) );
  XOR2_X1 SBOX_s5_mul2_0_0_U25 ( .A(SBOX_stage4Out[5]), .B(SBOX_stage4Out[7]), 
        .Z(SBOX_s5_mul2_0_0_n67) );
  XNOR2_X1 SBOX_s5_mul2_0_0_U24 ( .A(SBOX_stage4Out[4]), .B(SBOX_stage4Out[6]), 
        .ZN(SBOX_s5_mul2_0_0_n66) );
  AOI221_X1 SBOX_s5_mul2_0_0_U23 ( .B1(SBOX_stage4Out[0]), .B2(
        SBOX_stage4Out[1]), .C1(SBOX_stage4Out[4]), .C2(SBOX_stage4Out[5]), 
        .A(SBOX_s5_mul2_0_0_n61), .ZN(SBOX_s5_mul2_0_0_n72) );
  OAI22_X1 SBOX_s5_mul2_0_0_U22 ( .A1(SBOX_stage4Out[0]), .A2(
        SBOX_stage4Out[1]), .B1(SBOX_stage4Out[5]), .B2(SBOX_stage4Out[4]), 
        .ZN(SBOX_s5_mul2_0_0_n61) );
  XNOR2_X1 SBOX_s5_mul2_0_0_U21 ( .A(SBOX_s5_mul2_0_0_n59), .B(
        SBOX_s5_mul2_0_0_n60), .ZN(SBOX_s5_concat[7]) );
  XOR2_X1 SBOX_s5_mul2_0_0_U20 ( .A(SBOX_s5_mul2_0_0_n76), .B(
        SBOX_s5_mul2_0_0_n75), .Z(SBOX_s5_mul2_0_0_n60) );
  NAND2_X1 SBOX_s5_mul2_0_0_U19 ( .A1(SBOX_stage4Out[3]), .A2(
        SBOX_stage4Out[7]), .ZN(SBOX_s5_mul2_0_0_n59) );
  XNOR2_X1 SBOX_s5_mul2_0_0_U18 ( .A(SBOX_s5_mul2_0_0_n57), .B(
        SBOX_s5_mul2_0_0_n58), .ZN(SBOX_s5_concat[5]) );
  XOR2_X1 SBOX_s5_mul2_0_0_U17 ( .A(SBOX_s5_mul2_0_0_n76), .B(
        SBOX_s5_mul2_0_0_n72), .Z(SBOX_s5_mul2_0_0_n58) );
  NAND2_X1 SBOX_s5_mul2_0_0_U16 ( .A1(SBOX_stage4Out[1]), .A2(
        SBOX_stage4Out[5]), .ZN(SBOX_s5_mul2_0_0_n57) );
  XNOR2_X1 SBOX_s5_mul2_0_0_U15 ( .A(SBOX_s5_mul2_0_0_n55), .B(
        SBOX_s5_mul2_0_0_n56), .ZN(SBOX_s5_concat[6]) );
  XOR2_X1 SBOX_s5_mul2_0_0_U14 ( .A(SBOX_s5_mul2_0_0_n74), .B(
        SBOX_s5_mul2_0_0_n75), .Z(SBOX_s5_mul2_0_0_n56) );
  NAND2_X1 SBOX_s5_mul2_0_0_U13 ( .A1(SBOX_stage4Out[2]), .A2(
        SBOX_stage4Out[6]), .ZN(SBOX_s5_mul2_0_0_n55) );
  XNOR2_X1 SBOX_s5_mul2_0_0_U12 ( .A(SBOX_s5_mul2_0_0_n53), .B(
        SBOX_s5_mul2_0_0_n54), .ZN(SBOX_s5_concat[4]) );
  XOR2_X1 SBOX_s5_mul2_0_0_U11 ( .A(SBOX_s5_mul2_0_0_n72), .B(
        SBOX_s5_mul2_0_0_n74), .Z(SBOX_s5_mul2_0_0_n54) );
  NAND2_X1 SBOX_s5_mul2_0_0_U10 ( .A1(SBOX_stage4Out[0]), .A2(
        SBOX_stage4Out[4]), .ZN(SBOX_s5_mul2_0_0_n53) );
  NAND2_X1 SBOX_s5_mul2_0_0_U9 ( .A1(SBOX_s5_mul2_0_0_n67), .A2(
        SBOX_s5_mul2_0_0_n69), .ZN(SBOX_s5_mul2_0_0_n65) );
  INV_X1 SBOX_s5_mul2_0_0_U8 ( .A(SBOX_s5_mul2_0_0_n64), .ZN(
        SBOX_s5_mul2_0_0_n71) );
  XNOR2_X1 SBOX_s5_mul2_0_0_U7 ( .A(SBOX_s5_mul2_0_0_n66), .B(
        SBOX_s5_mul2_0_0_n65), .ZN(SBOX_s5_mul2_0_0_n70) );
  NAND2_X1 SBOX_s5_mul2_0_0_U6 ( .A1(SBOX_s5_mul2_0_0_n67), .A2(
        SBOX_s5_mul2_0_0_n71), .ZN(SBOX_s5_mul2_0_0_n68) );
  OAI22_X1 SBOX_s5_mul2_0_0_U5 ( .A1(SBOX_s5_mul2_0_0_n71), .A2(
        SBOX_s5_mul2_0_0_n70), .B1(SBOX_s5_mul2_0_0_n69), .B2(
        SBOX_s5_mul2_0_0_n68), .ZN(SBOX_s5_mul2_0_0_n76) );
  NAND2_X1 SBOX_s5_mul2_0_0_U4 ( .A1(SBOX_s5_mul2_0_0_n67), .A2(
        SBOX_s5_mul2_0_0_n64), .ZN(SBOX_s5_mul2_0_0_n62) );
  NOR2_X1 SBOX_s5_mul2_0_0_U3 ( .A1(SBOX_s5_mul2_0_0_n69), .A2(
        SBOX_s5_mul2_0_0_n66), .ZN(SBOX_s5_mul2_0_0_n63) );
  XNOR2_X1 SBOX_s5_mul2_0_0_U2 ( .A(SBOX_stage4Out[0]), .B(SBOX_stage4Out[2]), 
        .ZN(SBOX_s5_mul2_0_0_n69) );
  XOR2_X1 SBOX_s5_mul2_0_0_U1 ( .A(SBOX_stage4Out[1]), .B(SBOX_stage4Out[3]), 
        .Z(SBOX_s5_mul2_0_0_n64) );
  XOR2_X1 SBOX_s5_compr_0_0_U8 ( .A(SBOX_s5_regOut[7]), .B(SBOX_s5_regOut[15]), 
        .Z(SBOX_stage5Out[7]) );
  XOR2_X1 SBOX_s5_compr_0_0_U7 ( .A(SBOX_s5_regOut[6]), .B(SBOX_s5_regOut[14]), 
        .Z(SBOX_stage5Out[6]) );
  XOR2_X1 SBOX_s5_compr_0_0_U6 ( .A(SBOX_s5_regOut[5]), .B(SBOX_s5_regOut[13]), 
        .Z(SBOX_stage5Out[5]) );
  XOR2_X1 SBOX_s5_compr_0_0_U5 ( .A(SBOX_s5_regOut[4]), .B(SBOX_s5_regOut[12]), 
        .Z(SBOX_stage5Out[4]) );
  XOR2_X1 SBOX_s5_compr_0_0_U4 ( .A(SBOX_s5_regOut[3]), .B(SBOX_s5_regOut[11]), 
        .Z(SBOX_stage5Out[3]) );
  XOR2_X1 SBOX_s5_compr_0_0_U3 ( .A(SBOX_s5_regOut[1]), .B(SBOX_s5_regOut[9]), 
        .Z(SBOX_stage5Out[1]) );
  XOR2_X1 SBOX_s5_compr_0_0_U2 ( .A(SBOX_s5_regOut[0]), .B(SBOX_s5_regOut[8]), 
        .Z(SBOX_stage5Out[0]) );
  XOR2_X1 SBOX_s5_compr_0_0_U1 ( .A(SBOX_s5_regOut[2]), .B(SBOX_s5_regOut[10]), 
        .Z(SBOX_stage5Out[2]) );
  XOR2_X1 SBOX_s5_compr_1_0_U8 ( .A(SBOX_s5_regOut[23]), .B(SBOX_s5_regOut[31]), .Z(SBOX_stage5Out[15]) );
  XOR2_X1 SBOX_s5_compr_1_0_U7 ( .A(SBOX_s5_regOut[22]), .B(SBOX_s5_regOut[30]), .Z(SBOX_stage5Out[14]) );
  XOR2_X1 SBOX_s5_compr_1_0_U6 ( .A(SBOX_s5_regOut[21]), .B(SBOX_s5_regOut[29]), .Z(SBOX_stage5Out[13]) );
  XOR2_X1 SBOX_s5_compr_1_0_U5 ( .A(SBOX_s5_regOut[20]), .B(SBOX_s5_regOut[28]), .Z(SBOX_stage5Out[12]) );
  XOR2_X1 SBOX_s5_compr_1_0_U4 ( .A(SBOX_s5_regOut[19]), .B(SBOX_s5_regOut[27]), .Z(SBOX_stage5Out[11]) );
  XOR2_X1 SBOX_s5_compr_1_0_U3 ( .A(SBOX_s5_regOut[17]), .B(SBOX_s5_regOut[25]), .Z(SBOX_stage5Out[9]) );
  XOR2_X1 SBOX_s5_compr_1_0_U2 ( .A(SBOX_s5_regOut[16]), .B(SBOX_s5_regOut[24]), .Z(SBOX_stage5Out[8]) );
  XOR2_X1 SBOX_s5_compr_1_0_U1 ( .A(SBOX_s5_regOut[18]), .B(SBOX_s5_regOut[26]), .Z(SBOX_stage5Out[10]) );
  XOR2_X1 SBOX_s6_1_U11 ( .A(SBOX_stage5Out[14]), .B(SBOX_stage5Out[8]), .Z(
        SBOX_stage6Out[13]) );
  XNOR2_X1 SBOX_s6_1_U10 ( .A(SBOX_s6_1_n8), .B(SBOX_stage5Out[9]), .ZN(
        SBOX_stage6Out[9]) );
  XNOR2_X1 SBOX_s6_1_U9 ( .A(SBOX_stage5Out[13]), .B(SBOX_stage5Out[12]), .ZN(
        SBOX_s6_1_n8) );
  XNOR2_X1 SBOX_s6_1_U8 ( .A(SBOX_s6_1_n7), .B(SBOX_stage6Out[13]), .ZN(
        SBOX_stage6Out[10]) );
  XNOR2_X1 SBOX_s6_1_U7 ( .A(SBOX_stage6Out[15]), .B(SBOX_stage5Out[10]), .ZN(
        SBOX_s6_1_n7) );
  XOR2_X1 SBOX_s6_1_U6 ( .A(SBOX_stage5Out[11]), .B(SBOX_stage5Out[13]), .Z(
        SBOX_stage6Out[15]) );
  XOR2_X1 SBOX_s6_1_U5 ( .A(SBOX_stage5Out[11]), .B(SBOX_stage5Out[15]), .Z(
        SBOX_stage6Out[14]) );
  XOR2_X1 SBOX_s6_1_U4 ( .A(SBOX_stage6Out[15]), .B(SBOX_stage5Out[15]), .Z(
        SBOX_stage6Out[12]) );
  XNOR2_X1 SBOX_s6_1_U3 ( .A(SBOX_stage6Out[12]), .B(SBOX_s6_1_n9), .ZN(
        SBOX_stage6Out[11]) );
  XNOR2_X1 SBOX_s6_1_U2 ( .A(SBOX_stage5Out[9]), .B(SBOX_s6_1_n9), .ZN(
        SBOX_stage6Out[8]) );
  XNOR2_X1 SBOX_s6_1_U1 ( .A(SBOX_stage5Out[14]), .B(SBOX_stage5Out[12]), .ZN(
        SBOX_s6_1_n9) );
  XOR2_X1 SBOX_s6_0_U11 ( .A(SBOX_stage5Out[6]), .B(SBOX_stage5Out[0]), .Z(
        SBOX_stage6Out[5]) );
  XNOR2_X1 SBOX_s6_0_U10 ( .A(SBOX_s6_0_n8), .B(SBOX_stage5Out[1]), .ZN(
        SBOX_stage6Out[1]) );
  XNOR2_X1 SBOX_s6_0_U9 ( .A(SBOX_stage5Out[5]), .B(SBOX_stage5Out[4]), .ZN(
        SBOX_s6_0_n8) );
  XNOR2_X1 SBOX_s6_0_U8 ( .A(SBOX_s6_0_n7), .B(SBOX_stage6Out[5]), .ZN(
        SBOX_stage6Out[2]) );
  XNOR2_X1 SBOX_s6_0_U7 ( .A(SBOX_stage6Out[7]), .B(SBOX_stage5Out[2]), .ZN(
        SBOX_s6_0_n7) );
  XOR2_X1 SBOX_s6_0_U6 ( .A(SBOX_stage5Out[3]), .B(SBOX_stage5Out[5]), .Z(
        SBOX_stage6Out[7]) );
  XOR2_X1 SBOX_s6_0_U5 ( .A(SBOX_stage5Out[3]), .B(SBOX_stage5Out[7]), .Z(
        SBOX_stage6Out[6]) );
  XOR2_X1 SBOX_s6_0_U4 ( .A(SBOX_stage6Out[7]), .B(SBOX_stage5Out[7]), .Z(
        SBOX_stage6Out[4]) );
  XNOR2_X1 SBOX_s6_0_U3 ( .A(SBOX_stage6Out[4]), .B(SBOX_s6_0_n9), .ZN(
        SBOX_stage6Out[3]) );
  XNOR2_X1 SBOX_s6_0_U2 ( .A(SBOX_stage5Out[1]), .B(SBOX_s6_0_n9), .ZN(
        SBOX_stage6Out[0]) );
  XNOR2_X1 SBOX_s6_0_U1 ( .A(SBOX_stage5Out[6]), .B(SBOX_stage5Out[4]), .ZN(
        SBOX_s6_0_n9) );
  BUF_X1 aes_key_regs_1_U3 ( .A(n114), .Z(aes_key_regs_1_n4) );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_0_ ( .D(aes_key_regs_1_K00xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[8]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_0_ ( .D(aes_key_regs_1_K10xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_0_ ( .D(aes_key_regs_1_K20xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_0_ ( .D(aes_key_regs_1_K01xDP_0_), .SI(
        KeyOutxD[8]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_0_ ( .D(aes_key_regs_1_K01xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_0_ ( .D(aes_key_regs_1_K11xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_0_ ( .D(aes_key_regs_1_K21xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_0_ ( .D(aes_key_regs_1_K02xDP_0_), .SI(
        aes_key_regs_1_K01xDP_0_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_0_ ( .D(aes_key_regs_1_K02xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_0_ ( .D(aes_key_regs_1_K12xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_0_ ( .D(aes_key_regs_1_K22xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_0_ ( .D(K03xD[8]), .SI(
        aes_key_regs_1_K02xDP_0_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_1_ ( .D(aes_key_regs_1_K00xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[9]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_1_ ( .D(aes_key_regs_1_K10xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_1_ ( .D(aes_key_regs_1_K20xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_1_ ( .D(aes_key_regs_1_K01xDP_1_), .SI(
        KeyOutxD[9]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K20xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_1_ ( .D(aes_key_regs_1_K01xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_1_ ( .D(aes_key_regs_1_K11xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_1_ ( .D(aes_key_regs_1_K21xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_1_ ( .D(aes_key_regs_1_K02xDP_1_), .SI(
        aes_key_regs_1_K01xDP_1_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K21xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_1_ ( .D(aes_key_regs_1_K02xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_1_ ( .D(aes_key_regs_1_K12xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_1_ ( .D(aes_key_regs_1_K22xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_1_ ( .D(K03xD[9]), .SI(
        aes_key_regs_1_K02xDP_1_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K22xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_2_ ( .D(aes_key_regs_1_K00xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[10]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_2_ ( .D(aes_key_regs_1_K10xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_2_ ( .D(aes_key_regs_1_K20xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_2_ ( .D(aes_key_regs_1_K01xDP_2_), .SI(
        KeyOutxD[10]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_2_ ( .D(aes_key_regs_1_K01xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_2_ ( .D(aes_key_regs_1_K11xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_2_ ( .D(aes_key_regs_1_K21xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_2_ ( .D(aes_key_regs_1_K02xDP_2_), .SI(
        aes_key_regs_1_K01xDP_2_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K21xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_2_ ( .D(aes_key_regs_1_K02xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_2_ ( .D(aes_key_regs_1_K12xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_2_ ( .D(aes_key_regs_1_K22xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_2_ ( .D(K03xD[10]), .SI(
        aes_key_regs_1_K02xDP_2_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K22xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_3_ ( .D(aes_key_regs_1_K00xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[11]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_3_ ( .D(aes_key_regs_1_K10xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_3_ ( .D(aes_key_regs_1_K20xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_3_ ( .D(aes_key_regs_1_K01xDP_3_), .SI(
        KeyOutxD[11]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K20xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_3_ ( .D(aes_key_regs_1_K01xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_3_ ( .D(aes_key_regs_1_K11xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_3_ ( .D(aes_key_regs_1_K21xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_3_ ( .D(aes_key_regs_1_K02xDP_3_), .SI(
        aes_key_regs_1_K01xDP_3_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K21xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_3_ ( .D(aes_key_regs_1_K02xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_3_ ( .D(aes_key_regs_1_K12xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_3_ ( .D(aes_key_regs_1_K22xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_3_ ( .D(K03xD[11]), .SI(
        aes_key_regs_1_K02xDP_3_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K22xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_4_ ( .D(aes_key_regs_1_K00xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[12]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_4_ ( .D(aes_key_regs_1_K10xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_4_ ( .D(aes_key_regs_1_K20xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_4_ ( .D(aes_key_regs_1_K01xDP_4_), .SI(
        KeyOutxD[12]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_4_ ( .D(aes_key_regs_1_K01xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_4_ ( .D(aes_key_regs_1_K11xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_4_ ( .D(aes_key_regs_1_K21xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_4_ ( .D(aes_key_regs_1_K02xDP_4_), .SI(
        aes_key_regs_1_K01xDP_4_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_4_ ( .D(aes_key_regs_1_K02xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_4_ ( .D(aes_key_regs_1_K12xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_4_ ( .D(aes_key_regs_1_K22xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_4_ ( .D(K03xD[12]), .SI(
        aes_key_regs_1_K02xDP_4_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_5_ ( .D(aes_key_regs_1_K00xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[13]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_5_ ( .D(aes_key_regs_1_K10xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_5_ ( .D(aes_key_regs_1_K20xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_5_ ( .D(aes_key_regs_1_K01xDP_5_), .SI(
        KeyOutxD[13]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K20xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_5_ ( .D(aes_key_regs_1_K01xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_5_ ( .D(aes_key_regs_1_K11xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_5_ ( .D(aes_key_regs_1_K21xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_5_ ( .D(aes_key_regs_1_K02xDP_5_), .SI(
        aes_key_regs_1_K01xDP_5_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K21xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_5_ ( .D(aes_key_regs_1_K02xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_5_ ( .D(aes_key_regs_1_K12xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_5_ ( .D(aes_key_regs_1_K22xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_5_ ( .D(K03xD[13]), .SI(
        aes_key_regs_1_K02xDP_5_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_6_ ( .D(aes_key_regs_1_K00xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[14]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_6_ ( .D(aes_key_regs_1_K10xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_6_ ( .D(aes_key_regs_1_K20xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_6_ ( .D(aes_key_regs_1_K01xDP_6_), .SI(
        KeyOutxD[14]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_6_ ( .D(aes_key_regs_1_K01xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_6_ ( .D(aes_key_regs_1_K11xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_6_ ( .D(aes_key_regs_1_K21xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_6_ ( .D(aes_key_regs_1_K02xDP_6_), .SI(
        aes_key_regs_1_K01xDP_6_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_6_ ( .D(aes_key_regs_1_K02xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_6_ ( .D(aes_key_regs_1_K12xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_6_ ( .D(aes_key_regs_1_K22xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_6_ ( .D(K03xD[14]), .SI(
        aes_key_regs_1_K02xDP_6_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_7_ ( .D(aes_key_regs_1_K00xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[15]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_7_ ( .D(aes_key_regs_1_K10xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_7_ ( .D(aes_key_regs_1_K20xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_7_ ( .D(aes_key_regs_1_K01xDP_7_), .SI(
        KeyOutxD[15]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_7_ ( .D(aes_key_regs_1_K01xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_7_ ( .D(aes_key_regs_1_K11xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_7_ ( .D(aes_key_regs_1_K21xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_7_ ( .D(aes_key_regs_1_K02xDP_7_), .SI(
        aes_key_regs_1_K01xDP_7_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_7_ ( .D(aes_key_regs_1_K02xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_7_ ( .D(aes_key_regs_1_K12xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_7_ ( .D(aes_key_regs_1_K22xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_7_ ( .D(K03xD[15]), .SI(
        aes_key_regs_1_K02xDP_7_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K22xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_0_ ( .D(KeyInxD[8]), .SI(K03xD[8]), .SE(
        aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_0_ ( .D(KeyToSboxOutxD[8]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[8]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_0_ ( .D(aes_key_regs_1_K13xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[8]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_0_ ( .D(aes_key_regs_1_K23xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_1_ ( .D(KeyInxD[9]), .SI(K03xD[9]), .SE(
        aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_1_ ( .D(KeyToSboxOutxD[9]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[9]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_1_ ( .D(aes_key_regs_1_K13xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[9]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_1_ ( .D(aes_key_regs_1_K23xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_2_ ( .D(KeyInxD[10]), .SI(K03xD[10]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_2_ ( .D(KeyToSboxOutxD[10]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[10]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_2_ ( .D(aes_key_regs_1_K13xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[10]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_2_ ( .D(aes_key_regs_1_K23xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_3_ ( .D(KeyInxD[11]), .SI(K03xD[11]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_3_ ( .D(KeyToSboxOutxD[11]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[11]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_3_ ( .D(aes_key_regs_1_K13xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[11]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_3_ ( .D(aes_key_regs_1_K23xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_4_ ( .D(KeyInxD[12]), .SI(K03xD[12]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_4_ ( .D(KeyToSboxOutxD[12]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[12]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_4_ ( .D(aes_key_regs_1_K13xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[12]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_4_ ( .D(aes_key_regs_1_K23xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_5_ ( .D(KeyInxD[13]), .SI(K03xD[13]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_5_ ( .D(KeyToSboxOutxD[13]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[13]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_5_ ( .D(aes_key_regs_1_K13xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[13]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_5_ ( .D(aes_key_regs_1_K23xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_6_ ( .D(KeyInxD[14]), .SI(K03xD[14]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_6_ ( .D(KeyToSboxOutxD[14]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[14]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_6_ ( .D(aes_key_regs_1_K13xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[14]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_6_ ( .D(aes_key_regs_1_K23xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_7_ ( .D(KeyInxD[15]), .SI(K03xD[15]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_7_ ( .D(KeyToSboxOutxD[15]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[15]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_7_ ( .D(aes_key_regs_1_K13xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[15]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_7_ ( .D(aes_key_regs_1_K23xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[7]), .QN() );
  OAI222_X1 aes_state_regs_1_U55 ( .A1(aes_state_regs_1_n79), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n80), .B2(
        aes_state_regs_1_n98), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n47), .ZN(aes_state_regs_1_S10xDN[7]) );
  INV_X1 aes_state_regs_1_U54 ( .A(aes_state_regs_1_MixColumnsS2xD[7]), .ZN(
        aes_state_regs_1_n79) );
  OAI222_X1 aes_state_regs_1_U53 ( .A1(aes_state_regs_1_n78), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n80), .B2(
        aes_state_regs_1_n99), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n48), .ZN(aes_state_regs_1_S10xDN[6]) );
  INV_X1 aes_state_regs_1_U52 ( .A(aes_state_regs_1_MixColumnsS2xD[6]), .ZN(
        aes_state_regs_1_n78) );
  OAI222_X1 aes_state_regs_1_U51 ( .A1(aes_state_regs_1_n77), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n80), .B2(
        aes_state_regs_1_n100), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n49), .ZN(aes_state_regs_1_S10xDN[5]) );
  INV_X1 aes_state_regs_1_U50 ( .A(aes_state_regs_1_MixColumnsS2xD[5]), .ZN(
        aes_state_regs_1_n77) );
  OAI222_X1 aes_state_regs_1_U49 ( .A1(aes_state_regs_1_n76), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n80), .B2(
        aes_state_regs_1_n101), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n50), .ZN(aes_state_regs_1_S10xDN[4]) );
  INV_X1 aes_state_regs_1_U48 ( .A(aes_state_regs_1_MixColumnsS2xD[4]), .ZN(
        aes_state_regs_1_n76) );
  OAI222_X1 aes_state_regs_1_U47 ( .A1(aes_state_regs_1_n75), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n80), .B2(
        aes_state_regs_1_n102), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n51), .ZN(aes_state_regs_1_S10xDN[3]) );
  INV_X1 aes_state_regs_1_U46 ( .A(aes_state_regs_1_MixColumnsS2xD[3]), .ZN(
        aes_state_regs_1_n75) );
  INV_X1 aes_state_regs_1_U45 ( .A(nextRCONxS), .ZN(aes_state_regs_1_n74) );
  INV_X4 aes_state_regs_1_U44 ( .A(aes_state_regs_1_n74), .ZN(
        aes_state_regs_1_n73) );
  OAI222_X1 aes_state_regs_1_U43 ( .A1(aes_state_regs_1_n70), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n62), .C1(aes_state_regs_1_n80), .C2(
        aes_state_regs_1_n97), .ZN(aes_state_regs_1_S20xDN[0]) );
  INV_X1 aes_state_regs_1_U42 ( .A(aes_state_regs_1_MixColumnsS3xD[0]), .ZN(
        aes_state_regs_1_n70) );
  OAI222_X1 aes_state_regs_1_U41 ( .A1(aes_state_regs_1_n69), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n80), .B2(
        aes_state_regs_1_n105), .C1(aes_state_regs_1_n54), .C2(
        aes_state_regs_1_n74), .ZN(aes_state_regs_1_S10xDN[0]) );
  INV_X1 aes_state_regs_1_U40 ( .A(aes_state_regs_1_MixColumnsS2xD[0]), .ZN(
        aes_state_regs_1_n69) );
  OAI222_X1 aes_state_regs_1_U39 ( .A1(aes_state_regs_1_n68), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n60), .C1(aes_state_regs_1_n80), .C2(
        aes_state_regs_1_n95), .ZN(aes_state_regs_1_S20xDN[2]) );
  INV_X1 aes_state_regs_1_U38 ( .A(aes_state_regs_1_MixColumnsS3xD[2]), .ZN(
        aes_state_regs_1_n68) );
  OAI21_X1 aes_state_regs_1_U37 ( .B1(aes_state_regs_1_n91), .B2(
        aes_state_regs_1_n80), .A(aes_state_regs_1_n67), .ZN(
        aes_state_regs_1_S20xDN[6]) );
  AOI22_X1 aes_state_regs_1_U36 ( .A1(aes_state_regs_1_MixColumnsS3xD[6]), 
        .A2(aes_state_regs_1_n71), .B1(aes_state_regs_1_n8), .B2(
        aes_state_regs_1_n73), .ZN(aes_state_regs_1_n67) );
  OAI222_X1 aes_state_regs_1_U35 ( .A1(aes_state_regs_1_n66), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n61), .C1(aes_state_regs_1_n80), .C2(
        aes_state_regs_1_n96), .ZN(aes_state_regs_1_S20xDN[1]) );
  INV_X1 aes_state_regs_1_U34 ( .A(aes_state_regs_1_MixColumnsS3xD[1]), .ZN(
        aes_state_regs_1_n66) );
  OAI222_X1 aes_state_regs_1_U33 ( .A1(aes_state_regs_1_n65), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n59), .C1(aes_state_regs_1_n80), .C2(
        aes_state_regs_1_n94), .ZN(aes_state_regs_1_S20xDN[3]) );
  INV_X1 aes_state_regs_1_U32 ( .A(aes_state_regs_1_MixColumnsS3xD[3]), .ZN(
        aes_state_regs_1_n65) );
  OAI222_X1 aes_state_regs_1_U31 ( .A1(aes_state_regs_1_n64), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n58), .C1(aes_state_regs_1_n80), .C2(
        aes_state_regs_1_n93), .ZN(aes_state_regs_1_S20xDN[4]) );
  INV_X1 aes_state_regs_1_U30 ( .A(aes_state_regs_1_MixColumnsS3xD[4]), .ZN(
        aes_state_regs_1_n64) );
  OAI222_X1 aes_state_regs_1_U29 ( .A1(aes_state_regs_1_n63), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n57), .C1(aes_state_regs_1_n80), .C2(
        aes_state_regs_1_n92), .ZN(aes_state_regs_1_S20xDN[5]) );
  INV_X1 aes_state_regs_1_U28 ( .A(aes_state_regs_1_MixColumnsS3xD[5]), .ZN(
        aes_state_regs_1_n63) );
  OAI222_X1 aes_state_regs_1_U27 ( .A1(aes_state_regs_1_n56), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n55), .C1(aes_state_regs_1_n80), .C2(
        aes_state_regs_1_n90), .ZN(aes_state_regs_1_S20xDN[7]) );
  INV_X1 aes_state_regs_1_U26 ( .A(aes_state_regs_1_MixColumnsS3xD[7]), .ZN(
        aes_state_regs_1_n56) );
  OAI222_X1 aes_state_regs_1_U25 ( .A1(aes_state_regs_1_n46), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n53), .C1(aes_state_regs_1_n104), .C2(
        aes_state_regs_1_n80), .ZN(aes_state_regs_1_S10xDN[1]) );
  INV_X1 aes_state_regs_1_U24 ( .A(aes_state_regs_1_MixColumnsS2xD[1]), .ZN(
        aes_state_regs_1_n46) );
  OAI222_X1 aes_state_regs_1_U23 ( .A1(aes_state_regs_1_n45), .A2(
        aes_state_regs_1_n72), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n52), .C1(aes_state_regs_1_n80), .C2(
        aes_state_regs_1_n103), .ZN(aes_state_regs_1_S10xDN[2]) );
  INV_X1 aes_state_regs_1_U22 ( .A(aes_state_regs_1_MixColumnsS2xD[2]), .ZN(
        aes_state_regs_1_n45) );
  INV_X2 aes_state_regs_1_U21 ( .A(aes_state_regs_1_n71), .ZN(
        aes_state_regs_1_n72) );
  NAND2_X1 aes_state_regs_1_U20 ( .A1(aes_state_regs_1_n71), .A2(
        aes_state_regs_1_MixColumnsS0xD[7]), .ZN(aes_state_regs_1_n81) );
  OAI21_X1 aes_state_regs_1_U19 ( .B1(aes_state_regs_1_n71), .B2(
        aes_state_regs_1_n82), .A(aes_state_regs_1_n81), .ZN(StateOutxD[15])
         );
  NAND2_X1 aes_state_regs_1_U18 ( .A1(aes_state_regs_1_n71), .A2(
        aes_state_regs_1_MixColumnsS0xD[4]), .ZN(aes_state_regs_1_n108) );
  OAI21_X1 aes_state_regs_1_U17 ( .B1(aes_state_regs_1_n71), .B2(
        aes_state_regs_1_n86), .A(aes_state_regs_1_n108), .ZN(StateOutxD[12])
         );
  NAND2_X1 aes_state_regs_1_U16 ( .A1(aes_state_regs_1_n71), .A2(
        aes_state_regs_1_MixColumnsS0xD[3]), .ZN(aes_state_regs_1_n109) );
  OAI21_X1 aes_state_regs_1_U15 ( .B1(aes_state_regs_1_n71), .B2(
        aes_state_regs_1_n85), .A(aes_state_regs_1_n109), .ZN(StateOutxD[11])
         );
  NAND2_X1 aes_state_regs_1_U14 ( .A1(aes_state_regs_1_n71), .A2(
        aes_state_regs_1_MixColumnsS0xD[2]), .ZN(aes_state_regs_1_n110) );
  OAI21_X1 aes_state_regs_1_U13 ( .B1(aes_state_regs_1_n71), .B2(
        aes_state_regs_1_n84), .A(aes_state_regs_1_n110), .ZN(StateOutxD[10])
         );
  NAND2_X1 aes_state_regs_1_U12 ( .A1(aes_state_regs_1_n71), .A2(
        aes_state_regs_1_MixColumnsS0xD[1]), .ZN(aes_state_regs_1_n111) );
  OAI21_X1 aes_state_regs_1_U11 ( .B1(aes_state_regs_1_n71), .B2(
        aes_state_regs_1_n83), .A(aes_state_regs_1_n111), .ZN(StateOutxD[9])
         );
  OR2_X1 aes_state_regs_1_U10 ( .A1(aes_state_regs_1_n73), .A2(doMixColumnsxS), 
        .ZN(aes_state_regs_1_n80) );
  AND2_X2 aes_state_regs_1_U9 ( .A1(doMixColumnsxS), .A2(aes_state_regs_1_n74), 
        .ZN(aes_state_regs_1_n71) );
  NAND2_X1 aes_state_regs_1_U8 ( .A1(aes_state_regs_1_n71), .A2(
        aes_state_regs_1_MixColumnsS0xD[0]), .ZN(aes_state_regs_1_n112) );
  OAI21_X1 aes_state_regs_1_U7 ( .B1(aes_state_regs_1_n71), .B2(
        aes_state_regs_1_n89), .A(aes_state_regs_1_n112), .ZN(StateOutxD[8])
         );
  NAND2_X1 aes_state_regs_1_U6 ( .A1(aes_state_regs_1_n71), .A2(
        aes_state_regs_1_MixColumnsS0xD[6]), .ZN(aes_state_regs_1_n106) );
  OAI21_X1 aes_state_regs_1_U5 ( .B1(aes_state_regs_1_n71), .B2(
        aes_state_regs_1_n88), .A(aes_state_regs_1_n106), .ZN(StateOutxD[14])
         );
  NAND2_X1 aes_state_regs_1_U4 ( .A1(aes_state_regs_1_n71), .A2(
        aes_state_regs_1_MixColumnsS0xD[5]), .ZN(aes_state_regs_1_n107) );
  OAI21_X1 aes_state_regs_1_U3 ( .B1(aes_state_regs_1_n71), .B2(
        aes_state_regs_1_n87), .A(aes_state_regs_1_n107), .ZN(StateOutxD[13])
         );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_7_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[7]), .SI(aes_state_regs_1_S10xDP_7_), 
        .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[7]), .QN(aes_state_regs_1_n82) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_6_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[6]), .SI(aes_state_regs_1_S10xDP_6_), 
        .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[6]), .QN(aes_state_regs_1_n88) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_5_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[5]), .SI(aes_state_regs_1_S10xDP_5_), 
        .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[5]), .QN(aes_state_regs_1_n87) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_4_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[4]), .SI(aes_state_regs_1_S10xDP_4_), 
        .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[4]), .QN(aes_state_regs_1_n86) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_3_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[3]), .SI(aes_state_regs_1_S10xDP_3_), 
        .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[3]), .QN(aes_state_regs_1_n85) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_2_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[2]), .SI(aes_state_regs_1_S10xDP_2_), 
        .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[2]), .QN(aes_state_regs_1_n84) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_1_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[1]), .SI(aes_state_regs_1_S10xDP_1_), 
        .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[1]), .QN(aes_state_regs_1_n83) );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_7_ ( .D(aes_state_regs_1_S10xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_7_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_6_ ( .D(aes_state_regs_1_S10xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_6_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_5_ ( .D(aes_state_regs_1_S10xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_5_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_4_ ( .D(aes_state_regs_1_S10xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_4_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_3_ ( .D(aes_state_regs_1_S10xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_3_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_2_ ( .D(aes_state_regs_1_S10xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_2_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_1_ ( .D(aes_state_regs_1_S10xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_7_ ( .D(aes_state_regs_1_S01xDO_7_), 
        .SI(StateInxD[15]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_7_), .QN(aes_state_regs_1_n90) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_7_ ( .D(aes_state_regs_1_n1), .SI(
        aes_state_regs_1_n4), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[7]), .QN(aes_state_regs_1_n47) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_7_ ( .D(aes_state_regs_1_S02xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_7_ ( .D(aes_state_regs_1_n2), .SI(
        aes_state_regs_1_S23xDP_7_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_7_ ( .D(aes_state_regs_1_n4), .SI(
        aes_state_regs_1_n1), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_7_ ( .D(aes_state_regs_1_S02xDP_7_), 
        .SI(aes_state_regs_1_S01xDO_7_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n1), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_7_ ( .D(aes_state_regs_1_S01xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_7_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_7_ ( .D(aes_state_regs_1_S21xDP[7]), 
        .SI(aes_state_regs_1_n2), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S01xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_7_ ( .D(aes_state_regs_1_n3), .SI(
        aes_state_regs_1_S30xDP_7_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n2), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_7_ ( .D(aes_state_regs_1_n5), .SI(
        aes_state_regs_1_S02xDP_7_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n3), .QN(aes_state_regs_1_n55) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_7_ ( .D(StateInxD[15]), .SI(
        aes_state_regs_1_n5), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n4), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_7_ ( .D(aes_state_regs_1_S03xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n5), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_7_ ( .D(aes_state_regs_1_S23xDP_7_), 
        .SI(aes_state_regs_1_S20xDP_7_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[7]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_7_ ( .D(aes_state_regs_1_S20xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_7_), .QN(
        aes_state_regs_1_n98) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_6_ ( .D(aes_state_regs_1_S01xDO_6_), 
        .SI(StateInxD[14]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_6_), .QN(aes_state_regs_1_n91) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_6_ ( .D(aes_state_regs_1_n6), .SI(
        aes_state_regs_1_n9), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[6]), .QN(aes_state_regs_1_n48) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_6_ ( .D(aes_state_regs_1_S02xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_6_ ( .D(aes_state_regs_1_n7), .SI(
        aes_state_regs_1_S23xDP_6_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_6_ ( .D(aes_state_regs_1_n9), .SI(
        aes_state_regs_1_n6), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_6_ ( .D(aes_state_regs_1_S02xDP_6_), 
        .SI(aes_state_regs_1_S01xDO_6_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n6), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_6_ ( .D(aes_state_regs_1_S01xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_6_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_6_ ( .D(aes_state_regs_1_S21xDP[6]), 
        .SI(aes_state_regs_1_n7), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S01xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_6_ ( .D(aes_state_regs_1_n8), .SI(
        aes_state_regs_1_S30xDP_6_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n7), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_6_ ( .D(aes_state_regs_1_n10), .SI(
        aes_state_regs_1_S02xDP_6_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n8), .QN() );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_6_ ( .D(StateInxD[14]), .SI(
        aes_state_regs_1_n10), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n9), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_6_ ( .D(aes_state_regs_1_S03xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n10), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_6_ ( .D(aes_state_regs_1_S23xDP_6_), 
        .SI(aes_state_regs_1_S20xDP_6_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[6]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_6_ ( .D(aes_state_regs_1_S20xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_6_), .QN(
        aes_state_regs_1_n99) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_5_ ( .D(aes_state_regs_1_S01xDO_5_), 
        .SI(StateInxD[13]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_5_), .QN(aes_state_regs_1_n92) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_5_ ( .D(aes_state_regs_1_n11), .SI(
        aes_state_regs_1_n14), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[5]), .QN(aes_state_regs_1_n49) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_5_ ( .D(aes_state_regs_1_S02xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_5_ ( .D(aes_state_regs_1_n12), .SI(
        aes_state_regs_1_S23xDP_5_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_5_ ( .D(aes_state_regs_1_n14), .SI(
        aes_state_regs_1_n11), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_5_ ( .D(aes_state_regs_1_S02xDP_5_), 
        .SI(aes_state_regs_1_S01xDO_5_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n11), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_5_ ( .D(aes_state_regs_1_S01xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_5_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_5_ ( .D(aes_state_regs_1_S21xDP[5]), 
        .SI(aes_state_regs_1_n12), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_5_ ( .D(aes_state_regs_1_n13), .SI(
        aes_state_regs_1_S30xDP_5_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n12), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_5_ ( .D(aes_state_regs_1_n15), .SI(
        aes_state_regs_1_S02xDP_5_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n13), .QN(aes_state_regs_1_n57) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_5_ ( .D(StateInxD[13]), .SI(
        aes_state_regs_1_n15), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n14), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_5_ ( .D(aes_state_regs_1_S03xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n15), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_5_ ( .D(aes_state_regs_1_S23xDP_5_), 
        .SI(aes_state_regs_1_S20xDP_5_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[5]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_5_ ( .D(aes_state_regs_1_S20xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_5_), .QN(
        aes_state_regs_1_n100) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_4_ ( .D(aes_state_regs_1_S01xDO_4_), 
        .SI(StateInxD[12]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_4_), .QN(aes_state_regs_1_n93) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_4_ ( .D(aes_state_regs_1_n16), .SI(
        aes_state_regs_1_n19), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[4]), .QN(aes_state_regs_1_n50) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_4_ ( .D(aes_state_regs_1_S02xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_4_ ( .D(aes_state_regs_1_n17), .SI(
        aes_state_regs_1_S23xDP_4_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_4_ ( .D(aes_state_regs_1_n19), .SI(
        aes_state_regs_1_n16), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_4_ ( .D(aes_state_regs_1_S02xDP_4_), 
        .SI(aes_state_regs_1_S01xDO_4_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n16), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_4_ ( .D(aes_state_regs_1_S01xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_4_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_4_ ( .D(aes_state_regs_1_S21xDP[4]), 
        .SI(aes_state_regs_1_n17), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_4_ ( .D(aes_state_regs_1_n18), .SI(
        aes_state_regs_1_S30xDP_4_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n17), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_4_ ( .D(aes_state_regs_1_n20), .SI(
        aes_state_regs_1_S02xDP_4_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n18), .QN(aes_state_regs_1_n58) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_4_ ( .D(StateInxD[12]), .SI(
        aes_state_regs_1_n20), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n19), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_4_ ( .D(aes_state_regs_1_S03xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n20), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_4_ ( .D(aes_state_regs_1_S23xDP_4_), 
        .SI(aes_state_regs_1_S20xDP_4_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[4]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_4_ ( .D(aes_state_regs_1_S20xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_4_), .QN(
        aes_state_regs_1_n101) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_3_ ( .D(aes_state_regs_1_S01xDO_3_), 
        .SI(StateInxD[11]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_3_), .QN(aes_state_regs_1_n94) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_3_ ( .D(aes_state_regs_1_n21), .SI(
        aes_state_regs_1_n24), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[3]), .QN(aes_state_regs_1_n51) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_3_ ( .D(aes_state_regs_1_S02xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_3_ ( .D(aes_state_regs_1_n22), .SI(
        aes_state_regs_1_S23xDP_3_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_3_ ( .D(aes_state_regs_1_n24), .SI(
        aes_state_regs_1_n21), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_3_ ( .D(aes_state_regs_1_S02xDP_3_), 
        .SI(aes_state_regs_1_S01xDO_3_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n21), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_3_ ( .D(aes_state_regs_1_S01xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_3_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_3_ ( .D(aes_state_regs_1_S21xDP[3]), 
        .SI(aes_state_regs_1_n22), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_3_ ( .D(aes_state_regs_1_n23), .SI(
        aes_state_regs_1_S30xDP_3_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n22), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_3_ ( .D(aes_state_regs_1_n25), .SI(
        aes_state_regs_1_S02xDP_3_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n23), .QN(aes_state_regs_1_n59) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_3_ ( .D(StateInxD[11]), .SI(
        aes_state_regs_1_n25), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n24), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_3_ ( .D(aes_state_regs_1_S03xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n25), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_3_ ( .D(aes_state_regs_1_S23xDP_3_), 
        .SI(aes_state_regs_1_S20xDP_3_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[3]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_3_ ( .D(aes_state_regs_1_S20xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_3_), .QN(
        aes_state_regs_1_n102) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_2_ ( .D(aes_state_regs_1_S01xDO_2_), 
        .SI(StateInxD[10]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_2_), .QN(aes_state_regs_1_n95) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_2_ ( .D(aes_state_regs_1_n26), .SI(
        aes_state_regs_1_n29), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[2]), .QN(aes_state_regs_1_n52) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_2_ ( .D(aes_state_regs_1_S02xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_2_ ( .D(aes_state_regs_1_n27), .SI(
        aes_state_regs_1_S23xDP_2_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_2_ ( .D(aes_state_regs_1_n29), .SI(
        aes_state_regs_1_n26), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_2_ ( .D(aes_state_regs_1_S02xDP_2_), 
        .SI(aes_state_regs_1_S01xDO_2_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n26), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_2_ ( .D(aes_state_regs_1_S01xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_2_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_2_ ( .D(aes_state_regs_1_S21xDP[2]), 
        .SI(aes_state_regs_1_n27), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_2_ ( .D(aes_state_regs_1_n28), .SI(
        aes_state_regs_1_S30xDP_2_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n27), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_2_ ( .D(aes_state_regs_1_n30), .SI(
        aes_state_regs_1_S02xDP_2_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n28), .QN(aes_state_regs_1_n60) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_2_ ( .D(StateInxD[10]), .SI(
        aes_state_regs_1_n30), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n29), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_2_ ( .D(aes_state_regs_1_S03xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n30), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_2_ ( .D(aes_state_regs_1_S23xDP_2_), 
        .SI(aes_state_regs_1_S20xDP_2_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[2]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_2_ ( .D(aes_state_regs_1_S20xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_2_), .QN(
        aes_state_regs_1_n103) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_1_ ( .D(aes_state_regs_1_S01xDO_1_), 
        .SI(StateInxD[9]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), 
        .Q(aes_state_regs_1_S30xDP_1_), .QN(aes_state_regs_1_n96) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_1_ ( .D(aes_state_regs_1_n31), .SI(
        aes_state_regs_1_n34), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[1]), .QN(aes_state_regs_1_n53) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_1_ ( .D(aes_state_regs_1_S02xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_1_ ( .D(aes_state_regs_1_n32), .SI(
        aes_state_regs_1_S23xDP_1_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_1_ ( .D(aes_state_regs_1_n34), .SI(
        aes_state_regs_1_n31), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_1_ ( .D(aes_state_regs_1_S02xDP_1_), 
        .SI(aes_state_regs_1_S01xDO_1_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n31), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_1_ ( .D(aes_state_regs_1_S01xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_1_ ( .D(aes_state_regs_1_S21xDP[1]), 
        .SI(aes_state_regs_1_n32), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_1_ ( .D(aes_state_regs_1_n33), .SI(
        aes_state_regs_1_S30xDP_1_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n32), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_1_ ( .D(aes_state_regs_1_n35), .SI(
        aes_state_regs_1_S02xDP_1_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n33), .QN(aes_state_regs_1_n61) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_1_ ( .D(StateInxD[9]), .SI(
        aes_state_regs_1_n35), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n34), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_1_ ( .D(aes_state_regs_1_S03xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n35), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_1_ ( .D(aes_state_regs_1_S23xDP_1_), 
        .SI(aes_state_regs_1_S20xDP_1_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[1]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_1_ ( .D(aes_state_regs_1_S20xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_1_), .QN(
        aes_state_regs_1_n104) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_0_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[0]), .SI(aes_state_regs_1_S10xDP_0_), 
        .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[0]), .QN(aes_state_regs_1_n89) );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_0_ ( .D(aes_state_regs_1_S10xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_0_ ( .D(aes_state_regs_1_n37), .SI(
        aes_state_regs_1_S31xDP_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S23xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_0_ ( .D(aes_state_regs_1_S02xDP_0_), 
        .SI(aes_state_regs_1_S01xDO_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S31xDP_0_), .QN() );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_0_ ( .D(aes_state_regs_1_S02xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_0_ ( .D(aes_state_regs_1_S22xDP_0_), 
        .SI(aes_state_regs_1_S23xDP_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_0_ ( .D(aes_state_regs_1_n38), .SI(
        aes_state_regs_1_S30xDP_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S22xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_0_ ( .D(aes_state_regs_1_S01xDO_0_), 
        .SI(StateInxD[8]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), 
        .Q(aes_state_regs_1_S30xDP_0_), .QN(aes_state_regs_1_n97) );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_0_ ( .D(aes_state_regs_1_S01xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_0_ ( .D(aes_state_regs_1_n36), .SI(
        aes_state_regs_1_S22xDP_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_0_ ( .D(aes_state_regs_1_S31xDP_0_), 
        .SI(aes_state_regs_1_n37), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n36), .QN(aes_state_regs_1_n54) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_0_ ( .D(StateInxD[8]), .SI(
        aes_state_regs_1_S03xDP_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n37), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_0_ ( .D(aes_state_regs_1_S03xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_0_ ( .D(aes_state_regs_1_S23xDP_0_), 
        .SI(aes_state_regs_1_S20xDP_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[0]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_0_ ( .D(aes_state_regs_1_S20xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_0_), .QN(
        aes_state_regs_1_n105) );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_0_ ( .D(aes_state_regs_1_S03xDP_0_), 
        .SI(aes_state_regs_1_S02xDP_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n38), .QN(aes_state_regs_1_n62) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U119 ( .A(
        aes_state_regs_1_mix_columns_1_n209), .B(
        aes_state_regs_1_mix_columns_1_n208), .ZN(
        aes_state_regs_1_mix_columns_1_n217) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U118 ( .A(
        aes_state_regs_1_mix_columns_1_n195), .B(
        aes_state_regs_1_mix_columns_1_n233), .ZN(
        aes_state_regs_1_MixColumnsS3xD[0]) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U117 ( .A1(
        aes_state_regs_1_S20xDP_0_), .A2(aes_state_regs_1_mix_columns_1_n232), 
        .B1(aes_state_regs_1_mix_columns_1_n231), .B2(
        aes_state_regs_1_mix_columns_1_n230), .ZN(
        aes_state_regs_1_mix_columns_1_n195) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U116 ( .A(
        aes_state_regs_1_mix_columns_1_n193), .B(
        aes_state_regs_1_mix_columns_1_n194), .ZN(
        aes_state_regs_1_MixColumnsS1xD[2]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U115 ( .A(aes_state_regs_1_S20xDP_1_), .B(aes_state_regs_1_S10xDP_1_), .ZN(aes_state_regs_1_mix_columns_1_n194) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U114 ( .A(
        aes_state_regs_1_mix_columns_1_n215), .B(aes_state_regs_1_S20xDP_2_), 
        .Z(aes_state_regs_1_mix_columns_1_n193) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U113 ( .A(
        aes_state_regs_1_mix_columns_1_n192), .B(
        aes_state_regs_1_mix_columns_1_n217), .ZN(
        aes_state_regs_1_MixColumnsS1xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U112 ( .A(aes_state_regs_1_S20xDP_3_), .B(aes_state_regs_1_mix_columns_1_n206), .ZN(
        aes_state_regs_1_mix_columns_1_n192) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U111 ( .A(
        aes_state_regs_1_mix_columns_1_n190), .B(
        aes_state_regs_1_mix_columns_1_n191), .ZN(
        aes_state_regs_1_MixColumnsS1xD[5]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U110 ( .A(aes_state_regs_1_S20xDP_4_), .B(aes_state_regs_1_S10xDP_4_), .ZN(aes_state_regs_1_mix_columns_1_n191) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U109 ( .A(aes_state_regs_1_S00xDP[5]), 
        .B(aes_state_regs_1_mix_columns_1_n225), .Z(
        aes_state_regs_1_mix_columns_1_n190) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U108 ( .A(
        aes_state_regs_1_mix_columns_1_n189), .B(
        aes_state_regs_1_mix_columns_1_n233), .ZN(
        aes_state_regs_1_MixColumnsS2xD[0]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U107 ( .A(aes_state_regs_1_S20xDP_7_), .B(aes_state_regs_1_mix_columns_1_n213), .ZN(
        aes_state_regs_1_mix_columns_1_n189) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U106 ( .A(
        aes_state_regs_1_mix_columns_1_n187), .B(
        aes_state_regs_1_mix_columns_1_n188), .ZN(
        aes_state_regs_1_MixColumnsS1xD[6]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U105 ( .A(aes_state_regs_1_S20xDP_5_), .B(aes_state_regs_1_S10xDP_5_), .ZN(aes_state_regs_1_mix_columns_1_n188) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U104 ( .A(aes_state_regs_1_S00xDP[6]), 
        .B(aes_state_regs_1_mix_columns_1_n229), .Z(
        aes_state_regs_1_mix_columns_1_n187) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U103 ( .A(
        aes_state_regs_1_mix_columns_1_n186), .B(
        aes_state_regs_1_mix_columns_1_n223), .ZN(
        aes_state_regs_1_mix_columns_1_n210) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U102 ( .A(aes_state_regs_1_S10xDP_7_), .B(aes_state_regs_1_S10xDP_3_), .ZN(aes_state_regs_1_mix_columns_1_n186) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U101 ( .A(
        aes_state_regs_1_mix_columns_1_n185), .B(
        aes_state_regs_1_mix_columns_1_n244), .ZN(
        aes_state_regs_1_MixColumnsS1xD[0]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U100 ( .A(
        aes_state_regs_1_mix_columns_1_n204), .B(aes_state_regs_1_S00xDP[0]), 
        .ZN(aes_state_regs_1_mix_columns_1_n185) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U99 ( .A(
        aes_state_regs_1_mix_columns_1_n183), .B(
        aes_state_regs_1_mix_columns_1_n184), .ZN(
        aes_state_regs_1_MixColumnsS3xD[2]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U98 ( .A(aes_state_regs_1_S30xDP_1_), 
        .B(aes_state_regs_1_S00xDP[2]), .ZN(
        aes_state_regs_1_mix_columns_1_n184) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U97 ( .A(
        aes_state_regs_1_mix_columns_1_n236), .B(aes_state_regs_1_S00xDP[1]), 
        .Z(aes_state_regs_1_mix_columns_1_n183) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U96 ( .A(
        aes_state_regs_1_mix_columns_1_n221), .B(
        aes_state_regs_1_mix_columns_1_n182), .ZN(
        aes_state_regs_1_mix_columns_1_n240) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U95 ( .A1(aes_state_regs_1_S30xDP_3_), .A2(aes_state_regs_1_mix_columns_1_n220), .B1(aes_state_regs_1_S30xDP_7_), 
        .B2(aes_state_regs_1_mix_columns_1_n181), .ZN(
        aes_state_regs_1_mix_columns_1_n182) );
  INV_X1 aes_state_regs_1_mix_columns_1_U94 ( .A(aes_state_regs_1_S30xDP_3_), 
        .ZN(aes_state_regs_1_mix_columns_1_n181) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U93 ( .A(
        aes_state_regs_1_mix_columns_1_n180), .B(
        aes_state_regs_1_mix_columns_1_n179), .ZN(
        aes_state_regs_1_MixColumnsS3xD[6]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U92 ( .A(aes_state_regs_1_S30xDP_5_), 
        .B(aes_state_regs_1_S00xDP[5]), .ZN(
        aes_state_regs_1_mix_columns_1_n180) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U91 ( .A1(
        aes_state_regs_1_mix_columns_1_n243), .A2(aes_state_regs_1_S20xDP_6_), 
        .B1(aes_state_regs_1_mix_columns_1_n242), .B2(
        aes_state_regs_1_mix_columns_1_n178), .ZN(
        aes_state_regs_1_mix_columns_1_n179) );
  INV_X1 aes_state_regs_1_mix_columns_1_U90 ( .A(
        aes_state_regs_1_mix_columns_1_n243), .ZN(
        aes_state_regs_1_mix_columns_1_n178) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U89 ( .A(
        aes_state_regs_1_mix_columns_1_n177), .B(
        aes_state_regs_1_mix_columns_1_n212), .ZN(
        aes_state_regs_1_MixColumnsS1xD[1]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U88 ( .A(
        aes_state_regs_1_mix_columns_1_n205), .B(aes_state_regs_1_S00xDP[1]), 
        .ZN(aes_state_regs_1_mix_columns_1_n177) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U87 ( .A1(aes_state_regs_1_S30xDP_2_), .A2(aes_state_regs_1_S30xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n220), 
        .B2(aes_state_regs_1_mix_columns_1_n176), .ZN(
        aes_state_regs_1_mix_columns_1_n238) );
  INV_X1 aes_state_regs_1_mix_columns_1_U86 ( .A(aes_state_regs_1_S30xDP_2_), 
        .ZN(aes_state_regs_1_mix_columns_1_n176) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U85 ( .A(
        aes_state_regs_1_mix_columns_1_n175), .B(
        aes_state_regs_1_mix_columns_1_n235), .ZN(
        aes_state_regs_1_MixColumnsS3xD[1]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U84 ( .A(
        aes_state_regs_1_mix_columns_1_n234), .B(aes_state_regs_1_S20xDP_1_), 
        .ZN(aes_state_regs_1_mix_columns_1_n175) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U83 ( .A(
        aes_state_regs_1_mix_columns_1_n174), .B(
        aes_state_regs_1_mix_columns_1_n219), .ZN(
        aes_state_regs_1_MixColumnsS1xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U82 ( .A(
        aes_state_regs_1_mix_columns_1_n210), .B(aes_state_regs_1_S00xDP[4]), 
        .ZN(aes_state_regs_1_mix_columns_1_n174) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U81 ( .A(
        aes_state_regs_1_mix_columns_1_n173), .B(
        aes_state_regs_1_mix_columns_1_n238), .ZN(
        aes_state_regs_1_MixColumnsS3xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U80 ( .A(
        aes_state_regs_1_mix_columns_1_n237), .B(aes_state_regs_1_S00xDP[3]), 
        .ZN(aes_state_regs_1_mix_columns_1_n173) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U79 ( .A(
        aes_state_regs_1_mix_columns_1_n172), .B(
        aes_state_regs_1_mix_columns_1_n205), .ZN(
        aes_state_regs_1_MixColumnsS0xD[1]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U78 ( .A(aes_state_regs_1_S10xDP_1_), 
        .B(aes_state_regs_1_mix_columns_1_n234), .ZN(
        aes_state_regs_1_mix_columns_1_n172) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U77 ( .A(
        aes_state_regs_1_mix_columns_1_n171), .B(
        aes_state_regs_1_mix_columns_1_n240), .ZN(
        aes_state_regs_1_MixColumnsS3xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U76 ( .A(
        aes_state_regs_1_mix_columns_1_n239), .B(aes_state_regs_1_S20xDP_4_), 
        .ZN(aes_state_regs_1_mix_columns_1_n171) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U75 ( .A1(aes_state_regs_1_S20xDP_3_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n211), 
        .B2(aes_state_regs_1_mix_columns_1_n170), .ZN(
        aes_state_regs_1_mix_columns_1_n219) );
  INV_X1 aes_state_regs_1_mix_columns_1_U74 ( .A(aes_state_regs_1_S20xDP_3_), 
        .ZN(aes_state_regs_1_mix_columns_1_n170) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U73 ( .A(
        aes_state_regs_1_mix_columns_1_n168), .B(
        aes_state_regs_1_mix_columns_1_n169), .ZN(
        aes_state_regs_1_MixColumnsS3xD[5]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U72 ( .A(
        aes_state_regs_1_mix_columns_1_n241), .B(aes_state_regs_1_S20xDP_5_), 
        .ZN(aes_state_regs_1_mix_columns_1_n169) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U71 ( .A(aes_state_regs_1_S00xDP[4]), 
        .B(aes_state_regs_1_S30xDP_4_), .Z(aes_state_regs_1_mix_columns_1_n168) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U70 ( .A(
        aes_state_regs_1_mix_columns_1_n166), .B(
        aes_state_regs_1_mix_columns_1_n167), .ZN(
        aes_state_regs_1_MixColumnsS1xD[7]) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U69 ( .A1(aes_state_regs_1_S20xDP_6_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n211), 
        .B2(aes_state_regs_1_mix_columns_1_n242), .ZN(
        aes_state_regs_1_mix_columns_1_n167) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U68 ( .A(aes_state_regs_1_S10xDP_6_), 
        .B(aes_state_regs_1_mix_columns_1_n231), .ZN(
        aes_state_regs_1_mix_columns_1_n166) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U67 ( .A(
        aes_state_regs_1_mix_columns_1_n165), .B(
        aes_state_regs_1_mix_columns_1_n164), .ZN(
        aes_state_regs_1_MixColumnsS3xD[7]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U66 ( .A(
        aes_state_regs_1_mix_columns_1_n244), .B(aes_state_regs_1_S30xDP_6_), 
        .ZN(aes_state_regs_1_mix_columns_1_n165) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U65 ( .A1(aes_state_regs_1_S00xDP[6]), .A2(aes_state_regs_1_S00xDP[7]), .B1(aes_state_regs_1_mix_columns_1_n245), 
        .B2(aes_state_regs_1_mix_columns_1_n163), .ZN(
        aes_state_regs_1_mix_columns_1_n164) );
  INV_X1 aes_state_regs_1_mix_columns_1_U64 ( .A(aes_state_regs_1_S00xDP[6]), 
        .ZN(aes_state_regs_1_mix_columns_1_n163) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U63 ( .A(
        aes_state_regs_1_mix_columns_1_n162), .B(
        aes_state_regs_1_mix_columns_1_n235), .ZN(
        aes_state_regs_1_MixColumnsS2xD[1]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U62 ( .A(aes_state_regs_1_S30xDP_1_), 
        .B(aes_state_regs_1_mix_columns_1_n212), .ZN(
        aes_state_regs_1_mix_columns_1_n162) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U61 ( .A(
        aes_state_regs_1_mix_columns_1_n160), .B(
        aes_state_regs_1_mix_columns_1_n161), .ZN(
        aes_state_regs_1_mix_columns_1_n237) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U60 ( .A(aes_state_regs_1_S20xDP_3_), 
        .B(aes_state_regs_1_S00xDP[7]), .ZN(
        aes_state_regs_1_mix_columns_1_n161) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U59 ( .A(aes_state_regs_1_S00xDP[2]), 
        .B(aes_state_regs_1_S10xDP_3_), .Z(aes_state_regs_1_mix_columns_1_n160) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U58 ( .A(
        aes_state_regs_1_mix_columns_1_n215), .B(
        aes_state_regs_1_mix_columns_1_n159), .ZN(
        aes_state_regs_1_MixColumnsS2xD[2]) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U57 ( .A(
        aes_state_regs_1_mix_columns_1_n216), .B(aes_state_regs_1_S10xDP_2_), 
        .Z(aes_state_regs_1_mix_columns_1_n159) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U56 ( .A(aes_state_regs_1_S10xDP_3_), 
        .B(aes_state_regs_1_mix_columns_1_n217), .ZN(
        aes_state_regs_1_mix_columns_1_n218) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U55 ( .A(
        aes_state_regs_1_mix_columns_1_n218), .B(
        aes_state_regs_1_mix_columns_1_n238), .ZN(
        aes_state_regs_1_MixColumnsS2xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U54 ( .A(aes_state_regs_1_S30xDP_4_), 
        .B(aes_state_regs_1_mix_columns_1_n219), .ZN(
        aes_state_regs_1_mix_columns_1_n222) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U53 ( .A(
        aes_state_regs_1_mix_columns_1_n222), .B(
        aes_state_regs_1_mix_columns_1_n240), .ZN(
        aes_state_regs_1_MixColumnsS2xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U52 ( .A(
        aes_state_regs_1_mix_columns_1_n223), .B(aes_state_regs_1_S30xDP_5_), 
        .ZN(aes_state_regs_1_mix_columns_1_n224) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U51 ( .A(
        aes_state_regs_1_mix_columns_1_n224), .B(
        aes_state_regs_1_mix_columns_1_n241), .ZN(
        aes_state_regs_1_MixColumnsS2xD[5]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U50 ( .A(
        aes_state_regs_1_mix_columns_1_n225), .B(aes_state_regs_1_S30xDP_6_), 
        .ZN(aes_state_regs_1_mix_columns_1_n226) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U49 ( .A(
        aes_state_regs_1_mix_columns_1_n226), .B(
        aes_state_regs_1_mix_columns_1_n243), .ZN(
        aes_state_regs_1_MixColumnsS2xD[6]) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U48 ( .A1(aes_state_regs_1_S10xDP_7_), .A2(aes_state_regs_1_mix_columns_1_n232), .B1(
        aes_state_regs_1_mix_columns_1_n231), .B2(
        aes_state_regs_1_mix_columns_1_n227), .ZN(
        aes_state_regs_1_mix_columns_1_n228) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U47 ( .A(
        aes_state_regs_1_mix_columns_1_n229), .B(
        aes_state_regs_1_mix_columns_1_n228), .ZN(
        aes_state_regs_1_MixColumnsS2xD[7]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U46 ( .A(
        aes_state_regs_1_mix_columns_1_n244), .B(
        aes_state_regs_1_mix_columns_1_n243), .ZN(
        aes_state_regs_1_mix_columns_1_n203) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U45 ( .A(
        aes_state_regs_1_mix_columns_1_n203), .B(aes_state_regs_1_S30xDP_7_), 
        .ZN(aes_state_regs_1_MixColumnsS0xD[7]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U44 ( .A(aes_state_regs_1_S10xDP_4_), 
        .B(aes_state_regs_1_mix_columns_1_n239), .ZN(
        aes_state_regs_1_mix_columns_1_n200) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U43 ( .A(
        aes_state_regs_1_mix_columns_1_n200), .B(
        aes_state_regs_1_mix_columns_1_n210), .ZN(
        aes_state_regs_1_MixColumnsS0xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U42 ( .A(aes_state_regs_1_S30xDP_3_), 
        .B(aes_state_regs_1_mix_columns_1_n237), .ZN(
        aes_state_regs_1_mix_columns_1_n199) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U41 ( .A(
        aes_state_regs_1_mix_columns_1_n199), .B(
        aes_state_regs_1_mix_columns_1_n206), .ZN(
        aes_state_regs_1_MixColumnsS0xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U40 ( .A(aes_state_regs_1_S30xDP_2_), 
        .B(aes_state_regs_1_mix_columns_1_n236), .ZN(
        aes_state_regs_1_mix_columns_1_n198) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U39 ( .A(
        aes_state_regs_1_mix_columns_1_n198), .B(
        aes_state_regs_1_mix_columns_1_n214), .ZN(
        aes_state_regs_1_MixColumnsS0xD[2]) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U38 ( .A(aes_state_regs_1_S10xDP_0_), 
        .B(aes_state_regs_1_S00xDP[0]), .Z(aes_state_regs_1_mix_columns_1_n233) );
  INV_X1 aes_state_regs_1_mix_columns_1_U37 ( .A(
        aes_state_regs_1_mix_columns_1_n231), .ZN(
        aes_state_regs_1_mix_columns_1_n232) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U36 ( .A1(aes_state_regs_1_S00xDP[7]), .A2(aes_state_regs_1_S30xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n220), 
        .B2(aes_state_regs_1_mix_columns_1_n245), .ZN(
        aes_state_regs_1_mix_columns_1_n231) );
  INV_X1 aes_state_regs_1_mix_columns_1_U35 ( .A(aes_state_regs_1_S20xDP_0_), 
        .ZN(aes_state_regs_1_mix_columns_1_n230) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U34 ( .A(aes_state_regs_1_S30xDP_0_), 
        .B(aes_state_regs_1_mix_columns_1_n220), .ZN(
        aes_state_regs_1_mix_columns_1_n213) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U33 ( .A(aes_state_regs_1_S30xDP_0_), 
        .B(aes_state_regs_1_S20xDP_0_), .Z(aes_state_regs_1_mix_columns_1_n204) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U32 ( .A1(aes_state_regs_1_S10xDP_7_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n211), 
        .B2(aes_state_regs_1_mix_columns_1_n227), .ZN(
        aes_state_regs_1_mix_columns_1_n244) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U31 ( .A(
        aes_state_regs_1_mix_columns_1_n214), .B(
        aes_state_regs_1_mix_columns_1_n213), .Z(
        aes_state_regs_1_mix_columns_1_n235) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U30 ( .A(aes_state_regs_1_S00xDP[7]), 
        .B(aes_state_regs_1_S00xDP[0]), .Z(aes_state_regs_1_mix_columns_1_n234) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U29 ( .A(aes_state_regs_1_S10xDP_2_), 
        .B(aes_state_regs_1_S20xDP_2_), .Z(aes_state_regs_1_mix_columns_1_n236) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U28 ( .A(aes_state_regs_1_S00xDP[7]), 
        .B(aes_state_regs_1_S00xDP[3]), .Z(aes_state_regs_1_mix_columns_1_n239) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U27 ( .A(aes_state_regs_1_S10xDP_5_), 
        .B(aes_state_regs_1_S00xDP[5]), .Z(aes_state_regs_1_mix_columns_1_n241) );
  INV_X1 aes_state_regs_1_mix_columns_1_U26 ( .A(aes_state_regs_1_S20xDP_6_), 
        .ZN(aes_state_regs_1_mix_columns_1_n242) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U25 ( .A(aes_state_regs_1_S10xDP_6_), 
        .B(aes_state_regs_1_S00xDP[6]), .Z(aes_state_regs_1_mix_columns_1_n243) );
  INV_X1 aes_state_regs_1_mix_columns_1_U24 ( .A(aes_state_regs_1_S00xDP[7]), 
        .ZN(aes_state_regs_1_mix_columns_1_n245) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U23 ( .A1(aes_state_regs_1_S20xDP_0_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n211), 
        .B2(aes_state_regs_1_mix_columns_1_n230), .ZN(
        aes_state_regs_1_mix_columns_1_n212) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U22 ( .A(aes_state_regs_1_S30xDP_2_), 
        .B(aes_state_regs_1_S00xDP[2]), .Z(aes_state_regs_1_mix_columns_1_n215) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U21 ( .A(aes_state_regs_1_S30xDP_1_), 
        .B(aes_state_regs_1_S20xDP_1_), .ZN(
        aes_state_regs_1_mix_columns_1_n216) );
  INV_X1 aes_state_regs_1_mix_columns_1_U20 ( .A(aes_state_regs_1_S00xDP[3]), 
        .ZN(aes_state_regs_1_mix_columns_1_n207) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U19 ( .A1(aes_state_regs_1_S00xDP[3]), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n211), 
        .B2(aes_state_regs_1_mix_columns_1_n207), .ZN(
        aes_state_regs_1_mix_columns_1_n208) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U18 ( .A(aes_state_regs_1_S20xDP_2_), 
        .B(aes_state_regs_1_S30xDP_3_), .ZN(
        aes_state_regs_1_mix_columns_1_n209) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U17 ( .A(aes_state_regs_1_S30xDP_4_), 
        .B(aes_state_regs_1_S20xDP_4_), .Z(aes_state_regs_1_mix_columns_1_n223) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U16 ( .A(aes_state_regs_1_S30xDP_5_), 
        .B(aes_state_regs_1_S20xDP_5_), .Z(aes_state_regs_1_mix_columns_1_n225) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U15 ( .A(aes_state_regs_1_S30xDP_6_), 
        .B(aes_state_regs_1_S20xDP_6_), .Z(aes_state_regs_1_mix_columns_1_n229) );
  INV_X1 aes_state_regs_1_mix_columns_1_U14 ( .A(aes_state_regs_1_S10xDP_7_), 
        .ZN(aes_state_regs_1_mix_columns_1_n227) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U13 ( .A(
        aes_state_regs_1_mix_columns_1_n197), .B(
        aes_state_regs_1_mix_columns_1_n216), .ZN(
        aes_state_regs_1_mix_columns_1_n205) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U12 ( .A(aes_state_regs_1_S10xDP_7_), 
        .B(aes_state_regs_1_S10xDP_2_), .Z(aes_state_regs_1_mix_columns_1_n206) );
  INV_X1 aes_state_regs_1_mix_columns_1_U11 ( .A(aes_state_regs_1_S20xDP_7_), 
        .ZN(aes_state_regs_1_mix_columns_1_n211) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U10 ( .A(aes_state_regs_1_S00xDP[7]), 
        .B(aes_state_regs_1_mix_columns_1_n197), .ZN(
        aes_state_regs_1_mix_columns_1_n196) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U9 ( .A(
        aes_state_regs_1_mix_columns_1_n196), .B(
        aes_state_regs_1_mix_columns_1_n204), .ZN(
        aes_state_regs_1_MixColumnsS0xD[0]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U8 ( .A(aes_state_regs_1_S10xDP_6_), 
        .B(aes_state_regs_1_mix_columns_1_n241), .ZN(
        aes_state_regs_1_mix_columns_1_n202) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U7 ( .A(
        aes_state_regs_1_mix_columns_1_n202), .B(
        aes_state_regs_1_mix_columns_1_n229), .ZN(
        aes_state_regs_1_MixColumnsS0xD[6]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U6 ( .A(aes_state_regs_1_S10xDP_5_), 
        .B(aes_state_regs_1_mix_columns_1_n221), .ZN(
        aes_state_regs_1_mix_columns_1_n201) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U5 ( .A(
        aes_state_regs_1_mix_columns_1_n201), .B(
        aes_state_regs_1_mix_columns_1_n225), .ZN(
        aes_state_regs_1_MixColumnsS0xD[5]) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U4 ( .A(aes_state_regs_1_S10xDP_1_), 
        .B(aes_state_regs_1_S00xDP[1]), .Z(aes_state_regs_1_mix_columns_1_n214) );
  INV_X1 aes_state_regs_1_mix_columns_1_U3 ( .A(aes_state_regs_1_S30xDP_7_), 
        .ZN(aes_state_regs_1_mix_columns_1_n220) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U2 ( .A(aes_state_regs_1_S10xDP_4_), 
        .B(aes_state_regs_1_S00xDP[4]), .Z(aes_state_regs_1_mix_columns_1_n221) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U1 ( .A(aes_state_regs_1_S10xDP_7_), 
        .B(aes_state_regs_1_S10xDP_0_), .Z(aes_state_regs_1_mix_columns_1_n197) );
  BUF_X1 aes_key_regs_0_U3 ( .A(n114), .Z(aes_key_regs_0_n4) );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_0_ ( .D(aes_key_regs_0_K00xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_0_ ( .D(aes_key_regs_0_K10xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_0_ ( .D(aes_key_regs_0_K20xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_0_ ( .D(aes_key_regs_0_K01xDP_0_), .SI(
        KeyOutxD[0]), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K20xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_0_ ( .D(aes_key_regs_0_K01xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_0_ ( .D(aes_key_regs_0_K11xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_0_ ( .D(aes_key_regs_0_K21xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_0_ ( .D(aes_key_regs_0_K02xDP_0_), .SI(
        aes_key_regs_0_K01xDP_0_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K21xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_0_ ( .D(aes_key_regs_0_K02xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_0_ ( .D(aes_key_regs_0_K12xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_0_ ( .D(aes_key_regs_0_K22xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_0_ ( .D(K03xD[0]), .SI(
        aes_key_regs_0_K02xDP_0_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_1_ ( .D(aes_key_regs_0_K00xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_1_ ( .D(aes_key_regs_0_K10xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_1_ ( .D(aes_key_regs_0_K20xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_1_ ( .D(aes_key_regs_0_K01xDP_1_), .SI(
        KeyOutxD[1]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_1_ ( .D(aes_key_regs_0_K01xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_1_ ( .D(aes_key_regs_0_K11xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_1_ ( .D(aes_key_regs_0_K21xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_1_ ( .D(aes_key_regs_0_K02xDP_1_), .SI(
        aes_key_regs_0_K01xDP_1_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_1_ ( .D(aes_key_regs_0_K02xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_1_ ( .D(aes_key_regs_0_K12xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_1_ ( .D(aes_key_regs_0_K22xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_1_ ( .D(K03xD[1]), .SI(
        aes_key_regs_0_K02xDP_1_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_2_ ( .D(aes_key_regs_0_K00xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_2_ ( .D(aes_key_regs_0_K10xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_2_ ( .D(aes_key_regs_0_K20xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_2_ ( .D(aes_key_regs_0_K01xDP_2_), .SI(
        KeyOutxD[2]), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K20xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_2_ ( .D(aes_key_regs_0_K01xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_2_ ( .D(aes_key_regs_0_K11xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_2_ ( .D(aes_key_regs_0_K21xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_2_ ( .D(aes_key_regs_0_K02xDP_2_), .SI(
        aes_key_regs_0_K01xDP_2_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_2_ ( .D(aes_key_regs_0_K02xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_2_ ( .D(aes_key_regs_0_K12xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_2_ ( .D(aes_key_regs_0_K22xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_2_ ( .D(K03xD[2]), .SI(
        aes_key_regs_0_K02xDP_2_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_3_ ( .D(aes_key_regs_0_K00xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_3_ ( .D(aes_key_regs_0_K10xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_3_ ( .D(aes_key_regs_0_K20xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_3_ ( .D(aes_key_regs_0_K01xDP_3_), .SI(
        KeyOutxD[3]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_3_ ( .D(aes_key_regs_0_K01xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_3_ ( .D(aes_key_regs_0_K11xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_3_ ( .D(aes_key_regs_0_K21xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_3_ ( .D(aes_key_regs_0_K02xDP_3_), .SI(
        aes_key_regs_0_K01xDP_3_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_3_ ( .D(aes_key_regs_0_K02xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_3_ ( .D(aes_key_regs_0_K12xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_3_ ( .D(aes_key_regs_0_K22xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_3_ ( .D(K03xD[3]), .SI(
        aes_key_regs_0_K02xDP_3_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_4_ ( .D(aes_key_regs_0_K00xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_4_ ( .D(aes_key_regs_0_K10xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_4_ ( .D(aes_key_regs_0_K20xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_4_ ( .D(aes_key_regs_0_K01xDP_4_), .SI(
        KeyOutxD[4]), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K20xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_4_ ( .D(aes_key_regs_0_K01xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_4_ ( .D(aes_key_regs_0_K11xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_4_ ( .D(aes_key_regs_0_K21xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_4_ ( .D(aes_key_regs_0_K02xDP_4_), .SI(
        aes_key_regs_0_K01xDP_4_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K21xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_4_ ( .D(aes_key_regs_0_K02xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_4_ ( .D(aes_key_regs_0_K12xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_4_ ( .D(aes_key_regs_0_K22xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_4_ ( .D(K03xD[4]), .SI(
        aes_key_regs_0_K02xDP_4_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K22xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_5_ ( .D(aes_key_regs_0_K00xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_5_ ( .D(aes_key_regs_0_K10xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_5_ ( .D(aes_key_regs_0_K20xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_5_ ( .D(aes_key_regs_0_K01xDP_5_), .SI(
        KeyOutxD[5]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_5_ ( .D(aes_key_regs_0_K01xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_5_ ( .D(aes_key_regs_0_K11xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_5_ ( .D(aes_key_regs_0_K21xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_5_ ( .D(aes_key_regs_0_K02xDP_5_), .SI(
        aes_key_regs_0_K01xDP_5_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_5_ ( .D(aes_key_regs_0_K02xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_5_ ( .D(aes_key_regs_0_K12xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_5_ ( .D(aes_key_regs_0_K22xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_5_ ( .D(K03xD[5]), .SI(
        aes_key_regs_0_K02xDP_5_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_6_ ( .D(aes_key_regs_0_K00xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_6_ ( .D(aes_key_regs_0_K10xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_6_ ( .D(aes_key_regs_0_K20xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_6_ ( .D(aes_key_regs_0_K01xDP_6_), .SI(
        KeyOutxD[6]), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K20xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_6_ ( .D(aes_key_regs_0_K01xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_6_ ( .D(aes_key_regs_0_K11xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_6_ ( .D(aes_key_regs_0_K21xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_6_ ( .D(aes_key_regs_0_K02xDP_6_), .SI(
        aes_key_regs_0_K01xDP_6_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K21xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_6_ ( .D(aes_key_regs_0_K02xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_6_ ( .D(aes_key_regs_0_K12xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_6_ ( .D(aes_key_regs_0_K22xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_6_ ( .D(K03xD[6]), .SI(
        aes_key_regs_0_K02xDP_6_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K22xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_7_ ( .D(aes_key_regs_0_K00xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_7_ ( .D(aes_key_regs_0_K10xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_7_ ( .D(aes_key_regs_0_K20xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_7_ ( .D(aes_key_regs_0_K01xDP_7_), .SI(
        KeyOutxD[7]), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K20xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_7_ ( .D(aes_key_regs_0_K01xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_7_ ( .D(aes_key_regs_0_K11xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_7_ ( .D(aes_key_regs_0_K21xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_7_ ( .D(aes_key_regs_0_K02xDP_7_), .SI(
        aes_key_regs_0_K01xDP_7_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K21xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_7_ ( .D(aes_key_regs_0_K02xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_7_ ( .D(aes_key_regs_0_K12xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_7_ ( .D(aes_key_regs_0_K22xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_7_ ( .D(K03xD[7]), .SI(
        aes_key_regs_0_K02xDP_7_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K22xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_0_ ( .D(KeyInxD[0]), .SI(K03xD[0]), .SE(
        n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[0]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_0_ ( .D(KeyToSboxOutxD[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_0_ ( .D(aes_key_regs_0_K13xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_0_ ( .D(aes_key_regs_0_K23xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_1_ ( .D(KeyInxD[1]), .SI(K03xD[1]), .SE(
        n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[1]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_1_ ( .D(KeyToSboxOutxD[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_1_ ( .D(aes_key_regs_0_K13xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_1_ ( .D(aes_key_regs_0_K23xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_2_ ( .D(KeyInxD[2]), .SI(K03xD[2]), .SE(
        n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[2]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_2_ ( .D(KeyToSboxOutxD[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_2_ ( .D(aes_key_regs_0_K13xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_2_ ( .D(aes_key_regs_0_K23xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_3_ ( .D(KeyInxD[3]), .SI(K03xD[3]), .SE(
        n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[3]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_3_ ( .D(KeyToSboxOutxD[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_3_ ( .D(aes_key_regs_0_K13xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_3_ ( .D(aes_key_regs_0_K23xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_4_ ( .D(KeyInxD[4]), .SI(K03xD[4]), .SE(
        n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[4]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_4_ ( .D(KeyToSboxOutxD[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_4_ ( .D(aes_key_regs_0_K13xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_4_ ( .D(aes_key_regs_0_K23xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_5_ ( .D(KeyInxD[5]), .SI(K03xD[5]), .SE(
        n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[5]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_5_ ( .D(KeyToSboxOutxD[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_5_ ( .D(aes_key_regs_0_K13xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_5_ ( .D(aes_key_regs_0_K23xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_6_ ( .D(KeyInxD[6]), .SI(K03xD[6]), .SE(
        n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[6]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_6_ ( .D(KeyToSboxOutxD[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_6_ ( .D(aes_key_regs_0_K13xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_6_ ( .D(aes_key_regs_0_K23xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_7_ ( .D(KeyInxD[7]), .SI(K03xD[7]), .SE(
        n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[7]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_7_ ( .D(KeyToSboxOutxD[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_7_ ( .D(aes_key_regs_0_K13xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_7_ ( .D(aes_key_regs_0_K23xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[7]), .QN() );
  INV_X1 aes_state_regs_0_U56 ( .A(aes_state_regs_0_MixColumnsS2xD[7]), .ZN(
        aes_state_regs_0_n186) );
  INV_X1 aes_state_regs_0_U55 ( .A(aes_state_regs_0_MixColumnsS2xD[6]), .ZN(
        aes_state_regs_0_n185) );
  INV_X1 aes_state_regs_0_U54 ( .A(aes_state_regs_0_MixColumnsS2xD[5]), .ZN(
        aes_state_regs_0_n184) );
  INV_X1 aes_state_regs_0_U53 ( .A(aes_state_regs_0_MixColumnsS2xD[4]), .ZN(
        aes_state_regs_0_n183) );
  INV_X1 aes_state_regs_0_U52 ( .A(aes_state_regs_0_MixColumnsS2xD[3]), .ZN(
        aes_state_regs_0_n182) );
  INV_X1 aes_state_regs_0_U51 ( .A(aes_state_regs_0_MixColumnsS2xD[2]), .ZN(
        aes_state_regs_0_n181) );
  INV_X1 aes_state_regs_0_U50 ( .A(aes_state_regs_0_MixColumnsS2xD[1]), .ZN(
        aes_state_regs_0_n180) );
  INV_X2 aes_state_regs_0_U49 ( .A(aes_state_regs_0_n178), .ZN(
        aes_state_regs_0_n177) );
  INV_X4 aes_state_regs_0_U48 ( .A(aes_state_regs_0_n178), .ZN(
        aes_state_regs_0_n176) );
  INV_X1 aes_state_regs_0_U47 ( .A(nextRCONxS), .ZN(aes_state_regs_0_n178) );
  OAI21_X1 aes_state_regs_0_U46 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n34), .A(aes_state_regs_0_n175), .ZN(StateOutxD[6])
         );
  NAND2_X1 aes_state_regs_0_U45 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[6]), .ZN(aes_state_regs_0_n175) );
  OAI21_X1 aes_state_regs_0_U44 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n33), .A(aes_state_regs_0_n174), .ZN(StateOutxD[5])
         );
  NAND2_X1 aes_state_regs_0_U43 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[5]), .ZN(aes_state_regs_0_n174) );
  AOI22_X1 aes_state_regs_0_U42 ( .A1(aes_state_regs_0_n177), .A2(
        aes_state_regs_0_n136), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[0]), .ZN(aes_state_regs_0_n187) );
  OAI21_X1 aes_state_regs_0_U41 ( .B1(aes_state_regs_0_n43), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n187), .ZN(
        aes_state_regs_0_S20xDN[0]) );
  AOI22_X1 aes_state_regs_0_U40 ( .A1(aes_state_regs_0_n177), .A2(
        aes_state_regs_0_n138), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS2xD[0]), .ZN(aes_state_regs_0_n179) );
  OAI21_X1 aes_state_regs_0_U39 ( .B1(aes_state_regs_0_n51), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n179), .ZN(
        aes_state_regs_0_S10xDN[0]) );
  NAND2_X2 aes_state_regs_0_U38 ( .A1(doMixColumnsxS), .A2(
        aes_state_regs_0_n178), .ZN(aes_state_regs_0_n109) );
  AOI22_X1 aes_state_regs_0_U37 ( .A1(aes_state_regs_0_n177), .A2(
        aes_state_regs_0_n141), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[1]), .ZN(aes_state_regs_0_n188) );
  OAI21_X1 aes_state_regs_0_U36 ( .B1(aes_state_regs_0_n42), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n188), .ZN(
        aes_state_regs_0_S20xDN[1]) );
  AOI22_X1 aes_state_regs_0_U35 ( .A1(aes_state_regs_0_n177), .A2(
        aes_state_regs_0_n146), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[2]), .ZN(aes_state_regs_0_n189) );
  OAI21_X1 aes_state_regs_0_U34 ( .B1(aes_state_regs_0_n41), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n189), .ZN(
        aes_state_regs_0_S20xDN[2]) );
  AOI22_X1 aes_state_regs_0_U33 ( .A1(aes_state_regs_0_n177), .A2(
        aes_state_regs_0_n151), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[3]), .ZN(aes_state_regs_0_n190) );
  OAI21_X1 aes_state_regs_0_U32 ( .B1(aes_state_regs_0_n40), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n190), .ZN(
        aes_state_regs_0_S20xDN[3]) );
  AOI22_X1 aes_state_regs_0_U31 ( .A1(aes_state_regs_0_n176), .A2(
        aes_state_regs_0_n156), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[4]), .ZN(aes_state_regs_0_n191) );
  OAI21_X1 aes_state_regs_0_U30 ( .B1(aes_state_regs_0_n39), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n191), .ZN(
        aes_state_regs_0_S20xDN[4]) );
  AOI22_X1 aes_state_regs_0_U29 ( .A1(aes_state_regs_0_n176), .A2(
        aes_state_regs_0_n161), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[5]), .ZN(aes_state_regs_0_n192) );
  OAI21_X1 aes_state_regs_0_U28 ( .B1(aes_state_regs_0_n38), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n192), .ZN(
        aes_state_regs_0_S20xDN[5]) );
  AOI22_X1 aes_state_regs_0_U27 ( .A1(aes_state_regs_0_n176), .A2(
        aes_state_regs_0_n166), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[6]), .ZN(aes_state_regs_0_n193) );
  OAI21_X1 aes_state_regs_0_U26 ( .B1(aes_state_regs_0_n37), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n193), .ZN(
        aes_state_regs_0_S20xDN[6]) );
  AOI22_X1 aes_state_regs_0_U25 ( .A1(aes_state_regs_0_n176), .A2(
        aes_state_regs_0_n171), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[7]), .ZN(aes_state_regs_0_n194) );
  OAI21_X1 aes_state_regs_0_U24 ( .B1(aes_state_regs_0_n36), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n194), .ZN(
        aes_state_regs_0_S20xDN[7]) );
  OAI222_X1 aes_state_regs_0_U23 ( .A1(aes_state_regs_0_n180), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n50), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n121), .ZN(aes_state_regs_0_S10xDN[1]) );
  OAI222_X1 aes_state_regs_0_U22 ( .A1(aes_state_regs_0_n181), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n49), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n122), .ZN(aes_state_regs_0_S10xDN[2]) );
  OAI222_X1 aes_state_regs_0_U21 ( .A1(aes_state_regs_0_n182), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n48), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n123), .ZN(aes_state_regs_0_S10xDN[3]) );
  OAI222_X1 aes_state_regs_0_U20 ( .A1(aes_state_regs_0_n183), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n47), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n124), .ZN(aes_state_regs_0_S10xDN[4]) );
  OAI222_X1 aes_state_regs_0_U19 ( .A1(aes_state_regs_0_n184), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n46), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n125), .ZN(aes_state_regs_0_S10xDN[5]) );
  OAI222_X1 aes_state_regs_0_U18 ( .A1(aes_state_regs_0_n185), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n45), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n126), .ZN(aes_state_regs_0_S10xDN[6]) );
  OAI222_X1 aes_state_regs_0_U17 ( .A1(aes_state_regs_0_n186), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n44), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n127), .ZN(aes_state_regs_0_S10xDN[7]) );
  NAND2_X1 aes_state_regs_0_U16 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[0]), .ZN(aes_state_regs_0_n201) );
  OAI21_X1 aes_state_regs_0_U15 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n35), .A(aes_state_regs_0_n201), .ZN(StateOutxD[0])
         );
  NAND2_X1 aes_state_regs_0_U14 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[7]), .ZN(aes_state_regs_0_n196) );
  OAI21_X1 aes_state_regs_0_U13 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n28), .A(aes_state_regs_0_n196), .ZN(StateOutxD[7])
         );
  NAND2_X1 aes_state_regs_0_U12 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[4]), .ZN(aes_state_regs_0_n197) );
  OAI21_X1 aes_state_regs_0_U11 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n32), .A(aes_state_regs_0_n197), .ZN(StateOutxD[4])
         );
  NAND2_X1 aes_state_regs_0_U10 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[3]), .ZN(aes_state_regs_0_n198) );
  OAI21_X1 aes_state_regs_0_U9 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n31), .A(aes_state_regs_0_n198), .ZN(StateOutxD[3])
         );
  NAND2_X1 aes_state_regs_0_U8 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[2]), .ZN(aes_state_regs_0_n199) );
  OAI21_X1 aes_state_regs_0_U7 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n30), .A(aes_state_regs_0_n199), .ZN(StateOutxD[2])
         );
  NAND2_X1 aes_state_regs_0_U6 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[1]), .ZN(aes_state_regs_0_n200) );
  OAI21_X1 aes_state_regs_0_U5 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n29), .A(aes_state_regs_0_n200), .ZN(StateOutxD[1])
         );
  OR2_X1 aes_state_regs_0_U4 ( .A1(aes_state_regs_0_n177), .A2(doMixColumnsxS), 
        .ZN(aes_state_regs_0_n195) );
  INV_X2 aes_state_regs_0_U3 ( .A(aes_state_regs_0_n109), .ZN(
        aes_state_regs_0_n202) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_7_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[7]), .SI(aes_state_regs_0_S10xDP_7_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[7]), .QN(aes_state_regs_0_n28) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_6_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[6]), .SI(aes_state_regs_0_S10xDP_6_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[6]), .QN(aes_state_regs_0_n34) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_5_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[5]), .SI(aes_state_regs_0_S10xDP_5_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[5]), .QN(aes_state_regs_0_n33) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_4_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[4]), .SI(aes_state_regs_0_S10xDP_4_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[4]), .QN(aes_state_regs_0_n32) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_3_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[3]), .SI(aes_state_regs_0_S10xDP_3_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[3]), .QN(aes_state_regs_0_n31) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_2_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[2]), .SI(aes_state_regs_0_S10xDP_2_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[2]), .QN(aes_state_regs_0_n30) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_1_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[1]), .SI(aes_state_regs_0_S10xDP_1_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[1]), .QN(aes_state_regs_0_n29) );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_7_ ( .D(aes_state_regs_0_S10xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_7_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_6_ ( .D(aes_state_regs_0_S10xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_6_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_5_ ( .D(aes_state_regs_0_S10xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_5_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_4_ ( .D(aes_state_regs_0_S10xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_4_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_3_ ( .D(aes_state_regs_0_S10xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_3_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_2_ ( .D(aes_state_regs_0_S10xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_2_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_1_ ( .D(aes_state_regs_0_S10xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_7_ ( .D(aes_state_regs_0_S01xDO_7_), 
        .SI(StateInxD[7]), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_7_), .QN(aes_state_regs_0_n36) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_7_ ( .D(aes_state_regs_0_n173), .SI(
        aes_state_regs_0_n170), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[7]), .QN(aes_state_regs_0_n127) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_7_ ( .D(aes_state_regs_0_S02xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_7_ ( .D(aes_state_regs_0_n172), .SI(
        aes_state_regs_0_S23xDP_7_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_7_ ( .D(aes_state_regs_0_n170), .SI(
        aes_state_regs_0_n173), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_7_ ( .D(aes_state_regs_0_S02xDP_7_), 
        .SI(aes_state_regs_0_S01xDO_7_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n173), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_7_ ( .D(aes_state_regs_0_S01xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_7_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_7_ ( .D(aes_state_regs_0_S21xDP[7]), 
        .SI(aes_state_regs_0_n172), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_7_ ( .D(aes_state_regs_0_n171), .SI(
        aes_state_regs_0_S30xDP_7_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n172), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_7_ ( .D(aes_state_regs_0_n169), .SI(
        aes_state_regs_0_S02xDP_7_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n171), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_7_ ( .D(StateInxD[7]), .SI(
        aes_state_regs_0_n169), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n170), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_7_ ( .D(aes_state_regs_0_S03xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n169), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_7_ ( .D(aes_state_regs_0_S23xDP_7_), 
        .SI(aes_state_regs_0_S20xDP_7_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[7]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_7_ ( .D(aes_state_regs_0_S20xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_7_), .QN(
        aes_state_regs_0_n44) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_6_ ( .D(aes_state_regs_0_S01xDO_6_), 
        .SI(StateInxD[6]), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_6_), .QN(aes_state_regs_0_n37) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_6_ ( .D(aes_state_regs_0_n168), .SI(
        aes_state_regs_0_n165), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[6]), .QN(aes_state_regs_0_n126) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_6_ ( .D(aes_state_regs_0_S02xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_6_ ( .D(aes_state_regs_0_n167), .SI(
        aes_state_regs_0_S23xDP_6_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_6_ ( .D(aes_state_regs_0_n165), .SI(
        aes_state_regs_0_n168), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_6_ ( .D(aes_state_regs_0_S02xDP_6_), 
        .SI(aes_state_regs_0_S01xDO_6_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n168), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_6_ ( .D(aes_state_regs_0_S01xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_6_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_6_ ( .D(aes_state_regs_0_S21xDP[6]), 
        .SI(aes_state_regs_0_n167), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_6_ ( .D(aes_state_regs_0_n166), .SI(
        aes_state_regs_0_S30xDP_6_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n167), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_6_ ( .D(aes_state_regs_0_n164), .SI(
        aes_state_regs_0_S02xDP_6_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n166), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_6_ ( .D(StateInxD[6]), .SI(
        aes_state_regs_0_n164), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n165), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_6_ ( .D(aes_state_regs_0_S03xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n164), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_6_ ( .D(aes_state_regs_0_S23xDP_6_), 
        .SI(aes_state_regs_0_S20xDP_6_), .SE(aes_state_regs_0_n177), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[6]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_6_ ( .D(aes_state_regs_0_S20xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_6_), .QN(
        aes_state_regs_0_n45) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_5_ ( .D(aes_state_regs_0_S01xDO_5_), 
        .SI(StateInxD[5]), .SE(nextRCONxS), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S30xDP_5_), .QN(aes_state_regs_0_n38) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_5_ ( .D(aes_state_regs_0_n163), .SI(
        aes_state_regs_0_n160), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[5]), .QN(aes_state_regs_0_n125) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_5_ ( .D(aes_state_regs_0_S02xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_5_ ( .D(aes_state_regs_0_n162), .SI(
        aes_state_regs_0_S23xDP_5_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_5_ ( .D(aes_state_regs_0_n160), .SI(
        aes_state_regs_0_n163), .SE(nextRCONxS), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S23xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_5_ ( .D(aes_state_regs_0_S02xDP_5_), 
        .SI(aes_state_regs_0_S01xDO_5_), .SE(aes_state_regs_0_n177), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n163), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_5_ ( .D(aes_state_regs_0_S01xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_5_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_5_ ( .D(aes_state_regs_0_S21xDP[5]), 
        .SI(aes_state_regs_0_n162), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_5_ ( .D(aes_state_regs_0_n161), .SI(
        aes_state_regs_0_S30xDP_5_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n162), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_5_ ( .D(aes_state_regs_0_n159), .SI(
        aes_state_regs_0_S02xDP_5_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n161), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_5_ ( .D(StateInxD[5]), .SI(
        aes_state_regs_0_n159), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n160), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_5_ ( .D(aes_state_regs_0_S03xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n159), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_5_ ( .D(aes_state_regs_0_S23xDP_5_), 
        .SI(aes_state_regs_0_S20xDP_5_), .SE(aes_state_regs_0_n177), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[5]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_5_ ( .D(aes_state_regs_0_S20xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_5_), .QN(
        aes_state_regs_0_n46) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_4_ ( .D(aes_state_regs_0_S01xDO_4_), 
        .SI(StateInxD[4]), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_4_), .QN(aes_state_regs_0_n39) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_4_ ( .D(aes_state_regs_0_n158), .SI(
        aes_state_regs_0_n155), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[4]), .QN(aes_state_regs_0_n124) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_4_ ( .D(aes_state_regs_0_S02xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_4_ ( .D(aes_state_regs_0_n157), .SI(
        aes_state_regs_0_S23xDP_4_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_4_ ( .D(aes_state_regs_0_n155), .SI(
        aes_state_regs_0_n158), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_4_ ( .D(aes_state_regs_0_S02xDP_4_), 
        .SI(aes_state_regs_0_S01xDO_4_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n158), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_4_ ( .D(aes_state_regs_0_S01xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_4_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_4_ ( .D(aes_state_regs_0_S21xDP[4]), 
        .SI(aes_state_regs_0_n157), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_4_ ( .D(aes_state_regs_0_n156), .SI(
        aes_state_regs_0_S30xDP_4_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n157), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_4_ ( .D(aes_state_regs_0_n154), .SI(
        aes_state_regs_0_S02xDP_4_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n156), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_4_ ( .D(StateInxD[4]), .SI(
        aes_state_regs_0_n154), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n155), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_4_ ( .D(aes_state_regs_0_S03xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n154), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_4_ ( .D(aes_state_regs_0_S23xDP_4_), 
        .SI(aes_state_regs_0_S20xDP_4_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[4]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_4_ ( .D(aes_state_regs_0_S20xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_4_), .QN(
        aes_state_regs_0_n47) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_3_ ( .D(aes_state_regs_0_S01xDO_3_), 
        .SI(StateInxD[3]), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_3_), .QN(aes_state_regs_0_n40) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_3_ ( .D(aes_state_regs_0_n153), .SI(
        aes_state_regs_0_n150), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[3]), .QN(aes_state_regs_0_n123) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_3_ ( .D(aes_state_regs_0_S02xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_3_ ( .D(aes_state_regs_0_n152), .SI(
        aes_state_regs_0_S23xDP_3_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_3_ ( .D(aes_state_regs_0_n150), .SI(
        aes_state_regs_0_n153), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_3_ ( .D(aes_state_regs_0_S02xDP_3_), 
        .SI(aes_state_regs_0_S01xDO_3_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n153), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_3_ ( .D(aes_state_regs_0_S01xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_3_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_3_ ( .D(aes_state_regs_0_S21xDP[3]), 
        .SI(aes_state_regs_0_n152), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_3_ ( .D(aes_state_regs_0_n151), .SI(
        aes_state_regs_0_S30xDP_3_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n152), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_3_ ( .D(aes_state_regs_0_n149), .SI(
        aes_state_regs_0_S02xDP_3_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n151), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_3_ ( .D(StateInxD[3]), .SI(
        aes_state_regs_0_n149), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n150), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_3_ ( .D(aes_state_regs_0_S03xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n149), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_3_ ( .D(aes_state_regs_0_S23xDP_3_), 
        .SI(aes_state_regs_0_S20xDP_3_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[3]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_3_ ( .D(aes_state_regs_0_S20xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_3_), .QN(
        aes_state_regs_0_n48) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_2_ ( .D(aes_state_regs_0_S01xDO_2_), 
        .SI(StateInxD[2]), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_2_), .QN(aes_state_regs_0_n41) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_2_ ( .D(aes_state_regs_0_n148), .SI(
        aes_state_regs_0_n145), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[2]), .QN(aes_state_regs_0_n122) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_2_ ( .D(aes_state_regs_0_S02xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_2_ ( .D(aes_state_regs_0_n147), .SI(
        aes_state_regs_0_S23xDP_2_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_2_ ( .D(aes_state_regs_0_n145), .SI(
        aes_state_regs_0_n148), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_2_ ( .D(aes_state_regs_0_S02xDP_2_), 
        .SI(aes_state_regs_0_S01xDO_2_), .SE(aes_state_regs_0_n177), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n148), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_2_ ( .D(aes_state_regs_0_S01xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_2_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_2_ ( .D(aes_state_regs_0_S21xDP[2]), 
        .SI(aes_state_regs_0_n147), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_2_ ( .D(aes_state_regs_0_n146), .SI(
        aes_state_regs_0_S30xDP_2_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n147), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_2_ ( .D(aes_state_regs_0_n144), .SI(
        aes_state_regs_0_S02xDP_2_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n146), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_2_ ( .D(StateInxD[2]), .SI(
        aes_state_regs_0_n144), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n145), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_2_ ( .D(aes_state_regs_0_S03xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n144), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_2_ ( .D(aes_state_regs_0_S23xDP_2_), 
        .SI(aes_state_regs_0_S20xDP_2_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[2]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_2_ ( .D(aes_state_regs_0_S20xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_2_), .QN(
        aes_state_regs_0_n49) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_1_ ( .D(aes_state_regs_0_S01xDO_1_), 
        .SI(StateInxD[1]), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_1_), .QN(aes_state_regs_0_n42) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_1_ ( .D(aes_state_regs_0_n143), .SI(
        aes_state_regs_0_n140), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[1]), .QN(aes_state_regs_0_n121) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_1_ ( .D(aes_state_regs_0_S02xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_1_ ( .D(aes_state_regs_0_n142), .SI(
        aes_state_regs_0_S23xDP_1_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_1_ ( .D(aes_state_regs_0_n140), .SI(
        aes_state_regs_0_n143), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_1_ ( .D(aes_state_regs_0_S02xDP_1_), 
        .SI(aes_state_regs_0_S01xDO_1_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n143), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_1_ ( .D(aes_state_regs_0_S01xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_1_ ( .D(aes_state_regs_0_S21xDP[1]), 
        .SI(aes_state_regs_0_n142), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_1_ ( .D(aes_state_regs_0_n141), .SI(
        aes_state_regs_0_S30xDP_1_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n142), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_1_ ( .D(aes_state_regs_0_n139), .SI(
        aes_state_regs_0_S02xDP_1_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n141), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_1_ ( .D(StateInxD[1]), .SI(
        aes_state_regs_0_n139), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n140), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_1_ ( .D(aes_state_regs_0_S03xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n139), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_1_ ( .D(aes_state_regs_0_S23xDP_1_), 
        .SI(aes_state_regs_0_S20xDP_1_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[1]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_1_ ( .D(aes_state_regs_0_S20xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_1_), .QN(
        aes_state_regs_0_n50) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_0_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[0]), .SI(aes_state_regs_0_S10xDP_0_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[0]), .QN(aes_state_regs_0_n35) );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_0_ ( .D(aes_state_regs_0_S10xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_0_ ( .D(aes_state_regs_0_n137), .SI(
        aes_state_regs_0_S31xDP_0_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S23xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_0_ ( .D(aes_state_regs_0_S02xDP_0_), 
        .SI(aes_state_regs_0_S01xDO_0_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S31xDP_0_), .QN() );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_0_ ( .D(aes_state_regs_0_S02xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_0_ ( .D(aes_state_regs_0_S22xDP_0_), 
        .SI(aes_state_regs_0_S23xDP_0_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_0_ ( .D(aes_state_regs_0_n136), .SI(
        aes_state_regs_0_S30xDP_0_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S22xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_0_ ( .D(aes_state_regs_0_S01xDO_0_), 
        .SI(StateInxD[0]), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_0_), .QN(aes_state_regs_0_n43) );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_0_ ( .D(aes_state_regs_0_S01xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_0_ ( .D(aes_state_regs_0_n138), .SI(
        aes_state_regs_0_S22xDP_0_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_0_ ( .D(aes_state_regs_0_S31xDP_0_), 
        .SI(aes_state_regs_0_n137), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n138), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_0_ ( .D(StateInxD[0]), .SI(
        aes_state_regs_0_S03xDP_0_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n137), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_0_ ( .D(aes_state_regs_0_S03xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_0_ ( .D(aes_state_regs_0_S23xDP_0_), 
        .SI(aes_state_regs_0_S20xDP_0_), .SE(aes_state_regs_0_n177), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[0]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_0_ ( .D(aes_state_regs_0_S20xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_0_), .QN(
        aes_state_regs_0_n51) );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_0_ ( .D(aes_state_regs_0_S03xDP_0_), 
        .SI(aes_state_regs_0_S02xDP_0_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n136), .QN() );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U119 ( .A(
        aes_state_regs_0_mix_columns_1_n245), .B(
        aes_state_regs_0_mix_columns_1_n244), .ZN(
        aes_state_regs_0_MixColumnsS3xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U118 ( .A(
        aes_state_regs_0_mix_columns_1_n240), .B(
        aes_state_regs_0_mix_columns_1_n239), .ZN(
        aes_state_regs_0_MixColumnsS3xD[6]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U117 ( .A(
        aes_state_regs_0_mix_columns_1_n235), .B(
        aes_state_regs_0_mix_columns_1_n234), .ZN(
        aes_state_regs_0_MixColumnsS3xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U116 ( .A(
        aes_state_regs_0_mix_columns_1_n226), .B(
        aes_state_regs_0_mix_columns_1_n225), .ZN(
        aes_state_regs_0_MixColumnsS3xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U115 ( .A(
        aes_state_regs_0_mix_columns_1_n182), .B(
        aes_state_regs_0_mix_columns_1_n241), .ZN(
        aes_state_regs_0_MixColumnsS1xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U114 ( .A(
        aes_state_regs_0_mix_columns_1_n190), .B(aes_state_regs_0_S00xDP[0]), 
        .ZN(aes_state_regs_0_mix_columns_1_n182) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U113 ( .A(
        aes_state_regs_0_mix_columns_1_n180), .B(
        aes_state_regs_0_mix_columns_1_n181), .ZN(
        aes_state_regs_0_MixColumnsS1xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U112 ( .A(aes_state_regs_0_S20xDP_1_), .B(aes_state_regs_0_S10xDP_1_), .ZN(aes_state_regs_0_mix_columns_1_n181) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U111 ( .A(
        aes_state_regs_0_mix_columns_1_n200), .B(aes_state_regs_0_S20xDP_2_), 
        .Z(aes_state_regs_0_mix_columns_1_n180) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U110 ( .A(
        aes_state_regs_0_mix_columns_1_n207), .B(
        aes_state_regs_0_mix_columns_1_n179), .ZN(
        aes_state_regs_0_mix_columns_1_n231) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U109 ( .A1(
        aes_state_regs_0_S30xDP_3_), .A2(aes_state_regs_0_mix_columns_1_n206), 
        .B1(aes_state_regs_0_S30xDP_7_), .B2(
        aes_state_regs_0_mix_columns_1_n178), .ZN(
        aes_state_regs_0_mix_columns_1_n179) );
  INV_X1 aes_state_regs_0_mix_columns_1_U108 ( .A(aes_state_regs_0_S30xDP_3_), 
        .ZN(aes_state_regs_0_mix_columns_1_n178) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U107 ( .A(
        aes_state_regs_0_mix_columns_1_n177), .B(
        aes_state_regs_0_mix_columns_1_n196), .ZN(
        aes_state_regs_0_MixColumnsS1xD[1]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U106 ( .A(
        aes_state_regs_0_mix_columns_1_n191), .B(aes_state_regs_0_S00xDP[1]), 
        .ZN(aes_state_regs_0_mix_columns_1_n177) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U105 ( .A(
        aes_state_regs_0_mix_columns_1_n176), .B(
        aes_state_regs_0_mix_columns_1_n203), .ZN(
        aes_state_regs_0_MixColumnsS1xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U104 ( .A(aes_state_regs_0_S20xDP_3_), .B(aes_state_regs_0_mix_columns_1_n192), .ZN(
        aes_state_regs_0_mix_columns_1_n176) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U103 ( .A(
        aes_state_regs_0_mix_columns_1_n175), .B(
        aes_state_regs_0_mix_columns_1_n205), .ZN(
        aes_state_regs_0_MixColumnsS1xD[4]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U102 ( .A(
        aes_state_regs_0_mix_columns_1_n193), .B(aes_state_regs_0_S00xDP[4]), 
        .ZN(aes_state_regs_0_mix_columns_1_n175) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U101 ( .A1(
        aes_state_regs_0_S30xDP_2_), .A2(aes_state_regs_0_S30xDP_7_), .B1(
        aes_state_regs_0_mix_columns_1_n206), .B2(
        aes_state_regs_0_mix_columns_1_n174), .ZN(
        aes_state_regs_0_mix_columns_1_n228) );
  INV_X1 aes_state_regs_0_mix_columns_1_U100 ( .A(aes_state_regs_0_S30xDP_2_), 
        .ZN(aes_state_regs_0_mix_columns_1_n174) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U99 ( .A(
        aes_state_regs_0_mix_columns_1_n172), .B(
        aes_state_regs_0_mix_columns_1_n173), .ZN(
        aes_state_regs_0_MixColumnsS1xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U98 ( .A(aes_state_regs_0_S20xDP_4_), 
        .B(aes_state_regs_0_S10xDP_4_), .ZN(
        aes_state_regs_0_mix_columns_1_n173) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U97 ( .A(aes_state_regs_0_S00xDP[5]), 
        .B(aes_state_regs_0_mix_columns_1_n211), .Z(
        aes_state_regs_0_mix_columns_1_n172) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U96 ( .A(
        aes_state_regs_0_mix_columns_1_n171), .B(
        aes_state_regs_0_mix_columns_1_n170), .ZN(
        aes_state_regs_0_MixColumnsS1xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U95 ( .A(aes_state_regs_0_S10xDP_6_), 
        .B(aes_state_regs_0_mix_columns_1_n217), .ZN(
        aes_state_regs_0_mix_columns_1_n171) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U94 ( .A1(aes_state_regs_0_S20xDP_6_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n236), .ZN(
        aes_state_regs_0_mix_columns_1_n170) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U93 ( .A(
        aes_state_regs_0_mix_columns_1_n168), .B(
        aes_state_regs_0_mix_columns_1_n169), .ZN(
        aes_state_regs_0_MixColumnsS1xD[6]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U92 ( .A(aes_state_regs_0_S20xDP_5_), 
        .B(aes_state_regs_0_S10xDP_5_), .ZN(
        aes_state_regs_0_mix_columns_1_n169) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U91 ( .A(aes_state_regs_0_S00xDP[6]), 
        .B(aes_state_regs_0_mix_columns_1_n215), .Z(
        aes_state_regs_0_mix_columns_1_n168) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U90 ( .A1(aes_state_regs_0_S20xDP_3_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n167), .ZN(
        aes_state_regs_0_mix_columns_1_n205) );
  INV_X1 aes_state_regs_0_mix_columns_1_U89 ( .A(aes_state_regs_0_S20xDP_3_), 
        .ZN(aes_state_regs_0_mix_columns_1_n167) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U88 ( .A(
        aes_state_regs_0_mix_columns_1_n165), .B(
        aes_state_regs_0_mix_columns_1_n166), .ZN(
        aes_state_regs_0_mix_columns_1_n227) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U87 ( .A(aes_state_regs_0_S20xDP_3_), 
        .B(aes_state_regs_0_S00xDP[7]), .ZN(
        aes_state_regs_0_mix_columns_1_n166) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U86 ( .A(aes_state_regs_0_S00xDP[2]), 
        .B(aes_state_regs_0_S10xDP_3_), .Z(aes_state_regs_0_mix_columns_1_n165) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U85 ( .A(
        aes_state_regs_0_mix_columns_1_n164), .B(
        aes_state_regs_0_mix_columns_1_n163), .ZN(
        aes_state_regs_0_mix_columns_1_n203) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U84 ( .A(aes_state_regs_0_S20xDP_2_), 
        .B(aes_state_regs_0_S30xDP_3_), .ZN(
        aes_state_regs_0_mix_columns_1_n164) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U83 ( .A1(aes_state_regs_0_S00xDP[3]), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n162), .ZN(
        aes_state_regs_0_mix_columns_1_n163) );
  INV_X1 aes_state_regs_0_mix_columns_1_U82 ( .A(aes_state_regs_0_S00xDP[3]), 
        .ZN(aes_state_regs_0_mix_columns_1_n162) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U81 ( .A(
        aes_state_regs_0_mix_columns_1_n161), .B(
        aes_state_regs_0_mix_columns_1_n209), .ZN(
        aes_state_regs_0_mix_columns_1_n193) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U80 ( .A(aes_state_regs_0_S10xDP_7_), 
        .B(aes_state_regs_0_S10xDP_3_), .ZN(
        aes_state_regs_0_mix_columns_1_n161) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U79 ( .A(
        aes_state_regs_0_mix_columns_1_n160), .B(
        aes_state_regs_0_mix_columns_1_n215), .ZN(
        aes_state_regs_0_MixColumnsS0xD[6]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U78 ( .A(aes_state_regs_0_S10xDP_6_), 
        .B(aes_state_regs_0_mix_columns_1_n233), .ZN(
        aes_state_regs_0_mix_columns_1_n160) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U77 ( .A(
        aes_state_regs_0_mix_columns_1_n159), .B(
        aes_state_regs_0_mix_columns_1_n211), .ZN(
        aes_state_regs_0_MixColumnsS0xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U76 ( .A(aes_state_regs_0_S10xDP_5_), 
        .B(aes_state_regs_0_mix_columns_1_n207), .ZN(
        aes_state_regs_0_mix_columns_1_n159) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U75 ( .A1(aes_state_regs_0_S20xDP_0_), .A2(aes_state_regs_0_mix_columns_1_n218), .B1(
        aes_state_regs_0_mix_columns_1_n217), .B2(
        aes_state_regs_0_mix_columns_1_n216), .ZN(
        aes_state_regs_0_mix_columns_1_n219) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U74 ( .A(
        aes_state_regs_0_mix_columns_1_n220), .B(
        aes_state_regs_0_mix_columns_1_n219), .ZN(
        aes_state_regs_0_MixColumnsS3xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U73 ( .A(aes_state_regs_0_S20xDP_7_), 
        .B(aes_state_regs_0_mix_columns_1_n197), .ZN(
        aes_state_regs_0_mix_columns_1_n195) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U72 ( .A(
        aes_state_regs_0_mix_columns_1_n195), .B(
        aes_state_regs_0_mix_columns_1_n220), .ZN(
        aes_state_regs_0_MixColumnsS2xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U71 ( .A(
        aes_state_regs_0_mix_columns_1_n221), .B(aes_state_regs_0_S20xDP_1_), 
        .ZN(aes_state_regs_0_mix_columns_1_n223) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U70 ( .A(
        aes_state_regs_0_mix_columns_1_n223), .B(
        aes_state_regs_0_mix_columns_1_n222), .ZN(
        aes_state_regs_0_MixColumnsS3xD[1]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U69 ( .A(aes_state_regs_0_S30xDP_1_), 
        .B(aes_state_regs_0_mix_columns_1_n224), .ZN(
        aes_state_regs_0_mix_columns_1_n225) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U68 ( .A(aes_state_regs_0_S00xDP[2]), 
        .B(aes_state_regs_0_S00xDP[1]), .Z(aes_state_regs_0_mix_columns_1_n226) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U67 ( .A(
        aes_state_regs_0_mix_columns_1_n227), .B(aes_state_regs_0_S00xDP[3]), 
        .ZN(aes_state_regs_0_mix_columns_1_n229) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U66 ( .A(
        aes_state_regs_0_mix_columns_1_n229), .B(
        aes_state_regs_0_mix_columns_1_n228), .ZN(
        aes_state_regs_0_MixColumnsS3xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U65 ( .A(
        aes_state_regs_0_mix_columns_1_n230), .B(aes_state_regs_0_S20xDP_4_), 
        .ZN(aes_state_regs_0_mix_columns_1_n232) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U64 ( .A(
        aes_state_regs_0_mix_columns_1_n232), .B(
        aes_state_regs_0_mix_columns_1_n231), .ZN(
        aes_state_regs_0_MixColumnsS3xD[4]) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U63 ( .A(
        aes_state_regs_0_mix_columns_1_n233), .B(aes_state_regs_0_S20xDP_5_), 
        .Z(aes_state_regs_0_mix_columns_1_n235) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U62 ( .A(aes_state_regs_0_S30xDP_4_), 
        .B(aes_state_regs_0_S00xDP[4]), .ZN(
        aes_state_regs_0_mix_columns_1_n234) );
  INV_X1 aes_state_regs_0_mix_columns_1_U61 ( .A(
        aes_state_regs_0_mix_columns_1_n238), .ZN(
        aes_state_regs_0_mix_columns_1_n237) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U60 ( .A1(aes_state_regs_0_S20xDP_6_), .A2(aes_state_regs_0_mix_columns_1_n238), .B1(
        aes_state_regs_0_mix_columns_1_n237), .B2(
        aes_state_regs_0_mix_columns_1_n236), .ZN(
        aes_state_regs_0_mix_columns_1_n239) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U59 ( .A(aes_state_regs_0_S30xDP_5_), 
        .B(aes_state_regs_0_S00xDP[5]), .ZN(
        aes_state_regs_0_mix_columns_1_n240) );
  INV_X1 aes_state_regs_0_mix_columns_1_U58 ( .A(aes_state_regs_0_S00xDP[6]), 
        .ZN(aes_state_regs_0_mix_columns_1_n243) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U57 ( .A(aes_state_regs_0_S30xDP_6_), 
        .B(aes_state_regs_0_mix_columns_1_n241), .ZN(
        aes_state_regs_0_mix_columns_1_n245) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U56 ( .A1(aes_state_regs_0_S00xDP[7]), .A2(aes_state_regs_0_S00xDP[6]), .B1(aes_state_regs_0_mix_columns_1_n243), 
        .B2(aes_state_regs_0_mix_columns_1_n242), .ZN(
        aes_state_regs_0_mix_columns_1_n244) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U55 ( .A(aes_state_regs_0_S30xDP_1_), 
        .B(aes_state_regs_0_mix_columns_1_n196), .ZN(
        aes_state_regs_0_mix_columns_1_n199) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U54 ( .A(
        aes_state_regs_0_mix_columns_1_n199), .B(
        aes_state_regs_0_mix_columns_1_n222), .ZN(
        aes_state_regs_0_MixColumnsS2xD[1]) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U53 ( .A(aes_state_regs_0_S10xDP_2_), 
        .B(aes_state_regs_0_mix_columns_1_n200), .Z(
        aes_state_regs_0_mix_columns_1_n201) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U52 ( .A(
        aes_state_regs_0_mix_columns_1_n202), .B(
        aes_state_regs_0_mix_columns_1_n201), .ZN(
        aes_state_regs_0_MixColumnsS2xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U51 ( .A(aes_state_regs_0_S10xDP_3_), 
        .B(aes_state_regs_0_mix_columns_1_n203), .ZN(
        aes_state_regs_0_mix_columns_1_n204) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U50 ( .A(
        aes_state_regs_0_mix_columns_1_n204), .B(
        aes_state_regs_0_mix_columns_1_n228), .ZN(
        aes_state_regs_0_MixColumnsS2xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U49 ( .A(aes_state_regs_0_S30xDP_4_), 
        .B(aes_state_regs_0_mix_columns_1_n205), .ZN(
        aes_state_regs_0_mix_columns_1_n208) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U48 ( .A(
        aes_state_regs_0_mix_columns_1_n208), .B(
        aes_state_regs_0_mix_columns_1_n231), .ZN(
        aes_state_regs_0_MixColumnsS2xD[4]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U47 ( .A(
        aes_state_regs_0_mix_columns_1_n209), .B(aes_state_regs_0_S30xDP_5_), 
        .ZN(aes_state_regs_0_mix_columns_1_n210) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U46 ( .A(
        aes_state_regs_0_mix_columns_1_n210), .B(
        aes_state_regs_0_mix_columns_1_n233), .ZN(
        aes_state_regs_0_MixColumnsS2xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U45 ( .A(
        aes_state_regs_0_mix_columns_1_n211), .B(aes_state_regs_0_S30xDP_6_), 
        .ZN(aes_state_regs_0_mix_columns_1_n212) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U44 ( .A(
        aes_state_regs_0_mix_columns_1_n212), .B(
        aes_state_regs_0_mix_columns_1_n238), .ZN(
        aes_state_regs_0_MixColumnsS2xD[6]) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U43 ( .A1(aes_state_regs_0_S10xDP_7_), .A2(aes_state_regs_0_mix_columns_1_n218), .B1(
        aes_state_regs_0_mix_columns_1_n217), .B2(
        aes_state_regs_0_mix_columns_1_n213), .ZN(
        aes_state_regs_0_mix_columns_1_n214) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U42 ( .A(
        aes_state_regs_0_mix_columns_1_n215), .B(
        aes_state_regs_0_mix_columns_1_n214), .ZN(
        aes_state_regs_0_MixColumnsS2xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U41 ( .A(aes_state_regs_0_S00xDP[7]), 
        .B(aes_state_regs_0_mix_columns_1_n184), .ZN(
        aes_state_regs_0_mix_columns_1_n183) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U40 ( .A(
        aes_state_regs_0_mix_columns_1_n183), .B(
        aes_state_regs_0_mix_columns_1_n190), .ZN(
        aes_state_regs_0_MixColumnsS0xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U39 ( .A(
        aes_state_regs_0_mix_columns_1_n241), .B(
        aes_state_regs_0_mix_columns_1_n238), .ZN(
        aes_state_regs_0_mix_columns_1_n189) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U38 ( .A(
        aes_state_regs_0_mix_columns_1_n189), .B(aes_state_regs_0_S30xDP_7_), 
        .ZN(aes_state_regs_0_MixColumnsS0xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U37 ( .A(aes_state_regs_0_S10xDP_4_), 
        .B(aes_state_regs_0_mix_columns_1_n230), .ZN(
        aes_state_regs_0_mix_columns_1_n188) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U36 ( .A(
        aes_state_regs_0_mix_columns_1_n188), .B(
        aes_state_regs_0_mix_columns_1_n193), .ZN(
        aes_state_regs_0_MixColumnsS0xD[4]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U35 ( .A(aes_state_regs_0_S30xDP_3_), 
        .B(aes_state_regs_0_mix_columns_1_n227), .ZN(
        aes_state_regs_0_mix_columns_1_n187) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U34 ( .A(
        aes_state_regs_0_mix_columns_1_n187), .B(
        aes_state_regs_0_mix_columns_1_n192), .ZN(
        aes_state_regs_0_MixColumnsS0xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U33 ( .A(aes_state_regs_0_S30xDP_2_), 
        .B(aes_state_regs_0_mix_columns_1_n224), .ZN(
        aes_state_regs_0_mix_columns_1_n186) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U32 ( .A(
        aes_state_regs_0_mix_columns_1_n186), .B(
        aes_state_regs_0_mix_columns_1_n198), .ZN(
        aes_state_regs_0_MixColumnsS0xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U31 ( .A(aes_state_regs_0_S10xDP_1_), 
        .B(aes_state_regs_0_mix_columns_1_n221), .ZN(
        aes_state_regs_0_mix_columns_1_n185) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U30 ( .A(
        aes_state_regs_0_mix_columns_1_n185), .B(
        aes_state_regs_0_mix_columns_1_n191), .ZN(
        aes_state_regs_0_MixColumnsS0xD[1]) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U29 ( .A(aes_state_regs_0_S10xDP_0_), 
        .B(aes_state_regs_0_S00xDP[0]), .Z(aes_state_regs_0_mix_columns_1_n220) );
  INV_X1 aes_state_regs_0_mix_columns_1_U28 ( .A(
        aes_state_regs_0_mix_columns_1_n217), .ZN(
        aes_state_regs_0_mix_columns_1_n218) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U27 ( .A1(aes_state_regs_0_S00xDP[7]), .A2(aes_state_regs_0_S30xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n206), 
        .B2(aes_state_regs_0_mix_columns_1_n242), .ZN(
        aes_state_regs_0_mix_columns_1_n217) );
  INV_X1 aes_state_regs_0_mix_columns_1_U26 ( .A(aes_state_regs_0_S20xDP_0_), 
        .ZN(aes_state_regs_0_mix_columns_1_n216) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U25 ( .A(aes_state_regs_0_S30xDP_0_), 
        .B(aes_state_regs_0_mix_columns_1_n206), .ZN(
        aes_state_regs_0_mix_columns_1_n197) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U24 ( .A1(aes_state_regs_0_S10xDP_7_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n213), .ZN(
        aes_state_regs_0_mix_columns_1_n241) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U23 ( .A(aes_state_regs_0_S30xDP_0_), 
        .B(aes_state_regs_0_S20xDP_0_), .Z(aes_state_regs_0_mix_columns_1_n190) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U22 ( .A(
        aes_state_regs_0_mix_columns_1_n198), .B(
        aes_state_regs_0_mix_columns_1_n197), .Z(
        aes_state_regs_0_mix_columns_1_n222) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U21 ( .A(aes_state_regs_0_S00xDP[7]), 
        .B(aes_state_regs_0_S00xDP[0]), .Z(aes_state_regs_0_mix_columns_1_n221) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U20 ( .A(aes_state_regs_0_S10xDP_2_), 
        .B(aes_state_regs_0_S20xDP_2_), .Z(aes_state_regs_0_mix_columns_1_n224) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U19 ( .A(aes_state_regs_0_S00xDP[7]), 
        .B(aes_state_regs_0_S00xDP[3]), .Z(aes_state_regs_0_mix_columns_1_n230) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U18 ( .A(aes_state_regs_0_S10xDP_5_), 
        .B(aes_state_regs_0_S00xDP[5]), .Z(aes_state_regs_0_mix_columns_1_n233) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U17 ( .A(aes_state_regs_0_S10xDP_6_), 
        .B(aes_state_regs_0_S00xDP[6]), .Z(aes_state_regs_0_mix_columns_1_n238) );
  INV_X1 aes_state_regs_0_mix_columns_1_U16 ( .A(aes_state_regs_0_S20xDP_6_), 
        .ZN(aes_state_regs_0_mix_columns_1_n236) );
  INV_X1 aes_state_regs_0_mix_columns_1_U15 ( .A(aes_state_regs_0_S00xDP[7]), 
        .ZN(aes_state_regs_0_mix_columns_1_n242) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U14 ( .A1(aes_state_regs_0_S20xDP_0_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n216), .ZN(
        aes_state_regs_0_mix_columns_1_n196) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U13 ( .A(aes_state_regs_0_S30xDP_2_), 
        .B(aes_state_regs_0_S00xDP[2]), .Z(aes_state_regs_0_mix_columns_1_n200) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U12 ( .A(aes_state_regs_0_S30xDP_1_), 
        .B(aes_state_regs_0_S20xDP_1_), .ZN(
        aes_state_regs_0_mix_columns_1_n202) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U11 ( .A(aes_state_regs_0_S30xDP_4_), 
        .B(aes_state_regs_0_S20xDP_4_), .Z(aes_state_regs_0_mix_columns_1_n209) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U10 ( .A(aes_state_regs_0_S30xDP_5_), 
        .B(aes_state_regs_0_S20xDP_5_), .Z(aes_state_regs_0_mix_columns_1_n211) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U9 ( .A(aes_state_regs_0_S30xDP_6_), 
        .B(aes_state_regs_0_S20xDP_6_), .Z(aes_state_regs_0_mix_columns_1_n215) );
  INV_X1 aes_state_regs_0_mix_columns_1_U8 ( .A(aes_state_regs_0_S10xDP_7_), 
        .ZN(aes_state_regs_0_mix_columns_1_n213) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U7 ( .A(
        aes_state_regs_0_mix_columns_1_n184), .B(
        aes_state_regs_0_mix_columns_1_n202), .ZN(
        aes_state_regs_0_mix_columns_1_n191) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U6 ( .A(aes_state_regs_0_S10xDP_7_), 
        .B(aes_state_regs_0_S10xDP_2_), .Z(aes_state_regs_0_mix_columns_1_n192) );
  INV_X1 aes_state_regs_0_mix_columns_1_U5 ( .A(aes_state_regs_0_S20xDP_7_), 
        .ZN(aes_state_regs_0_mix_columns_1_n194) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U4 ( .A(aes_state_regs_0_S10xDP_7_), 
        .B(aes_state_regs_0_S10xDP_0_), .Z(aes_state_regs_0_mix_columns_1_n184) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U3 ( .A(aes_state_regs_0_S10xDP_1_), 
        .B(aes_state_regs_0_S00xDP[1]), .Z(aes_state_regs_0_mix_columns_1_n198) );
  INV_X1 aes_state_regs_0_mix_columns_1_U2 ( .A(aes_state_regs_0_S30xDP_7_), 
        .ZN(aes_state_regs_0_mix_columns_1_n206) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U1 ( .A(aes_state_regs_0_S10xDP_4_), 
        .B(aes_state_regs_0_S00xDP[4]), .Z(aes_state_regs_0_mix_columns_1_n207) );
endmodule

