
module circuit ( CLK, RESET, DONE, MESSAGE1, MESSAGE2, RESULT1, RESULT2 );
  input [199:0] MESSAGE1;
  input [199:0] MESSAGE2;
  output [199:0] RESULT1;
  output [199:0] RESULT2;
  input CLK, RESET;
  output DONE;
  wire   RoundFunction_T1_n400, RoundFunction_T1_n399, RoundFunction_T1_n398,
         RoundFunction_T1_n397, RoundFunction_T1_n396, RoundFunction_T1_n395,
         RoundFunction_T1_n394, RoundFunction_T1_n393, RoundFunction_T1_n392,
         RoundFunction_T1_n391, RoundFunction_T1_n390, RoundFunction_T1_n389,
         RoundFunction_T1_n388, RoundFunction_T1_n387, RoundFunction_T1_n386,
         RoundFunction_T1_n385, RoundFunction_T1_n384, RoundFunction_T1_n383,
         RoundFunction_T1_n382, RoundFunction_T1_n381, RoundFunction_T1_n380,
         RoundFunction_T1_n379, RoundFunction_T1_n378, RoundFunction_T1_n377,
         RoundFunction_T1_n376, RoundFunction_T1_n375, RoundFunction_T1_n374,
         RoundFunction_T1_n373, RoundFunction_T1_n372, RoundFunction_T1_n371,
         RoundFunction_T1_n370, RoundFunction_T1_n369, RoundFunction_T1_n368,
         RoundFunction_T1_n367, RoundFunction_T1_n366, RoundFunction_T1_n365,
         RoundFunction_T1_n364, RoundFunction_T1_n363, RoundFunction_T1_n362,
         RoundFunction_T1_n361, RoundFunction_T1_n360, RoundFunction_T1_n359,
         RoundFunction_T1_n358, RoundFunction_T1_n357, RoundFunction_T1_n356,
         RoundFunction_T1_n355, RoundFunction_T1_n354, RoundFunction_T1_n353,
         RoundFunction_T1_n352, RoundFunction_T1_n351, RoundFunction_T1_n350,
         RoundFunction_T1_n349, RoundFunction_T1_n348, RoundFunction_T1_n347,
         RoundFunction_T1_n346, RoundFunction_T1_n345, RoundFunction_T1_n344,
         RoundFunction_T1_n343, RoundFunction_T1_n342, RoundFunction_T1_n341,
         RoundFunction_T1_n340, RoundFunction_T1_n339, RoundFunction_T1_n338,
         RoundFunction_T1_n337, RoundFunction_T1_n336, RoundFunction_T1_n335,
         RoundFunction_T1_n334, RoundFunction_T1_n333, RoundFunction_T1_n332,
         RoundFunction_T1_n331, RoundFunction_T1_n330, RoundFunction_T1_n329,
         RoundFunction_T1_n328, RoundFunction_T1_n327, RoundFunction_T1_n326,
         RoundFunction_T1_n325, RoundFunction_T1_n324, RoundFunction_T1_n323,
         RoundFunction_T1_n322, RoundFunction_T1_n321, RoundFunction_T1_n320,
         RoundFunction_T1_n319, RoundFunction_T1_n318, RoundFunction_T1_n317,
         RoundFunction_T1_n316, RoundFunction_T1_n315, RoundFunction_T1_n314,
         RoundFunction_T1_n313, RoundFunction_T1_n312, RoundFunction_T1_n311,
         RoundFunction_T1_n310, RoundFunction_T1_n309, RoundFunction_T1_n308,
         RoundFunction_T1_n307, RoundFunction_T1_n306, RoundFunction_T1_n305,
         RoundFunction_T1_n304, RoundFunction_T1_n303, RoundFunction_T1_n302,
         RoundFunction_T1_n301, RoundFunction_T1_n300, RoundFunction_T1_n299,
         RoundFunction_T1_n298, RoundFunction_T1_n297, RoundFunction_T1_n296,
         RoundFunction_T1_n295, RoundFunction_T1_n294, RoundFunction_T1_n293,
         RoundFunction_T1_n292, RoundFunction_T1_n291, RoundFunction_T1_n290,
         RoundFunction_T1_n289, RoundFunction_T1_n288, RoundFunction_T1_n287,
         RoundFunction_T1_n286, RoundFunction_T1_n285, RoundFunction_T1_n284,
         RoundFunction_T1_n283, RoundFunction_T1_n282, RoundFunction_T1_n281,
         RoundFunction_T1_n280, RoundFunction_T1_n279, RoundFunction_T1_n278,
         RoundFunction_T1_n277, RoundFunction_T1_n276, RoundFunction_T1_n275,
         RoundFunction_T1_n274, RoundFunction_T1_n273, RoundFunction_T1_n272,
         RoundFunction_T1_n271, RoundFunction_T1_n270, RoundFunction_T1_n269,
         RoundFunction_T1_n268, RoundFunction_T1_n267, RoundFunction_T1_n266,
         RoundFunction_T1_n265, RoundFunction_T1_n264, RoundFunction_T1_n263,
         RoundFunction_T1_n262, RoundFunction_T1_n261, RoundFunction_T1_n260,
         RoundFunction_T1_n259, RoundFunction_T1_n258, RoundFunction_T1_n257,
         RoundFunction_T1_n256, RoundFunction_T1_n255, RoundFunction_T1_n254,
         RoundFunction_T1_n253, RoundFunction_T1_n252, RoundFunction_T1_n251,
         RoundFunction_T1_n250, RoundFunction_T1_n249, RoundFunction_T1_n248,
         RoundFunction_T1_n247, RoundFunction_T1_n246, RoundFunction_T1_n245,
         RoundFunction_T1_n244, RoundFunction_T1_n243, RoundFunction_T1_n242,
         RoundFunction_T1_n241, RoundFunction_T1_n240, RoundFunction_T1_n239,
         RoundFunction_T1_n238, RoundFunction_T1_n237, RoundFunction_T1_n236,
         RoundFunction_T1_n235, RoundFunction_T1_n234, RoundFunction_T1_n233,
         RoundFunction_T1_n232, RoundFunction_T1_n231, RoundFunction_T1_n230,
         RoundFunction_T1_n229, RoundFunction_T1_n228, RoundFunction_T1_n227,
         RoundFunction_T1_n226, RoundFunction_T1_n225, RoundFunction_T1_n224,
         RoundFunction_T1_n223, RoundFunction_T1_n222, RoundFunction_T1_n221,
         RoundFunction_T1_n220, RoundFunction_T1_n219, RoundFunction_T1_n218,
         RoundFunction_T1_n217, RoundFunction_T1_n216, RoundFunction_T1_n215,
         RoundFunction_T1_n214, RoundFunction_T1_n213, RoundFunction_T1_n212,
         RoundFunction_T1_n211, RoundFunction_T1_n210, RoundFunction_T1_n209,
         RoundFunction_T1_n208, RoundFunction_T1_n207, RoundFunction_T1_n206,
         RoundFunction_T1_n205, RoundFunction_T1_n204, RoundFunction_T1_n203,
         RoundFunction_T1_n202, RoundFunction_T1_n201, RoundFunction_T2_n400,
         RoundFunction_T2_n399, RoundFunction_T2_n398, RoundFunction_T2_n397,
         RoundFunction_T2_n396, RoundFunction_T2_n395, RoundFunction_T2_n394,
         RoundFunction_T2_n393, RoundFunction_T2_n392, RoundFunction_T2_n391,
         RoundFunction_T2_n390, RoundFunction_T2_n389, RoundFunction_T2_n388,
         RoundFunction_T2_n387, RoundFunction_T2_n386, RoundFunction_T2_n385,
         RoundFunction_T2_n384, RoundFunction_T2_n383, RoundFunction_T2_n382,
         RoundFunction_T2_n381, RoundFunction_T2_n380, RoundFunction_T2_n379,
         RoundFunction_T2_n378, RoundFunction_T2_n377, RoundFunction_T2_n376,
         RoundFunction_T2_n375, RoundFunction_T2_n374, RoundFunction_T2_n373,
         RoundFunction_T2_n372, RoundFunction_T2_n371, RoundFunction_T2_n370,
         RoundFunction_T2_n369, RoundFunction_T2_n368, RoundFunction_T2_n367,
         RoundFunction_T2_n366, RoundFunction_T2_n365, RoundFunction_T2_n364,
         RoundFunction_T2_n363, RoundFunction_T2_n362, RoundFunction_T2_n361,
         RoundFunction_T2_n360, RoundFunction_T2_n359, RoundFunction_T2_n358,
         RoundFunction_T2_n357, RoundFunction_T2_n356, RoundFunction_T2_n355,
         RoundFunction_T2_n354, RoundFunction_T2_n353, RoundFunction_T2_n352,
         RoundFunction_T2_n351, RoundFunction_T2_n350, RoundFunction_T2_n349,
         RoundFunction_T2_n348, RoundFunction_T2_n347, RoundFunction_T2_n346,
         RoundFunction_T2_n345, RoundFunction_T2_n344, RoundFunction_T2_n343,
         RoundFunction_T2_n342, RoundFunction_T2_n341, RoundFunction_T2_n340,
         RoundFunction_T2_n339, RoundFunction_T2_n338, RoundFunction_T2_n337,
         RoundFunction_T2_n336, RoundFunction_T2_n335, RoundFunction_T2_n334,
         RoundFunction_T2_n333, RoundFunction_T2_n332, RoundFunction_T2_n331,
         RoundFunction_T2_n330, RoundFunction_T2_n329, RoundFunction_T2_n328,
         RoundFunction_T2_n327, RoundFunction_T2_n326, RoundFunction_T2_n325,
         RoundFunction_T2_n324, RoundFunction_T2_n323, RoundFunction_T2_n322,
         RoundFunction_T2_n321, RoundFunction_T2_n320, RoundFunction_T2_n319,
         RoundFunction_T2_n318, RoundFunction_T2_n317, RoundFunction_T2_n316,
         RoundFunction_T2_n315, RoundFunction_T2_n314, RoundFunction_T2_n313,
         RoundFunction_T2_n312, RoundFunction_T2_n311, RoundFunction_T2_n310,
         RoundFunction_T2_n309, RoundFunction_T2_n308, RoundFunction_T2_n307,
         RoundFunction_T2_n306, RoundFunction_T2_n305, RoundFunction_T2_n304,
         RoundFunction_T2_n303, RoundFunction_T2_n302, RoundFunction_T2_n301,
         RoundFunction_T2_n300, RoundFunction_T2_n299, RoundFunction_T2_n298,
         RoundFunction_T2_n297, RoundFunction_T2_n296, RoundFunction_T2_n295,
         RoundFunction_T2_n294, RoundFunction_T2_n293, RoundFunction_T2_n292,
         RoundFunction_T2_n291, RoundFunction_T2_n290, RoundFunction_T2_n289,
         RoundFunction_T2_n288, RoundFunction_T2_n287, RoundFunction_T2_n286,
         RoundFunction_T2_n285, RoundFunction_T2_n284, RoundFunction_T2_n283,
         RoundFunction_T2_n282, RoundFunction_T2_n281, RoundFunction_T2_n280,
         RoundFunction_T2_n279, RoundFunction_T2_n278, RoundFunction_T2_n277,
         RoundFunction_T2_n276, RoundFunction_T2_n275, RoundFunction_T2_n274,
         RoundFunction_T2_n273, RoundFunction_T2_n272, RoundFunction_T2_n271,
         RoundFunction_T2_n270, RoundFunction_T2_n269, RoundFunction_T2_n268,
         RoundFunction_T2_n267, RoundFunction_T2_n266, RoundFunction_T2_n265,
         RoundFunction_T2_n264, RoundFunction_T2_n263, RoundFunction_T2_n262,
         RoundFunction_T2_n261, RoundFunction_T2_n260, RoundFunction_T2_n259,
         RoundFunction_T2_n258, RoundFunction_T2_n257, RoundFunction_T2_n256,
         RoundFunction_T2_n255, RoundFunction_T2_n254, RoundFunction_T2_n253,
         RoundFunction_T2_n252, RoundFunction_T2_n251, RoundFunction_T2_n250,
         RoundFunction_T2_n249, RoundFunction_T2_n248, RoundFunction_T2_n247,
         RoundFunction_T2_n246, RoundFunction_T2_n245, RoundFunction_T2_n244,
         RoundFunction_T2_n243, RoundFunction_T2_n242, RoundFunction_T2_n241,
         RoundFunction_T2_n240, RoundFunction_T2_n239, RoundFunction_T2_n238,
         RoundFunction_T2_n237, RoundFunction_T2_n236, RoundFunction_T2_n235,
         RoundFunction_T2_n234, RoundFunction_T2_n233, RoundFunction_T2_n232,
         RoundFunction_T2_n231, RoundFunction_T2_n230, RoundFunction_T2_n229,
         RoundFunction_T2_n228, RoundFunction_T2_n227, RoundFunction_T2_n226,
         RoundFunction_T2_n225, RoundFunction_T2_n224, RoundFunction_T2_n223,
         RoundFunction_T2_n222, RoundFunction_T2_n221, RoundFunction_T2_n220,
         RoundFunction_T2_n219, RoundFunction_T2_n218, RoundFunction_T2_n217,
         RoundFunction_T2_n216, RoundFunction_T2_n215, RoundFunction_T2_n214,
         RoundFunction_T2_n213, RoundFunction_T2_n212, RoundFunction_T2_n211,
         RoundFunction_T2_n210, RoundFunction_T2_n209, RoundFunction_T2_n208,
         RoundFunction_T2_n207, RoundFunction_T2_n206, RoundFunction_T2_n205,
         RoundFunction_T2_n204, RoundFunction_T2_n203, RoundFunction_T2_n202,
         RoundFunction_T2_n201, RoundFunction_C_Inst_Chi_NoFresh_0_n1,
         RoundFunction_C_Inst_Chi_NoFresh_0_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_0_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_0_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_0_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_0_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_0_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_0_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_0_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_0_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_0_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_1_n1,
         RoundFunction_C_Inst_Chi_NoFresh_1_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_1_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_1_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_1_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_1_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_1_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_1_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_1_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_1_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_1_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_2_n1,
         RoundFunction_C_Inst_Chi_NoFresh_2_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_2_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_2_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_2_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_2_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_2_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_2_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_2_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_2_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_2_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_3_n1,
         RoundFunction_C_Inst_Chi_NoFresh_3_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_3_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_3_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_3_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_3_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_3_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_3_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_3_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_3_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_3_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_4_n1,
         RoundFunction_C_Inst_Chi_NoFresh_4_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_4_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_4_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_4_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_4_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_4_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_4_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_4_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_4_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_4_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_5_n1,
         RoundFunction_C_Inst_Chi_NoFresh_5_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_5_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_5_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_5_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_5_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_5_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_5_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_5_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_5_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_5_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_6_n1,
         RoundFunction_C_Inst_Chi_NoFresh_6_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_6_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_6_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_6_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_6_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_6_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_6_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_6_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_6_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_6_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_7_n1,
         RoundFunction_C_Inst_Chi_NoFresh_7_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_7_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_7_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_7_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_7_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_7_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_7_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_7_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_7_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_7_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_8_n1,
         RoundFunction_C_Inst_Chi_NoFresh_8_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_8_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_8_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_8_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_8_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_8_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_8_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_8_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_8_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_8_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_9_n1,
         RoundFunction_C_Inst_Chi_NoFresh_9_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_9_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_9_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_9_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_9_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_9_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_9_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_9_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_9_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_9_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_10_n1,
         RoundFunction_C_Inst_Chi_NoFresh_10_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_10_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_10_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_10_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_10_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_10_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_10_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_10_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_10_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_10_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_11_n1,
         RoundFunction_C_Inst_Chi_NoFresh_11_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_11_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_11_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_11_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_11_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_11_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_11_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_11_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_11_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_11_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_12_n1,
         RoundFunction_C_Inst_Chi_NoFresh_12_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_12_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_12_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_12_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_12_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_12_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_12_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_12_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_12_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_12_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_13_n1,
         RoundFunction_C_Inst_Chi_NoFresh_13_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_13_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_13_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_13_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_13_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_13_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_13_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_13_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_13_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_13_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_14_n1,
         RoundFunction_C_Inst_Chi_NoFresh_14_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_14_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_14_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_14_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_14_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_14_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_14_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_14_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_14_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_14_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_15_n1,
         RoundFunction_C_Inst_Chi_NoFresh_15_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_15_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_15_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_15_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_15_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_15_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_15_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_15_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_15_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_15_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_16_n1,
         RoundFunction_C_Inst_Chi_NoFresh_16_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_16_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_16_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_16_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_16_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_16_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_16_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_16_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_16_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_16_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_17_n1,
         RoundFunction_C_Inst_Chi_NoFresh_17_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_17_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_17_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_17_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_17_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_17_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_17_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_17_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_17_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_17_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_18_n1,
         RoundFunction_C_Inst_Chi_NoFresh_18_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_18_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_18_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_18_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_18_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_18_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_18_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_18_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_18_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_18_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_19_n1,
         RoundFunction_C_Inst_Chi_NoFresh_19_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_19_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_19_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_19_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_19_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_19_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_19_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_19_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_19_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_19_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_20_n1,
         RoundFunction_C_Inst_Chi_NoFresh_20_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_20_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_20_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_20_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_20_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_20_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_20_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_20_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_20_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_20_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_21_n1,
         RoundFunction_C_Inst_Chi_NoFresh_21_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_21_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_21_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_21_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_21_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_21_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_21_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_21_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_21_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_21_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_22_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_22_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_22_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_22_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_22_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_22_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_22_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_22_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_22_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_22_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_23_n1,
         RoundFunction_C_Inst_Chi_NoFresh_23_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_23_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_23_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_23_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_23_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_23_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_23_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_23_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_23_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_23_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_24_n1,
         RoundFunction_C_Inst_Chi_NoFresh_24_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_24_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_24_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_24_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_24_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_24_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_24_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_24_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_24_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_24_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_25_n1,
         RoundFunction_C_Inst_Chi_NoFresh_25_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_25_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_25_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_25_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_25_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_25_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_25_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_25_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_25_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_25_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_26_n1,
         RoundFunction_C_Inst_Chi_NoFresh_26_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_26_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_26_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_26_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_26_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_26_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_26_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_26_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_26_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_26_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_27_n1,
         RoundFunction_C_Inst_Chi_NoFresh_27_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_27_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_27_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_27_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_27_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_27_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_27_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_27_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_27_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_27_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_28_n1,
         RoundFunction_C_Inst_Chi_NoFresh_28_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_28_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_28_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_28_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_28_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_28_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_28_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_28_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_28_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_28_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_29_n1,
         RoundFunction_C_Inst_Chi_NoFresh_29_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_29_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_29_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_29_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_29_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_29_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_29_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_29_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_29_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_29_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_30_n1,
         RoundFunction_C_Inst_Chi_NoFresh_30_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_30_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_30_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_30_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_30_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_30_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_30_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_30_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_30_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_30_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_31_n1,
         RoundFunction_C_Inst_Chi_NoFresh_31_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_31_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_31_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_31_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_31_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_31_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_31_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_31_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_31_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_31_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_32_n1,
         RoundFunction_C_Inst_Chi_NoFresh_32_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_32_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_32_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_32_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_32_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_32_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_32_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_32_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_32_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_32_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_33_n1,
         RoundFunction_C_Inst_Chi_NoFresh_33_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_33_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_33_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_33_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_33_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_33_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_33_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_33_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_33_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_33_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_34_n1,
         RoundFunction_C_Inst_Chi_NoFresh_34_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_34_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_34_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_34_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_34_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_34_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_34_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_34_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_34_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_34_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_35_n1,
         RoundFunction_C_Inst_Chi_NoFresh_35_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_35_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_35_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_35_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_35_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_35_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_35_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_35_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_35_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_35_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_36_n1,
         RoundFunction_C_Inst_Chi_NoFresh_36_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_36_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_36_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_36_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_36_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_36_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_36_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_36_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_36_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_36_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_37_n1,
         RoundFunction_C_Inst_Chi_NoFresh_37_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_37_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_37_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_37_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_37_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_37_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_37_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_37_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_37_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_37_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_38_n1,
         RoundFunction_C_Inst_Chi_NoFresh_38_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_38_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_38_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_38_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_38_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_38_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_38_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_38_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_38_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_38_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_39_n1,
         RoundFunction_C_Inst_Chi_NoFresh_39_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_39_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_39_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_39_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_39_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_39_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_39_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_39_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_39_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_39_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_2__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_2__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_5__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_6__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_7__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_7__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_13__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_13__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_16__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_17__CF_Inst_n2,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n4,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n4, FSM_n152,
         FSM_n151, FSM_n150, FSM_n149, FSM_n148, FSM_n147, FSM_n146, FSM_n145,
         FSM_n144, FSM_n143, FSM_n142, FSM_n141, FSM_n140, FSM_n139, FSM_n138,
         FSM_n137, FSM_n136, FSM_n135, FSM_n134, FSM_n133, FSM_n132, FSM_n131,
         FSM_n130, FSM_n129, FSM_n128, FSM_n127, FSM_n126, FSM_n125, FSM_n124,
         FSM_n123, FSM_n122, FSM_n121, FSM_n120, FSM_n119, FSM_n118, FSM_n117,
         FSM_n116, FSM_n115, FSM_n114, FSM_n113, FSM_n112, FSM_n111, FSM_n110,
         FSM_n109, FSM_n108, FSM_n107, FSM_n106, FSM_n105, FSM_n104, FSM_n103,
         FSM_n102, FSM_n101, FSM_n100, FSM_n99, FSM_n98, FSM_n97, FSM_n96,
         FSM_n95, FSM_n94, FSM_n93, FSM_n92, FSM_n91, FSM_n87, FSM_n86,
         FSM_n85, FSM_n19, FSM_n9, FSM_n6, FSM_n4, FSM_n2, FSM_n79, FSM_n78,
         FSM_n77, FSM_n76, FSM_n75, FSM_n74, FSM_n73, FSM_n72, FSM_n71,
         FSM_n70, FSM_n12, FSM_n8, FSM_n7, FSM_n3, FSM_CONST_internal_3,
         FSM_CONST_internal_7;
  wire   [7:0] CONST;
  wire   [199:0] RoundFunction_TMP3_2;
  wire   [7:0] RoundFunction_TMP4_1;
  wire   [199:0] RoundFunction_TMP3_1;
  wire   [199:0] RoundFunction_STATE2;
  wire   [199:0] RoundFunction_STATE1;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg;
  wire   [19:0] RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out;
  wire   [1:0] FSM_CONST_internal;

  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_0_ ( .D(RESULT1[192]), 
        .SI(MESSAGE1[192]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[0]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_1_ ( .D(RESULT1[193]), 
        .SI(MESSAGE1[193]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[1]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_2_ ( .D(RESULT1[194]), 
        .SI(MESSAGE1[194]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[2]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_3_ ( .D(RESULT1[195]), 
        .SI(MESSAGE1[195]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[3]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_4_ ( .D(RESULT1[196]), 
        .SI(MESSAGE1[196]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[4]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_5_ ( .D(RESULT1[197]), 
        .SI(MESSAGE1[197]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[5]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_6_ ( .D(RESULT1[198]), 
        .SI(MESSAGE1[198]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[6]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_7_ ( .D(RESULT1[199]), 
        .SI(MESSAGE1[199]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[7]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_8_ ( .D(RESULT1[184]), 
        .SI(MESSAGE1[184]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[8]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_9_ ( .D(RESULT1[185]), 
        .SI(MESSAGE1[185]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[9]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_10_ ( .D(RESULT1[186]), 
        .SI(MESSAGE1[186]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[10]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_11_ ( .D(RESULT1[187]), 
        .SI(MESSAGE1[187]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[11]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_12_ ( .D(RESULT1[188]), 
        .SI(MESSAGE1[188]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[12]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_13_ ( .D(RESULT1[189]), 
        .SI(MESSAGE1[189]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[13]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_14_ ( .D(RESULT1[190]), 
        .SI(MESSAGE1[190]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[14]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_15_ ( .D(RESULT1[191]), 
        .SI(MESSAGE1[191]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[15]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_16_ ( .D(RESULT1[176]), 
        .SI(MESSAGE1[176]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[16]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_17_ ( .D(RESULT1[177]), 
        .SI(MESSAGE1[177]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[17]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_18_ ( .D(RESULT1[178]), 
        .SI(MESSAGE1[178]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[18]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_19_ ( .D(RESULT1[179]), 
        .SI(MESSAGE1[179]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[19]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_20_ ( .D(RESULT1[180]), 
        .SI(MESSAGE1[180]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[20]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_21_ ( .D(RESULT1[181]), 
        .SI(MESSAGE1[181]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[21]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_22_ ( .D(RESULT1[182]), 
        .SI(MESSAGE1[182]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[22]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_23_ ( .D(RESULT1[183]), 
        .SI(MESSAGE1[183]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[23]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_24_ ( .D(RESULT1[168]), 
        .SI(MESSAGE1[168]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[24]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_25_ ( .D(RESULT1[169]), 
        .SI(MESSAGE1[169]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[25]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_26_ ( .D(RESULT1[170]), 
        .SI(MESSAGE1[170]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[26]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_27_ ( .D(RESULT1[171]), 
        .SI(MESSAGE1[171]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[27]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_28_ ( .D(RESULT1[172]), 
        .SI(MESSAGE1[172]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[28]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_29_ ( .D(RESULT1[173]), 
        .SI(MESSAGE1[173]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[29]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_30_ ( .D(RESULT1[174]), 
        .SI(MESSAGE1[174]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[30]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_31_ ( .D(RESULT1[175]), 
        .SI(MESSAGE1[175]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[31]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_32_ ( .D(RESULT1[160]), 
        .SI(MESSAGE1[160]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[32]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_33_ ( .D(RESULT1[161]), 
        .SI(MESSAGE1[161]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[33]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_34_ ( .D(RESULT1[162]), 
        .SI(MESSAGE1[162]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[34]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_35_ ( .D(RESULT1[163]), 
        .SI(MESSAGE1[163]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[35]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_36_ ( .D(RESULT1[164]), 
        .SI(MESSAGE1[164]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[36]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_37_ ( .D(RESULT1[165]), 
        .SI(MESSAGE1[165]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[37]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_38_ ( .D(RESULT1[166]), 
        .SI(MESSAGE1[166]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[38]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_39_ ( .D(RESULT1[167]), 
        .SI(MESSAGE1[167]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[39]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_40_ ( .D(RESULT1[152]), 
        .SI(MESSAGE1[152]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[40]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_41_ ( .D(RESULT1[153]), 
        .SI(MESSAGE1[153]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[41]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_42_ ( .D(RESULT1[154]), 
        .SI(MESSAGE1[154]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[42]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_43_ ( .D(RESULT1[155]), 
        .SI(MESSAGE1[155]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[43]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_44_ ( .D(RESULT1[156]), 
        .SI(MESSAGE1[156]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[44]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_45_ ( .D(RESULT1[157]), 
        .SI(MESSAGE1[157]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[45]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_46_ ( .D(RESULT1[158]), 
        .SI(MESSAGE1[158]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[46]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_47_ ( .D(RESULT1[159]), 
        .SI(MESSAGE1[159]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[47]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_48_ ( .D(RESULT1[144]), 
        .SI(MESSAGE1[144]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[48]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_49_ ( .D(RESULT1[145]), 
        .SI(MESSAGE1[145]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[49]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_50_ ( .D(RESULT1[146]), 
        .SI(MESSAGE1[146]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[50]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_51_ ( .D(RESULT1[147]), 
        .SI(MESSAGE1[147]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[51]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_52_ ( .D(RESULT1[148]), 
        .SI(MESSAGE1[148]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[52]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_53_ ( .D(RESULT1[149]), 
        .SI(MESSAGE1[149]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[53]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_54_ ( .D(RESULT1[150]), 
        .SI(MESSAGE1[150]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[54]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_55_ ( .D(RESULT1[151]), 
        .SI(MESSAGE1[151]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[55]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_56_ ( .D(RESULT1[136]), 
        .SI(MESSAGE1[136]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[56]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_57_ ( .D(RESULT1[137]), 
        .SI(MESSAGE1[137]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[57]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_58_ ( .D(RESULT1[138]), 
        .SI(MESSAGE1[138]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[58]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_59_ ( .D(RESULT1[139]), 
        .SI(MESSAGE1[139]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[59]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_60_ ( .D(RESULT1[140]), 
        .SI(MESSAGE1[140]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[60]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_61_ ( .D(RESULT1[141]), 
        .SI(MESSAGE1[141]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[61]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_62_ ( .D(RESULT1[142]), 
        .SI(MESSAGE1[142]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[62]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_63_ ( .D(RESULT1[143]), 
        .SI(MESSAGE1[143]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[63]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_64_ ( .D(RESULT1[128]), 
        .SI(MESSAGE1[128]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[64]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_65_ ( .D(RESULT1[129]), 
        .SI(MESSAGE1[129]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[65]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_66_ ( .D(RESULT1[130]), 
        .SI(MESSAGE1[130]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[66]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_67_ ( .D(RESULT1[131]), 
        .SI(MESSAGE1[131]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[67]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_68_ ( .D(RESULT1[132]), 
        .SI(MESSAGE1[132]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[68]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_69_ ( .D(RESULT1[133]), 
        .SI(MESSAGE1[133]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[69]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_70_ ( .D(RESULT1[134]), 
        .SI(MESSAGE1[134]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[70]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_71_ ( .D(RESULT1[135]), 
        .SI(MESSAGE1[135]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[71]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_72_ ( .D(RESULT1[120]), 
        .SI(MESSAGE1[120]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[72]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_73_ ( .D(RESULT1[121]), 
        .SI(MESSAGE1[121]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[73]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_74_ ( .D(RESULT1[122]), 
        .SI(MESSAGE1[122]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[74]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_75_ ( .D(RESULT1[123]), 
        .SI(MESSAGE1[123]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[75]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_76_ ( .D(RESULT1[124]), 
        .SI(MESSAGE1[124]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[76]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_77_ ( .D(RESULT1[125]), 
        .SI(MESSAGE1[125]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[77]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_78_ ( .D(RESULT1[126]), 
        .SI(MESSAGE1[126]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[78]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_79_ ( .D(RESULT1[127]), 
        .SI(MESSAGE1[127]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[79]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_80_ ( .D(RESULT1[112]), 
        .SI(MESSAGE1[112]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[80]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_81_ ( .D(RESULT1[113]), 
        .SI(MESSAGE1[113]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[81]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_82_ ( .D(RESULT1[114]), 
        .SI(MESSAGE1[114]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[82]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_83_ ( .D(RESULT1[115]), 
        .SI(MESSAGE1[115]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[83]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_84_ ( .D(RESULT1[116]), 
        .SI(MESSAGE1[116]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[84]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_85_ ( .D(RESULT1[117]), 
        .SI(MESSAGE1[117]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[85]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_86_ ( .D(RESULT1[118]), 
        .SI(MESSAGE1[118]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[86]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_87_ ( .D(RESULT1[119]), 
        .SI(MESSAGE1[119]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[87]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_88_ ( .D(RESULT1[104]), 
        .SI(MESSAGE1[104]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[88]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_89_ ( .D(RESULT1[105]), 
        .SI(MESSAGE1[105]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[89]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_90_ ( .D(RESULT1[106]), 
        .SI(MESSAGE1[106]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[90]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_91_ ( .D(RESULT1[107]), 
        .SI(MESSAGE1[107]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[91]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_92_ ( .D(RESULT1[108]), 
        .SI(MESSAGE1[108]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[92]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_93_ ( .D(RESULT1[109]), 
        .SI(MESSAGE1[109]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[93]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_94_ ( .D(RESULT1[110]), 
        .SI(MESSAGE1[110]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[94]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_95_ ( .D(RESULT1[111]), 
        .SI(MESSAGE1[111]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[95]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_96_ ( .D(RESULT1[96]), 
        .SI(MESSAGE1[96]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[96]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_97_ ( .D(RESULT1[97]), 
        .SI(MESSAGE1[97]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[97]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_98_ ( .D(RESULT1[98]), 
        .SI(MESSAGE1[98]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[98]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_99_ ( .D(RESULT1[99]), 
        .SI(MESSAGE1[99]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[99]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_100_ ( .D(RESULT1[100]), 
        .SI(MESSAGE1[100]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[100]), .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_101_ ( .D(RESULT1[101]), 
        .SI(MESSAGE1[101]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[101]), .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_102_ ( .D(RESULT1[102]), 
        .SI(MESSAGE1[102]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[102]), .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_103_ ( .D(RESULT1[103]), 
        .SI(MESSAGE1[103]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[103]), .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_104_ ( .D(RESULT1[88]), 
        .SI(MESSAGE1[88]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[104]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_105_ ( .D(RESULT1[89]), 
        .SI(MESSAGE1[89]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[105]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_106_ ( .D(RESULT1[90]), 
        .SI(MESSAGE1[90]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[106]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_107_ ( .D(RESULT1[91]), 
        .SI(MESSAGE1[91]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[107]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_108_ ( .D(RESULT1[92]), 
        .SI(MESSAGE1[92]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[108]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_109_ ( .D(RESULT1[93]), 
        .SI(MESSAGE1[93]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[109]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_110_ ( .D(RESULT1[94]), 
        .SI(MESSAGE1[94]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[110]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_111_ ( .D(RESULT1[95]), 
        .SI(MESSAGE1[95]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[111]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_112_ ( .D(RESULT1[80]), 
        .SI(MESSAGE1[80]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[112]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_113_ ( .D(RESULT1[81]), 
        .SI(MESSAGE1[81]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[113]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_114_ ( .D(RESULT1[82]), 
        .SI(MESSAGE1[82]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[114]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_115_ ( .D(RESULT1[83]), 
        .SI(MESSAGE1[83]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[115]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_116_ ( .D(RESULT1[84]), 
        .SI(MESSAGE1[84]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[116]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_117_ ( .D(RESULT1[85]), 
        .SI(MESSAGE1[85]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[117]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_118_ ( .D(RESULT1[86]), 
        .SI(MESSAGE1[86]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[118]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_119_ ( .D(RESULT1[87]), 
        .SI(MESSAGE1[87]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[119]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_120_ ( .D(RESULT1[72]), 
        .SI(MESSAGE1[72]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[120]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_121_ ( .D(RESULT1[73]), 
        .SI(MESSAGE1[73]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[121]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_122_ ( .D(RESULT1[74]), 
        .SI(MESSAGE1[74]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[122]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_123_ ( .D(RESULT1[75]), 
        .SI(MESSAGE1[75]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[123]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_124_ ( .D(RESULT1[76]), 
        .SI(MESSAGE1[76]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[124]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_125_ ( .D(RESULT1[77]), 
        .SI(MESSAGE1[77]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[125]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_126_ ( .D(RESULT1[78]), 
        .SI(MESSAGE1[78]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[126]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_127_ ( .D(RESULT1[79]), 
        .SI(MESSAGE1[79]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[127]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_128_ ( .D(RESULT1[64]), 
        .SI(MESSAGE1[64]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[128]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_129_ ( .D(RESULT1[65]), 
        .SI(MESSAGE1[65]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[129]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_130_ ( .D(RESULT1[66]), 
        .SI(MESSAGE1[66]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[130]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_131_ ( .D(RESULT1[67]), 
        .SI(MESSAGE1[67]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[131]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_132_ ( .D(RESULT1[68]), 
        .SI(MESSAGE1[68]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[132]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_133_ ( .D(RESULT1[69]), 
        .SI(MESSAGE1[69]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[133]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_134_ ( .D(RESULT1[70]), 
        .SI(MESSAGE1[70]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[134]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_135_ ( .D(RESULT1[71]), 
        .SI(MESSAGE1[71]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[135]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_136_ ( .D(RESULT1[56]), 
        .SI(MESSAGE1[56]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[136]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_137_ ( .D(RESULT1[57]), 
        .SI(MESSAGE1[57]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[137]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_138_ ( .D(RESULT1[58]), 
        .SI(MESSAGE1[58]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[138]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_139_ ( .D(RESULT1[59]), 
        .SI(MESSAGE1[59]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[139]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_140_ ( .D(RESULT1[60]), 
        .SI(MESSAGE1[60]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[140]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_141_ ( .D(RESULT1[61]), 
        .SI(MESSAGE1[61]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[141]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_142_ ( .D(RESULT1[62]), 
        .SI(MESSAGE1[62]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[142]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_143_ ( .D(RESULT1[63]), 
        .SI(MESSAGE1[63]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[143]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_144_ ( .D(RESULT1[48]), 
        .SI(MESSAGE1[48]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[144]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_145_ ( .D(RESULT1[49]), 
        .SI(MESSAGE1[49]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[145]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_146_ ( .D(RESULT1[50]), 
        .SI(MESSAGE1[50]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[146]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_147_ ( .D(RESULT1[51]), 
        .SI(MESSAGE1[51]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[147]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_148_ ( .D(RESULT1[52]), 
        .SI(MESSAGE1[52]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[148]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_149_ ( .D(RESULT1[53]), 
        .SI(MESSAGE1[53]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[149]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_150_ ( .D(RESULT1[54]), 
        .SI(MESSAGE1[54]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[150]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_151_ ( .D(RESULT1[55]), 
        .SI(MESSAGE1[55]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[151]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_152_ ( .D(RESULT1[40]), 
        .SI(MESSAGE1[40]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[152]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_153_ ( .D(RESULT1[41]), 
        .SI(MESSAGE1[41]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[153]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_154_ ( .D(RESULT1[42]), 
        .SI(MESSAGE1[42]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[154]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_155_ ( .D(RESULT1[43]), 
        .SI(MESSAGE1[43]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[155]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_156_ ( .D(RESULT1[44]), 
        .SI(MESSAGE1[44]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[156]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_157_ ( .D(RESULT1[45]), 
        .SI(MESSAGE1[45]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[157]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_158_ ( .D(RESULT1[46]), 
        .SI(MESSAGE1[46]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[158]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_159_ ( .D(RESULT1[47]), 
        .SI(MESSAGE1[47]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[159]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_160_ ( .D(RESULT1[32]), 
        .SI(MESSAGE1[32]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[160]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_161_ ( .D(RESULT1[33]), 
        .SI(MESSAGE1[33]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[161]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_162_ ( .D(RESULT1[34]), 
        .SI(MESSAGE1[34]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[162]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_163_ ( .D(RESULT1[35]), 
        .SI(MESSAGE1[35]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[163]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_164_ ( .D(RESULT1[36]), 
        .SI(MESSAGE1[36]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[164]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_165_ ( .D(RESULT1[37]), 
        .SI(MESSAGE1[37]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[165]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_166_ ( .D(RESULT1[38]), 
        .SI(MESSAGE1[38]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[166]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_167_ ( .D(RESULT1[39]), 
        .SI(MESSAGE1[39]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[167]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_168_ ( .D(RESULT1[24]), 
        .SI(MESSAGE1[24]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[168]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_169_ ( .D(RESULT1[25]), 
        .SI(MESSAGE1[25]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[169]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_170_ ( .D(RESULT1[26]), 
        .SI(MESSAGE1[26]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[170]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_171_ ( .D(RESULT1[27]), 
        .SI(MESSAGE1[27]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[171]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_172_ ( .D(RESULT1[28]), 
        .SI(MESSAGE1[28]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[172]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_173_ ( .D(RESULT1[29]), 
        .SI(MESSAGE1[29]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[173]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_174_ ( .D(RESULT1[30]), 
        .SI(MESSAGE1[30]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[174]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_175_ ( .D(RESULT1[31]), 
        .SI(MESSAGE1[31]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[175]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_176_ ( .D(RESULT1[16]), 
        .SI(MESSAGE1[16]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[176]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_177_ ( .D(RESULT1[17]), 
        .SI(MESSAGE1[17]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[177]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_178_ ( .D(RESULT1[18]), 
        .SI(MESSAGE1[18]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[178]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_179_ ( .D(RESULT1[19]), 
        .SI(MESSAGE1[19]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[179]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_180_ ( .D(RESULT1[20]), 
        .SI(MESSAGE1[20]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[180]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_181_ ( .D(RESULT1[21]), 
        .SI(MESSAGE1[21]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[181]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_182_ ( .D(RESULT1[22]), 
        .SI(MESSAGE1[22]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[182]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_183_ ( .D(RESULT1[23]), 
        .SI(MESSAGE1[23]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[183]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_184_ ( .D(RESULT1[8]), 
        .SI(MESSAGE1[8]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[184]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_185_ ( .D(RESULT1[9]), 
        .SI(MESSAGE1[9]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[185]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_186_ ( .D(RESULT1[10]), 
        .SI(MESSAGE1[10]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[186]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_187_ ( .D(RESULT1[11]), 
        .SI(MESSAGE1[11]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[187]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_188_ ( .D(RESULT1[12]), 
        .SI(MESSAGE1[12]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[188]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_189_ ( .D(RESULT1[13]), 
        .SI(MESSAGE1[13]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[189]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_190_ ( .D(RESULT1[14]), 
        .SI(MESSAGE1[14]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[190]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_191_ ( .D(RESULT1[15]), 
        .SI(MESSAGE1[15]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[191]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_192_ ( .D(RESULT1[0]), 
        .SI(MESSAGE1[0]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[192]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_193_ ( .D(RESULT1[1]), 
        .SI(MESSAGE1[1]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[193]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_194_ ( .D(RESULT1[2]), 
        .SI(MESSAGE1[2]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[194]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_195_ ( .D(RESULT1[3]), 
        .SI(MESSAGE1[3]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[195]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_196_ ( .D(RESULT1[4]), 
        .SI(MESSAGE1[4]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[196]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_197_ ( .D(RESULT1[5]), 
        .SI(MESSAGE1[5]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[197]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_198_ ( .D(RESULT1[6]), 
        .SI(MESSAGE1[6]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[198]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_199_ ( .D(RESULT1[7]), 
        .SI(MESSAGE1[7]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[199]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_0_ ( .D(RESULT2[192]), 
        .SI(MESSAGE2[192]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[0]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_1_ ( .D(RESULT2[193]), 
        .SI(MESSAGE2[193]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[1]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_2_ ( .D(RESULT2[194]), 
        .SI(MESSAGE2[194]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[2]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_3_ ( .D(RESULT2[195]), 
        .SI(MESSAGE2[195]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[3]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_4_ ( .D(RESULT2[196]), 
        .SI(MESSAGE2[196]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[4]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_5_ ( .D(RESULT2[197]), 
        .SI(MESSAGE2[197]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[5]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_6_ ( .D(RESULT2[198]), 
        .SI(MESSAGE2[198]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[6]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_7_ ( .D(RESULT2[199]), 
        .SI(MESSAGE2[199]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[7]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_8_ ( .D(RESULT2[184]), 
        .SI(MESSAGE2[184]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[8]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_9_ ( .D(RESULT2[185]), 
        .SI(MESSAGE2[185]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[9]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_10_ ( .D(RESULT2[186]), 
        .SI(MESSAGE2[186]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[10]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_11_ ( .D(RESULT2[187]), 
        .SI(MESSAGE2[187]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[11]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_12_ ( .D(RESULT2[188]), 
        .SI(MESSAGE2[188]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[12]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_13_ ( .D(RESULT2[189]), 
        .SI(MESSAGE2[189]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[13]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_14_ ( .D(RESULT2[190]), 
        .SI(MESSAGE2[190]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[14]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_15_ ( .D(RESULT2[191]), 
        .SI(MESSAGE2[191]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[15]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_16_ ( .D(RESULT2[176]), 
        .SI(MESSAGE2[176]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[16]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_17_ ( .D(RESULT2[177]), 
        .SI(MESSAGE2[177]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[17]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_18_ ( .D(RESULT2[178]), 
        .SI(MESSAGE2[178]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[18]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_19_ ( .D(RESULT2[179]), 
        .SI(MESSAGE2[179]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[19]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_20_ ( .D(RESULT2[180]), 
        .SI(MESSAGE2[180]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[20]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_21_ ( .D(RESULT2[181]), 
        .SI(MESSAGE2[181]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[21]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_22_ ( .D(RESULT2[182]), 
        .SI(MESSAGE2[182]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[22]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_23_ ( .D(RESULT2[183]), 
        .SI(MESSAGE2[183]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[23]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_24_ ( .D(RESULT2[168]), 
        .SI(MESSAGE2[168]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[24]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_25_ ( .D(RESULT2[169]), 
        .SI(MESSAGE2[169]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[25]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_26_ ( .D(RESULT2[170]), 
        .SI(MESSAGE2[170]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[26]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_27_ ( .D(RESULT2[171]), 
        .SI(MESSAGE2[171]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[27]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_28_ ( .D(RESULT2[172]), 
        .SI(MESSAGE2[172]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[28]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_29_ ( .D(RESULT2[173]), 
        .SI(MESSAGE2[173]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[29]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_30_ ( .D(RESULT2[174]), 
        .SI(MESSAGE2[174]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[30]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_31_ ( .D(RESULT2[175]), 
        .SI(MESSAGE2[175]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[31]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_32_ ( .D(RESULT2[160]), 
        .SI(MESSAGE2[160]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[32]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_33_ ( .D(RESULT2[161]), 
        .SI(MESSAGE2[161]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[33]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_34_ ( .D(RESULT2[162]), 
        .SI(MESSAGE2[162]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[34]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_35_ ( .D(RESULT2[163]), 
        .SI(MESSAGE2[163]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[35]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_36_ ( .D(RESULT2[164]), 
        .SI(MESSAGE2[164]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[36]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_37_ ( .D(RESULT2[165]), 
        .SI(MESSAGE2[165]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[37]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_38_ ( .D(RESULT2[166]), 
        .SI(MESSAGE2[166]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[38]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_39_ ( .D(RESULT2[167]), 
        .SI(MESSAGE2[167]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[39]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_40_ ( .D(RESULT2[152]), 
        .SI(MESSAGE2[152]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[40]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_41_ ( .D(RESULT2[153]), 
        .SI(MESSAGE2[153]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[41]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_42_ ( .D(RESULT2[154]), 
        .SI(MESSAGE2[154]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[42]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_43_ ( .D(RESULT2[155]), 
        .SI(MESSAGE2[155]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[43]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_44_ ( .D(RESULT2[156]), 
        .SI(MESSAGE2[156]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[44]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_45_ ( .D(RESULT2[157]), 
        .SI(MESSAGE2[157]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[45]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_46_ ( .D(RESULT2[158]), 
        .SI(MESSAGE2[158]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[46]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_47_ ( .D(RESULT2[159]), 
        .SI(MESSAGE2[159]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[47]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_48_ ( .D(RESULT2[144]), 
        .SI(MESSAGE2[144]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[48]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_49_ ( .D(RESULT2[145]), 
        .SI(MESSAGE2[145]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[49]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_50_ ( .D(RESULT2[146]), 
        .SI(MESSAGE2[146]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[50]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_51_ ( .D(RESULT2[147]), 
        .SI(MESSAGE2[147]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[51]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_52_ ( .D(RESULT2[148]), 
        .SI(MESSAGE2[148]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[52]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_53_ ( .D(RESULT2[149]), 
        .SI(MESSAGE2[149]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[53]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_54_ ( .D(RESULT2[150]), 
        .SI(MESSAGE2[150]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[54]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_55_ ( .D(RESULT2[151]), 
        .SI(MESSAGE2[151]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[55]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_56_ ( .D(RESULT2[136]), 
        .SI(MESSAGE2[136]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[56]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_57_ ( .D(RESULT2[137]), 
        .SI(MESSAGE2[137]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[57]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_58_ ( .D(RESULT2[138]), 
        .SI(MESSAGE2[138]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[58]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_59_ ( .D(RESULT2[139]), 
        .SI(MESSAGE2[139]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[59]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_60_ ( .D(RESULT2[140]), 
        .SI(MESSAGE2[140]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[60]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_61_ ( .D(RESULT2[141]), 
        .SI(MESSAGE2[141]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[61]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_62_ ( .D(RESULT2[142]), 
        .SI(MESSAGE2[142]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[62]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_63_ ( .D(RESULT2[143]), 
        .SI(MESSAGE2[143]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[63]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_64_ ( .D(RESULT2[128]), 
        .SI(MESSAGE2[128]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[64]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_65_ ( .D(RESULT2[129]), 
        .SI(MESSAGE2[129]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[65]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_66_ ( .D(RESULT2[130]), 
        .SI(MESSAGE2[130]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[66]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_67_ ( .D(RESULT2[131]), 
        .SI(MESSAGE2[131]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[67]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_68_ ( .D(RESULT2[132]), 
        .SI(MESSAGE2[132]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[68]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_69_ ( .D(RESULT2[133]), 
        .SI(MESSAGE2[133]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[69]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_70_ ( .D(RESULT2[134]), 
        .SI(MESSAGE2[134]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[70]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_71_ ( .D(RESULT2[135]), 
        .SI(MESSAGE2[135]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[71]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_72_ ( .D(RESULT2[120]), 
        .SI(MESSAGE2[120]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[72]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_73_ ( .D(RESULT2[121]), 
        .SI(MESSAGE2[121]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[73]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_74_ ( .D(RESULT2[122]), 
        .SI(MESSAGE2[122]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[74]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_75_ ( .D(RESULT2[123]), 
        .SI(MESSAGE2[123]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[75]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_76_ ( .D(RESULT2[124]), 
        .SI(MESSAGE2[124]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[76]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_77_ ( .D(RESULT2[125]), 
        .SI(MESSAGE2[125]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[77]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_78_ ( .D(RESULT2[126]), 
        .SI(MESSAGE2[126]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[78]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_79_ ( .D(RESULT2[127]), 
        .SI(MESSAGE2[127]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[79]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_80_ ( .D(RESULT2[112]), 
        .SI(MESSAGE2[112]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[80]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_81_ ( .D(RESULT2[113]), 
        .SI(MESSAGE2[113]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[81]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_82_ ( .D(RESULT2[114]), 
        .SI(MESSAGE2[114]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[82]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_83_ ( .D(RESULT2[115]), 
        .SI(MESSAGE2[115]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[83]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_84_ ( .D(RESULT2[116]), 
        .SI(MESSAGE2[116]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[84]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_85_ ( .D(RESULT2[117]), 
        .SI(MESSAGE2[117]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[85]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_86_ ( .D(RESULT2[118]), 
        .SI(MESSAGE2[118]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[86]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_87_ ( .D(RESULT2[119]), 
        .SI(MESSAGE2[119]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[87]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_88_ ( .D(RESULT2[104]), 
        .SI(MESSAGE2[104]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[88]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_89_ ( .D(RESULT2[105]), 
        .SI(MESSAGE2[105]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[89]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_90_ ( .D(RESULT2[106]), 
        .SI(MESSAGE2[106]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[90]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_91_ ( .D(RESULT2[107]), 
        .SI(MESSAGE2[107]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[91]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_92_ ( .D(RESULT2[108]), 
        .SI(MESSAGE2[108]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[92]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_93_ ( .D(RESULT2[109]), 
        .SI(MESSAGE2[109]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[93]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_94_ ( .D(RESULT2[110]), 
        .SI(MESSAGE2[110]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[94]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_95_ ( .D(RESULT2[111]), 
        .SI(MESSAGE2[111]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[95]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_96_ ( .D(RESULT2[96]), 
        .SI(MESSAGE2[96]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[96]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_97_ ( .D(RESULT2[97]), 
        .SI(MESSAGE2[97]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[97]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_98_ ( .D(RESULT2[98]), 
        .SI(MESSAGE2[98]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[98]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_99_ ( .D(RESULT2[99]), 
        .SI(MESSAGE2[99]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[99]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_100_ ( .D(RESULT2[100]), 
        .SI(MESSAGE2[100]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[100]), .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_101_ ( .D(RESULT2[101]), 
        .SI(MESSAGE2[101]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[101]), .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_102_ ( .D(RESULT2[102]), 
        .SI(MESSAGE2[102]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[102]), .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_103_ ( .D(RESULT2[103]), 
        .SI(MESSAGE2[103]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[103]), .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_104_ ( .D(RESULT2[88]), 
        .SI(MESSAGE2[88]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[104]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_105_ ( .D(RESULT2[89]), 
        .SI(MESSAGE2[89]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[105]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_106_ ( .D(RESULT2[90]), 
        .SI(MESSAGE2[90]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[106]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_107_ ( .D(RESULT2[91]), 
        .SI(MESSAGE2[91]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[107]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_108_ ( .D(RESULT2[92]), 
        .SI(MESSAGE2[92]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[108]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_109_ ( .D(RESULT2[93]), 
        .SI(MESSAGE2[93]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[109]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_110_ ( .D(RESULT2[94]), 
        .SI(MESSAGE2[94]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[110]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_111_ ( .D(RESULT2[95]), 
        .SI(MESSAGE2[95]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[111]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_112_ ( .D(RESULT2[80]), 
        .SI(MESSAGE2[80]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[112]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_113_ ( .D(RESULT2[81]), 
        .SI(MESSAGE2[81]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[113]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_114_ ( .D(RESULT2[82]), 
        .SI(MESSAGE2[82]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[114]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_115_ ( .D(RESULT2[83]), 
        .SI(MESSAGE2[83]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[115]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_116_ ( .D(RESULT2[84]), 
        .SI(MESSAGE2[84]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[116]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_117_ ( .D(RESULT2[85]), 
        .SI(MESSAGE2[85]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[117]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_118_ ( .D(RESULT2[86]), 
        .SI(MESSAGE2[86]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[118]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_119_ ( .D(RESULT2[87]), 
        .SI(MESSAGE2[87]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[119]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_120_ ( .D(RESULT2[72]), 
        .SI(MESSAGE2[72]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[120]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_121_ ( .D(RESULT2[73]), 
        .SI(MESSAGE2[73]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[121]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_122_ ( .D(RESULT2[74]), 
        .SI(MESSAGE2[74]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[122]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_123_ ( .D(RESULT2[75]), 
        .SI(MESSAGE2[75]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[123]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_124_ ( .D(RESULT2[76]), 
        .SI(MESSAGE2[76]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[124]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_125_ ( .D(RESULT2[77]), 
        .SI(MESSAGE2[77]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[125]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_126_ ( .D(RESULT2[78]), 
        .SI(MESSAGE2[78]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[126]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_127_ ( .D(RESULT2[79]), 
        .SI(MESSAGE2[79]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[127]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_128_ ( .D(RESULT2[64]), 
        .SI(MESSAGE2[64]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[128]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_129_ ( .D(RESULT2[65]), 
        .SI(MESSAGE2[65]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[129]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_130_ ( .D(RESULT2[66]), 
        .SI(MESSAGE2[66]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[130]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_131_ ( .D(RESULT2[67]), 
        .SI(MESSAGE2[67]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[131]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_132_ ( .D(RESULT2[68]), 
        .SI(MESSAGE2[68]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[132]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_133_ ( .D(RESULT2[69]), 
        .SI(MESSAGE2[69]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[133]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_134_ ( .D(RESULT2[70]), 
        .SI(MESSAGE2[70]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[134]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_135_ ( .D(RESULT2[71]), 
        .SI(MESSAGE2[71]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[135]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_136_ ( .D(RESULT2[56]), 
        .SI(MESSAGE2[56]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[136]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_137_ ( .D(RESULT2[57]), 
        .SI(MESSAGE2[57]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[137]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_138_ ( .D(RESULT2[58]), 
        .SI(MESSAGE2[58]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[138]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_139_ ( .D(RESULT2[59]), 
        .SI(MESSAGE2[59]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[139]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_140_ ( .D(RESULT2[60]), 
        .SI(MESSAGE2[60]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[140]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_141_ ( .D(RESULT2[61]), 
        .SI(MESSAGE2[61]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[141]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_142_ ( .D(RESULT2[62]), 
        .SI(MESSAGE2[62]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[142]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_143_ ( .D(RESULT2[63]), 
        .SI(MESSAGE2[63]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[143]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_144_ ( .D(RESULT2[48]), 
        .SI(MESSAGE2[48]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[144]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_145_ ( .D(RESULT2[49]), 
        .SI(MESSAGE2[49]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[145]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_146_ ( .D(RESULT2[50]), 
        .SI(MESSAGE2[50]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[146]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_147_ ( .D(RESULT2[51]), 
        .SI(MESSAGE2[51]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[147]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_148_ ( .D(RESULT2[52]), 
        .SI(MESSAGE2[52]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[148]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_149_ ( .D(RESULT2[53]), 
        .SI(MESSAGE2[53]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[149]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_150_ ( .D(RESULT2[54]), 
        .SI(MESSAGE2[54]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[150]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_151_ ( .D(RESULT2[55]), 
        .SI(MESSAGE2[55]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[151]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_152_ ( .D(RESULT2[40]), 
        .SI(MESSAGE2[40]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[152]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_153_ ( .D(RESULT2[41]), 
        .SI(MESSAGE2[41]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[153]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_154_ ( .D(RESULT2[42]), 
        .SI(MESSAGE2[42]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[154]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_155_ ( .D(RESULT2[43]), 
        .SI(MESSAGE2[43]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[155]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_156_ ( .D(RESULT2[44]), 
        .SI(MESSAGE2[44]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[156]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_157_ ( .D(RESULT2[45]), 
        .SI(MESSAGE2[45]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[157]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_158_ ( .D(RESULT2[46]), 
        .SI(MESSAGE2[46]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[158]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_159_ ( .D(RESULT2[47]), 
        .SI(MESSAGE2[47]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[159]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_160_ ( .D(RESULT2[32]), 
        .SI(MESSAGE2[32]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[160]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_161_ ( .D(RESULT2[33]), 
        .SI(MESSAGE2[33]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[161]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_162_ ( .D(RESULT2[34]), 
        .SI(MESSAGE2[34]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[162]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_163_ ( .D(RESULT2[35]), 
        .SI(MESSAGE2[35]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[163]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_164_ ( .D(RESULT2[36]), 
        .SI(MESSAGE2[36]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[164]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_165_ ( .D(RESULT2[37]), 
        .SI(MESSAGE2[37]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[165]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_166_ ( .D(RESULT2[38]), 
        .SI(MESSAGE2[38]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[166]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_167_ ( .D(RESULT2[39]), 
        .SI(MESSAGE2[39]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[167]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_168_ ( .D(RESULT2[24]), 
        .SI(MESSAGE2[24]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[168]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_169_ ( .D(RESULT2[25]), 
        .SI(MESSAGE2[25]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[169]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_170_ ( .D(RESULT2[26]), 
        .SI(MESSAGE2[26]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[170]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_171_ ( .D(RESULT2[27]), 
        .SI(MESSAGE2[27]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[171]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_172_ ( .D(RESULT2[28]), 
        .SI(MESSAGE2[28]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[172]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_173_ ( .D(RESULT2[29]), 
        .SI(MESSAGE2[29]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[173]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_174_ ( .D(RESULT2[30]), 
        .SI(MESSAGE2[30]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[174]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_175_ ( .D(RESULT2[31]), 
        .SI(MESSAGE2[31]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[175]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_176_ ( .D(RESULT2[16]), 
        .SI(MESSAGE2[16]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[176]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_177_ ( .D(RESULT2[17]), 
        .SI(MESSAGE2[17]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[177]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_178_ ( .D(RESULT2[18]), 
        .SI(MESSAGE2[18]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[178]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_179_ ( .D(RESULT2[19]), 
        .SI(MESSAGE2[19]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[179]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_180_ ( .D(RESULT2[20]), 
        .SI(MESSAGE2[20]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[180]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_181_ ( .D(RESULT2[21]), 
        .SI(MESSAGE2[21]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[181]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_182_ ( .D(RESULT2[22]), 
        .SI(MESSAGE2[22]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[182]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_183_ ( .D(RESULT2[23]), 
        .SI(MESSAGE2[23]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[183]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_184_ ( .D(RESULT2[8]), 
        .SI(MESSAGE2[8]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[184]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_185_ ( .D(RESULT2[9]), 
        .SI(MESSAGE2[9]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[185]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_186_ ( .D(RESULT2[10]), 
        .SI(MESSAGE2[10]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[186]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_187_ ( .D(RESULT2[11]), 
        .SI(MESSAGE2[11]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[187]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_188_ ( .D(RESULT2[12]), 
        .SI(MESSAGE2[12]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[188]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_189_ ( .D(RESULT2[13]), 
        .SI(MESSAGE2[13]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[189]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_190_ ( .D(RESULT2[14]), 
        .SI(MESSAGE2[14]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[190]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_191_ ( .D(RESULT2[15]), 
        .SI(MESSAGE2[15]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[191]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_192_ ( .D(RESULT2[0]), 
        .SI(MESSAGE2[0]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[192]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_193_ ( .D(RESULT2[1]), 
        .SI(MESSAGE2[1]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[193]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_194_ ( .D(RESULT2[2]), 
        .SI(MESSAGE2[2]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[194]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_195_ ( .D(RESULT2[3]), 
        .SI(MESSAGE2[3]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[195]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_196_ ( .D(RESULT2[4]), 
        .SI(MESSAGE2[4]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[196]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_197_ ( .D(RESULT2[5]), 
        .SI(MESSAGE2[5]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[197]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_198_ ( .D(RESULT2[6]), 
        .SI(MESSAGE2[6]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[198]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_199_ ( .D(RESULT2[7]), 
        .SI(MESSAGE2[7]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[199]), 
        .QN() );
  XNOR2_X1 RoundFunction_T1_U400 ( .A(RoundFunction_STATE1[9]), .B(
        RoundFunction_T1_n400), .ZN(RoundFunction_TMP3_1[82]) );
  XNOR2_X1 RoundFunction_T1_U399 ( .A(RoundFunction_STATE1[99]), .B(
        RoundFunction_T1_n399), .ZN(RoundFunction_TMP3_1[22]) );
  XNOR2_X1 RoundFunction_T1_U398 ( .A(RoundFunction_STATE1[98]), .B(
        RoundFunction_T1_n398), .ZN(RoundFunction_TMP3_1[21]) );
  XNOR2_X1 RoundFunction_T1_U397 ( .A(RoundFunction_STATE1[97]), .B(
        RoundFunction_T1_n397), .ZN(RoundFunction_TMP3_1[20]) );
  XNOR2_X1 RoundFunction_T1_U396 ( .A(RoundFunction_STATE1[96]), .B(
        RoundFunction_T1_n396), .ZN(RoundFunction_TMP3_1[19]) );
  XNOR2_X1 RoundFunction_T1_U395 ( .A(RoundFunction_STATE1[95]), .B(
        RoundFunction_T1_n395), .ZN(RoundFunction_TMP3_1[137]) );
  XNOR2_X1 RoundFunction_T1_U394 ( .A(RoundFunction_STATE1[94]), .B(
        RoundFunction_T1_n394), .ZN(RoundFunction_TMP3_1[136]) );
  XNOR2_X1 RoundFunction_T1_U393 ( .A(RoundFunction_STATE1[93]), .B(
        RoundFunction_T1_n393), .ZN(RoundFunction_TMP3_1[143]) );
  XNOR2_X1 RoundFunction_T1_U392 ( .A(RoundFunction_STATE1[92]), .B(
        RoundFunction_T1_n392), .ZN(RoundFunction_TMP3_1[142]) );
  XNOR2_X1 RoundFunction_T1_U391 ( .A(RoundFunction_STATE1[91]), .B(
        RoundFunction_T1_n391), .ZN(RoundFunction_TMP3_1[141]) );
  XNOR2_X1 RoundFunction_T1_U390 ( .A(RoundFunction_STATE1[90]), .B(
        RoundFunction_T1_n390), .ZN(RoundFunction_TMP3_1[140]) );
  XNOR2_X1 RoundFunction_T1_U389 ( .A(RoundFunction_STATE1[8]), .B(
        RoundFunction_T1_n389), .ZN(RoundFunction_TMP3_1[81]) );
  XNOR2_X1 RoundFunction_T1_U388 ( .A(RoundFunction_STATE1[89]), .B(
        RoundFunction_T1_n400), .ZN(RoundFunction_TMP3_1[139]) );
  XNOR2_X1 RoundFunction_T1_U387 ( .A(RoundFunction_STATE1[88]), .B(
        RoundFunction_T1_n389), .ZN(RoundFunction_TMP3_1[138]) );
  XNOR2_X1 RoundFunction_T1_U386 ( .A(RoundFunction_STATE1[87]), .B(
        RoundFunction_T1_n388), .ZN(RoundFunction_TMP3_1[58]) );
  XNOR2_X1 RoundFunction_T1_U385 ( .A(RoundFunction_STATE1[86]), .B(
        RoundFunction_T1_n387), .ZN(RoundFunction_TMP3_1[57]) );
  XNOR2_X1 RoundFunction_T1_U384 ( .A(RoundFunction_STATE1[85]), .B(
        RoundFunction_T1_n386), .ZN(RoundFunction_TMP3_1[56]) );
  XNOR2_X1 RoundFunction_T1_U383 ( .A(RoundFunction_STATE1[84]), .B(
        RoundFunction_T1_n385), .ZN(RoundFunction_TMP3_1[63]) );
  XNOR2_X1 RoundFunction_T1_U382 ( .A(RoundFunction_STATE1[83]), .B(
        RoundFunction_T1_n384), .ZN(RoundFunction_TMP3_1[62]) );
  XNOR2_X1 RoundFunction_T1_U381 ( .A(RoundFunction_STATE1[82]), .B(
        RoundFunction_T1_n383), .ZN(RoundFunction_TMP3_1[61]) );
  XNOR2_X1 RoundFunction_T1_U380 ( .A(RoundFunction_STATE1[81]), .B(
        RoundFunction_T1_n382), .ZN(RoundFunction_TMP3_1[60]) );
  XNOR2_X1 RoundFunction_T1_U379 ( .A(RoundFunction_STATE1[80]), .B(
        RoundFunction_T1_n381), .ZN(RoundFunction_TMP3_1[59]) );
  XNOR2_X1 RoundFunction_T1_U378 ( .A(RoundFunction_STATE1[7]), .B(
        RoundFunction_T1_n388), .ZN(RoundFunction_TMP3_1[7]) );
  XNOR2_X1 RoundFunction_T1_U377 ( .A(RoundFunction_STATE1[79]), .B(
        RoundFunction_T1_n380), .ZN(RoundFunction_TMP3_1[51]) );
  XNOR2_X1 RoundFunction_T1_U376 ( .A(RoundFunction_STATE1[78]), .B(
        RoundFunction_T1_n379), .ZN(RoundFunction_TMP3_1[50]) );
  XNOR2_X1 RoundFunction_T1_U375 ( .A(RoundFunction_STATE1[77]), .B(
        RoundFunction_T1_n378), .ZN(RoundFunction_TMP3_1[49]) );
  XNOR2_X1 RoundFunction_T1_U374 ( .A(RoundFunction_STATE1[76]), .B(
        RoundFunction_T1_n377), .ZN(RoundFunction_TMP3_1[48]) );
  XNOR2_X1 RoundFunction_T1_U373 ( .A(RoundFunction_STATE1[75]), .B(
        RoundFunction_T1_n376), .ZN(RoundFunction_TMP3_1[55]) );
  XNOR2_X1 RoundFunction_T1_U372 ( .A(RoundFunction_STATE1[74]), .B(
        RoundFunction_T1_n375), .ZN(RoundFunction_TMP3_1[54]) );
  XNOR2_X1 RoundFunction_T1_U371 ( .A(RoundFunction_STATE1[73]), .B(
        RoundFunction_T1_n374), .ZN(RoundFunction_TMP3_1[53]) );
  XNOR2_X1 RoundFunction_T1_U370 ( .A(RoundFunction_STATE1[72]), .B(
        RoundFunction_T1_n373), .ZN(RoundFunction_TMP3_1[52]) );
  XNOR2_X1 RoundFunction_T1_U369 ( .A(RoundFunction_STATE1[71]), .B(
        RoundFunction_T1_n372), .ZN(RoundFunction_TMP3_1[174]) );
  XNOR2_X1 RoundFunction_T1_U368 ( .A(RoundFunction_STATE1[70]), .B(
        RoundFunction_T1_n371), .ZN(RoundFunction_TMP3_1[173]) );
  XNOR2_X1 RoundFunction_T1_U367 ( .A(RoundFunction_STATE1[6]), .B(
        RoundFunction_T1_n387), .ZN(RoundFunction_TMP3_1[6]) );
  XNOR2_X1 RoundFunction_T1_U366 ( .A(RoundFunction_STATE1[69]), .B(
        RoundFunction_T1_n370), .ZN(RoundFunction_TMP3_1[172]) );
  XNOR2_X1 RoundFunction_T1_U365 ( .A(RoundFunction_STATE1[68]), .B(
        RoundFunction_T1_n369), .ZN(RoundFunction_TMP3_1[171]) );
  XNOR2_X1 RoundFunction_T1_U364 ( .A(RoundFunction_STATE1[67]), .B(
        RoundFunction_T1_n368), .ZN(RoundFunction_TMP3_1[170]) );
  XNOR2_X1 RoundFunction_T1_U363 ( .A(RoundFunction_STATE1[66]), .B(
        RoundFunction_T1_n367), .ZN(RoundFunction_TMP3_1[169]) );
  XNOR2_X1 RoundFunction_T1_U362 ( .A(RoundFunction_STATE1[65]), .B(
        RoundFunction_T1_n366), .ZN(RoundFunction_TMP3_1[168]) );
  XNOR2_X1 RoundFunction_T1_U361 ( .A(RoundFunction_STATE1[64]), .B(
        RoundFunction_T1_n365), .ZN(RoundFunction_TMP3_1[175]) );
  XNOR2_X1 RoundFunction_T1_U360 ( .A(RoundFunction_STATE1[63]), .B(
        RoundFunction_T1_n364), .ZN(RoundFunction_TMP3_1[93]) );
  XNOR2_X1 RoundFunction_T1_U359 ( .A(RoundFunction_STATE1[62]), .B(
        RoundFunction_T1_n363), .ZN(RoundFunction_TMP3_1[92]) );
  XNOR2_X1 RoundFunction_T1_U358 ( .A(RoundFunction_STATE1[61]), .B(
        RoundFunction_T1_n362), .ZN(RoundFunction_TMP3_1[91]) );
  XNOR2_X1 RoundFunction_T1_U357 ( .A(RoundFunction_STATE1[60]), .B(
        RoundFunction_T1_n361), .ZN(RoundFunction_TMP3_1[90]) );
  XNOR2_X1 RoundFunction_T1_U356 ( .A(RoundFunction_STATE1[5]), .B(
        RoundFunction_T1_n386), .ZN(RoundFunction_TMP3_1[5]) );
  XNOR2_X1 RoundFunction_T1_U355 ( .A(RoundFunction_STATE1[59]), .B(
        RoundFunction_T1_n399), .ZN(RoundFunction_TMP3_1[89]) );
  XNOR2_X1 RoundFunction_T1_U354 ( .A(RoundFunction_STATE1[58]), .B(
        RoundFunction_T1_n398), .ZN(RoundFunction_TMP3_1[88]) );
  XNOR2_X1 RoundFunction_T1_U353 ( .A(RoundFunction_STATE1[57]), .B(
        RoundFunction_T1_n397), .ZN(RoundFunction_TMP3_1[95]) );
  XNOR2_X1 RoundFunction_T1_U352 ( .A(RoundFunction_STATE1[56]), .B(
        RoundFunction_T1_n396), .ZN(RoundFunction_TMP3_1[94]) );
  XNOR2_X1 RoundFunction_T1_U351 ( .A(RoundFunction_STATE1[55]), .B(
        RoundFunction_T1_n395), .ZN(RoundFunction_TMP3_1[11]) );
  XNOR2_X1 RoundFunction_T1_U350 ( .A(RoundFunction_STATE1[54]), .B(
        RoundFunction_T1_n394), .ZN(RoundFunction_TMP3_1[10]) );
  XNOR2_X1 RoundFunction_T1_U349 ( .A(RoundFunction_STATE1[53]), .B(
        RoundFunction_T1_n393), .ZN(RoundFunction_TMP3_1[9]) );
  XNOR2_X1 RoundFunction_T1_U348 ( .A(RoundFunction_STATE1[52]), .B(
        RoundFunction_T1_n392), .ZN(RoundFunction_TMP3_1[8]) );
  XNOR2_X1 RoundFunction_T1_U347 ( .A(RoundFunction_STATE1[51]), .B(
        RoundFunction_T1_n391), .ZN(RoundFunction_TMP3_1[15]) );
  XNOR2_X1 RoundFunction_T1_U346 ( .A(RoundFunction_STATE1[50]), .B(
        RoundFunction_T1_n390), .ZN(RoundFunction_TMP3_1[14]) );
  XNOR2_X1 RoundFunction_T1_U345 ( .A(RoundFunction_STATE1[4]), .B(
        RoundFunction_T1_n385), .ZN(RoundFunction_TMP3_1[4]) );
  XNOR2_X1 RoundFunction_T1_U344 ( .A(RoundFunction_STATE1[49]), .B(
        RoundFunction_T1_n400), .ZN(RoundFunction_TMP3_1[13]) );
  XNOR2_X1 RoundFunction_T1_U343 ( .A(RoundFunction_STATE1[48]), .B(
        RoundFunction_T1_n389), .ZN(RoundFunction_TMP3_1[12]) );
  XNOR2_X1 RoundFunction_T1_U342 ( .A(RoundFunction_STATE1[47]), .B(
        RoundFunction_T1_n388), .ZN(RoundFunction_TMP3_1[131]) );
  XNOR2_X1 RoundFunction_T1_U341 ( .A(RoundFunction_STATE1[46]), .B(
        RoundFunction_T1_n387), .ZN(RoundFunction_TMP3_1[130]) );
  XNOR2_X1 RoundFunction_T1_U340 ( .A(RoundFunction_STATE1[45]), .B(
        RoundFunction_T1_n386), .ZN(RoundFunction_TMP3_1[129]) );
  XNOR2_X1 RoundFunction_T1_U339 ( .A(RoundFunction_STATE1[44]), .B(
        RoundFunction_T1_n385), .ZN(RoundFunction_TMP3_1[128]) );
  XNOR2_X1 RoundFunction_T1_U338 ( .A(RoundFunction_STATE1[43]), .B(
        RoundFunction_T1_n384), .ZN(RoundFunction_TMP3_1[135]) );
  XNOR2_X1 RoundFunction_T1_U337 ( .A(RoundFunction_STATE1[42]), .B(
        RoundFunction_T1_n383), .ZN(RoundFunction_TMP3_1[134]) );
  XNOR2_X1 RoundFunction_T1_U336 ( .A(RoundFunction_STATE1[41]), .B(
        RoundFunction_T1_n382), .ZN(RoundFunction_TMP3_1[133]) );
  XNOR2_X1 RoundFunction_T1_U335 ( .A(RoundFunction_STATE1[40]), .B(
        RoundFunction_T1_n381), .ZN(RoundFunction_TMP3_1[132]) );
  XNOR2_X1 RoundFunction_T1_U334 ( .A(RoundFunction_STATE1[3]), .B(
        RoundFunction_T1_n384), .ZN(RoundFunction_TMP3_1[3]) );
  XNOR2_X1 RoundFunction_T1_U333 ( .A(RoundFunction_STATE1[39]), .B(
        RoundFunction_T1_n380), .ZN(RoundFunction_TMP3_1[122]) );
  XNOR2_X1 RoundFunction_T1_U332 ( .A(RoundFunction_STATE1[38]), .B(
        RoundFunction_T1_n379), .ZN(RoundFunction_TMP3_1[121]) );
  XNOR2_X1 RoundFunction_T1_U331 ( .A(RoundFunction_STATE1[37]), .B(
        RoundFunction_T1_n378), .ZN(RoundFunction_TMP3_1[120]) );
  XNOR2_X1 RoundFunction_T1_U330 ( .A(RoundFunction_STATE1[36]), .B(
        RoundFunction_T1_n377), .ZN(RoundFunction_TMP3_1[127]) );
  XNOR2_X1 RoundFunction_T1_U329 ( .A(RoundFunction_STATE1[35]), .B(
        RoundFunction_T1_n376), .ZN(RoundFunction_TMP3_1[126]) );
  XNOR2_X1 RoundFunction_T1_U328 ( .A(RoundFunction_STATE1[34]), .B(
        RoundFunction_T1_n375), .ZN(RoundFunction_TMP3_1[125]) );
  XNOR2_X1 RoundFunction_T1_U327 ( .A(RoundFunction_STATE1[33]), .B(
        RoundFunction_T1_n374), .ZN(RoundFunction_TMP3_1[124]) );
  XNOR2_X1 RoundFunction_T1_U326 ( .A(RoundFunction_STATE1[32]), .B(
        RoundFunction_T1_n373), .ZN(RoundFunction_TMP3_1[123]) );
  XNOR2_X1 RoundFunction_T1_U325 ( .A(RoundFunction_STATE1[31]), .B(
        RoundFunction_T1_n372), .ZN(RoundFunction_TMP3_1[43]) );
  XNOR2_X1 RoundFunction_T1_U324 ( .A(RoundFunction_STATE1[30]), .B(
        RoundFunction_T1_n371), .ZN(RoundFunction_TMP3_1[42]) );
  XNOR2_X1 RoundFunction_T1_U323 ( .A(RoundFunction_STATE1[2]), .B(
        RoundFunction_T1_n383), .ZN(RoundFunction_TMP3_1[2]) );
  XNOR2_X1 RoundFunction_T1_U322 ( .A(RoundFunction_STATE1[29]), .B(
        RoundFunction_T1_n370), .ZN(RoundFunction_TMP3_1[41]) );
  XNOR2_X1 RoundFunction_T1_U321 ( .A(RoundFunction_STATE1[28]), .B(
        RoundFunction_T1_n369), .ZN(RoundFunction_TMP3_1[40]) );
  XNOR2_X1 RoundFunction_T1_U320 ( .A(RoundFunction_STATE1[27]), .B(
        RoundFunction_T1_n368), .ZN(RoundFunction_TMP3_1[47]) );
  XNOR2_X1 RoundFunction_T1_U319 ( .A(RoundFunction_STATE1[26]), .B(
        RoundFunction_T1_n367), .ZN(RoundFunction_TMP3_1[46]) );
  XNOR2_X1 RoundFunction_T1_U318 ( .A(RoundFunction_STATE1[25]), .B(
        RoundFunction_T1_n366), .ZN(RoundFunction_TMP3_1[45]) );
  XNOR2_X1 RoundFunction_T1_U317 ( .A(RoundFunction_STATE1[24]), .B(
        RoundFunction_T1_n365), .ZN(RoundFunction_TMP3_1[44]) );
  XNOR2_X1 RoundFunction_T1_U316 ( .A(RoundFunction_STATE1[23]), .B(
        RoundFunction_T1_n364), .ZN(RoundFunction_TMP3_1[165]) );
  XNOR2_X1 RoundFunction_T1_U315 ( .A(RoundFunction_STATE1[22]), .B(
        RoundFunction_T1_n363), .ZN(RoundFunction_TMP3_1[164]) );
  XNOR2_X1 RoundFunction_T1_U314 ( .A(RoundFunction_STATE1[21]), .B(
        RoundFunction_T1_n362), .ZN(RoundFunction_TMP3_1[163]) );
  XNOR2_X1 RoundFunction_T1_U313 ( .A(RoundFunction_STATE1[20]), .B(
        RoundFunction_T1_n361), .ZN(RoundFunction_TMP3_1[162]) );
  XNOR2_X1 RoundFunction_T1_U312 ( .A(RoundFunction_STATE1[1]), .B(
        RoundFunction_T1_n382), .ZN(RoundFunction_TMP3_1[1]) );
  XNOR2_X1 RoundFunction_T1_U311 ( .A(RoundFunction_STATE1[19]), .B(
        RoundFunction_T1_n399), .ZN(RoundFunction_TMP3_1[161]) );
  XNOR2_X1 RoundFunction_T1_U310 ( .A(RoundFunction_STATE1[199]), .B(
        RoundFunction_T1_n380), .ZN(RoundFunction_TMP3_1[37]) );
  XNOR2_X1 RoundFunction_T1_U309 ( .A(RoundFunction_STATE1[198]), .B(
        RoundFunction_T1_n379), .ZN(RoundFunction_TMP3_1[36]) );
  XNOR2_X1 RoundFunction_T1_U308 ( .A(RoundFunction_STATE1[197]), .B(
        RoundFunction_T1_n378), .ZN(RoundFunction_TMP3_1[35]) );
  XNOR2_X1 RoundFunction_T1_U307 ( .A(RoundFunction_STATE1[196]), .B(
        RoundFunction_T1_n377), .ZN(RoundFunction_TMP3_1[34]) );
  XNOR2_X1 RoundFunction_T1_U306 ( .A(RoundFunction_STATE1[195]), .B(
        RoundFunction_T1_n376), .ZN(RoundFunction_TMP3_1[33]) );
  XNOR2_X1 RoundFunction_T1_U305 ( .A(RoundFunction_STATE1[194]), .B(
        RoundFunction_T1_n375), .ZN(RoundFunction_TMP3_1[32]) );
  XNOR2_X1 RoundFunction_T1_U304 ( .A(RoundFunction_STATE1[193]), .B(
        RoundFunction_T1_n374), .ZN(RoundFunction_TMP3_1[39]) );
  XNOR2_X1 RoundFunction_T1_U303 ( .A(RoundFunction_STATE1[192]), .B(
        RoundFunction_T1_n373), .ZN(RoundFunction_TMP3_1[38]) );
  XNOR2_X1 RoundFunction_T1_U302 ( .A(RoundFunction_STATE1[191]), .B(
        RoundFunction_T1_n372), .ZN(RoundFunction_TMP3_1[159]) );
  XNOR2_X1 RoundFunction_T1_U301 ( .A(RoundFunction_STATE1[190]), .B(
        RoundFunction_T1_n371), .ZN(RoundFunction_TMP3_1[158]) );
  XNOR2_X1 RoundFunction_T1_U300 ( .A(RoundFunction_STATE1[18]), .B(
        RoundFunction_T1_n398), .ZN(RoundFunction_TMP3_1[160]) );
  XNOR2_X1 RoundFunction_T1_U299 ( .A(RoundFunction_STATE1[189]), .B(
        RoundFunction_T1_n370), .ZN(RoundFunction_TMP3_1[157]) );
  XNOR2_X1 RoundFunction_T1_U298 ( .A(RoundFunction_STATE1[188]), .B(
        RoundFunction_T1_n369), .ZN(RoundFunction_TMP3_1[156]) );
  XNOR2_X1 RoundFunction_T1_U297 ( .A(RoundFunction_STATE1[187]), .B(
        RoundFunction_T1_n368), .ZN(RoundFunction_TMP3_1[155]) );
  XNOR2_X1 RoundFunction_T1_U296 ( .A(RoundFunction_STATE1[186]), .B(
        RoundFunction_T1_n367), .ZN(RoundFunction_TMP3_1[154]) );
  XNOR2_X1 RoundFunction_T1_U295 ( .A(RoundFunction_STATE1[185]), .B(
        RoundFunction_T1_n366), .ZN(RoundFunction_TMP3_1[153]) );
  XNOR2_X1 RoundFunction_T1_U294 ( .A(RoundFunction_STATE1[184]), .B(
        RoundFunction_T1_n365), .ZN(RoundFunction_TMP3_1[152]) );
  XNOR2_X1 RoundFunction_T1_U293 ( .A(RoundFunction_STATE1[183]), .B(
        RoundFunction_T1_n364), .ZN(RoundFunction_TMP3_1[76]) );
  XNOR2_X1 RoundFunction_T1_U292 ( .A(RoundFunction_STATE1[182]), .B(
        RoundFunction_T1_n363), .ZN(RoundFunction_TMP3_1[75]) );
  XNOR2_X1 RoundFunction_T1_U291 ( .A(RoundFunction_STATE1[181]), .B(
        RoundFunction_T1_n362), .ZN(RoundFunction_TMP3_1[74]) );
  XNOR2_X1 RoundFunction_T1_U290 ( .A(RoundFunction_STATE1[180]), .B(
        RoundFunction_T1_n361), .ZN(RoundFunction_TMP3_1[73]) );
  XNOR2_X1 RoundFunction_T1_U289 ( .A(RoundFunction_STATE1[17]), .B(
        RoundFunction_T1_n397), .ZN(RoundFunction_TMP3_1[167]) );
  XNOR2_X1 RoundFunction_T1_U288 ( .A(RoundFunction_STATE1[179]), .B(
        RoundFunction_T1_n399), .ZN(RoundFunction_TMP3_1[72]) );
  XNOR2_X1 RoundFunction_T1_U287 ( .A(RoundFunction_STATE1[178]), .B(
        RoundFunction_T1_n398), .ZN(RoundFunction_TMP3_1[79]) );
  XNOR2_X1 RoundFunction_T1_U286 ( .A(RoundFunction_STATE1[177]), .B(
        RoundFunction_T1_n397), .ZN(RoundFunction_TMP3_1[78]) );
  XNOR2_X1 RoundFunction_T1_U285 ( .A(RoundFunction_STATE1[176]), .B(
        RoundFunction_T1_n396), .ZN(RoundFunction_TMP3_1[77]) );
  XNOR2_X1 RoundFunction_T1_U284 ( .A(RoundFunction_STATE1[175]), .B(
        RoundFunction_T1_n395), .ZN(RoundFunction_TMP3_1[193]) );
  XNOR2_X1 RoundFunction_T1_U283 ( .A(RoundFunction_STATE1[174]), .B(
        RoundFunction_T1_n394), .ZN(RoundFunction_TMP3_1[192]) );
  XNOR2_X1 RoundFunction_T1_U282 ( .A(RoundFunction_STATE1[173]), .B(
        RoundFunction_T1_n393), .ZN(RoundFunction_TMP3_1[199]) );
  XNOR2_X1 RoundFunction_T1_U281 ( .A(RoundFunction_STATE1[172]), .B(
        RoundFunction_T1_n392), .ZN(RoundFunction_TMP3_1[198]) );
  XNOR2_X1 RoundFunction_T1_U280 ( .A(RoundFunction_STATE1[171]), .B(
        RoundFunction_T1_n391), .ZN(RoundFunction_TMP3_1[197]) );
  XNOR2_X1 RoundFunction_T1_U279 ( .A(RoundFunction_STATE1[170]), .B(
        RoundFunction_T1_n390), .ZN(RoundFunction_TMP3_1[196]) );
  XNOR2_X1 RoundFunction_T1_U278 ( .A(RoundFunction_STATE1[16]), .B(
        RoundFunction_T1_n396), .ZN(RoundFunction_TMP3_1[166]) );
  XNOR2_X1 RoundFunction_T1_U277 ( .A(RoundFunction_STATE1[169]), .B(
        RoundFunction_T1_n400), .ZN(RoundFunction_TMP3_1[195]) );
  XNOR2_X1 RoundFunction_T1_U276 ( .A(RoundFunction_STATE1[168]), .B(
        RoundFunction_T1_n389), .ZN(RoundFunction_TMP3_1[194]) );
  XNOR2_X1 RoundFunction_T1_U275 ( .A(RoundFunction_STATE1[167]), .B(
        RoundFunction_T1_n388), .ZN(RoundFunction_TMP3_1[113]) );
  XNOR2_X1 RoundFunction_T1_U274 ( .A(RoundFunction_STATE1[166]), .B(
        RoundFunction_T1_n387), .ZN(RoundFunction_TMP3_1[112]) );
  XNOR2_X1 RoundFunction_T1_U273 ( .A(RoundFunction_STATE1[165]), .B(
        RoundFunction_T1_n386), .ZN(RoundFunction_TMP3_1[119]) );
  XNOR2_X1 RoundFunction_T1_U272 ( .A(RoundFunction_STATE1[164]), .B(
        RoundFunction_T1_n385), .ZN(RoundFunction_TMP3_1[118]) );
  XNOR2_X1 RoundFunction_T1_U271 ( .A(RoundFunction_STATE1[163]), .B(
        RoundFunction_T1_n384), .ZN(RoundFunction_TMP3_1[117]) );
  XNOR2_X1 RoundFunction_T1_U270 ( .A(RoundFunction_STATE1[162]), .B(
        RoundFunction_T1_n383), .ZN(RoundFunction_TMP3_1[116]) );
  XNOR2_X1 RoundFunction_T1_U269 ( .A(RoundFunction_STATE1[161]), .B(
        RoundFunction_T1_n382), .ZN(RoundFunction_TMP3_1[115]) );
  XNOR2_X1 RoundFunction_T1_U268 ( .A(RoundFunction_STATE1[160]), .B(
        RoundFunction_T1_n381), .ZN(RoundFunction_TMP3_1[114]) );
  XNOR2_X1 RoundFunction_T1_U267 ( .A(RoundFunction_STATE1[15]), .B(
        RoundFunction_T1_n395), .ZN(RoundFunction_TMP3_1[80]) );
  XNOR2_X1 RoundFunction_T1_U266 ( .A(RoundFunction_STATE1[159]), .B(
        RoundFunction_T1_n380), .ZN(RoundFunction_TMP3_1[111]) );
  XNOR2_X1 RoundFunction_T1_U265 ( .A(RoundFunction_STATE1[158]), .B(
        RoundFunction_T1_n379), .ZN(RoundFunction_TMP3_1[110]) );
  XNOR2_X1 RoundFunction_T1_U264 ( .A(RoundFunction_STATE1[157]), .B(
        RoundFunction_T1_n378), .ZN(RoundFunction_TMP3_1[109]) );
  XNOR2_X1 RoundFunction_T1_U263 ( .A(RoundFunction_STATE1[156]), .B(
        RoundFunction_T1_n377), .ZN(RoundFunction_TMP3_1[108]) );
  XNOR2_X1 RoundFunction_T1_U262 ( .A(RoundFunction_STATE1[155]), .B(
        RoundFunction_T1_n376), .ZN(RoundFunction_TMP3_1[107]) );
  XNOR2_X1 RoundFunction_T1_U261 ( .A(RoundFunction_STATE1[154]), .B(
        RoundFunction_T1_n375), .ZN(RoundFunction_TMP3_1[106]) );
  XNOR2_X1 RoundFunction_T1_U260 ( .A(RoundFunction_STATE1[153]), .B(
        RoundFunction_T1_n374), .ZN(RoundFunction_TMP3_1[105]) );
  XNOR2_X1 RoundFunction_T1_U259 ( .A(RoundFunction_STATE1[152]), .B(
        RoundFunction_T1_n373), .ZN(RoundFunction_TMP3_1[104]) );
  XNOR2_X1 RoundFunction_T1_U258 ( .A(RoundFunction_STATE1[151]), .B(
        RoundFunction_T1_n372), .ZN(RoundFunction_TMP3_1[28]) );
  XNOR2_X1 RoundFunction_T1_U257 ( .A(RoundFunction_STATE1[150]), .B(
        RoundFunction_T1_n371), .ZN(RoundFunction_TMP3_1[27]) );
  XNOR2_X1 RoundFunction_T1_U256 ( .A(RoundFunction_STATE1[14]), .B(
        RoundFunction_T1_n394), .ZN(RoundFunction_TMP3_1[87]) );
  XNOR2_X1 RoundFunction_T1_U255 ( .A(RoundFunction_STATE1[149]), .B(
        RoundFunction_T1_n370), .ZN(RoundFunction_TMP3_1[26]) );
  XNOR2_X1 RoundFunction_T1_U254 ( .A(RoundFunction_STATE1[148]), .B(
        RoundFunction_T1_n369), .ZN(RoundFunction_TMP3_1[25]) );
  XNOR2_X1 RoundFunction_T1_U253 ( .A(RoundFunction_STATE1[147]), .B(
        RoundFunction_T1_n368), .ZN(RoundFunction_TMP3_1[24]) );
  XNOR2_X1 RoundFunction_T1_U252 ( .A(RoundFunction_STATE1[146]), .B(
        RoundFunction_T1_n367), .ZN(RoundFunction_TMP3_1[31]) );
  XNOR2_X1 RoundFunction_T1_U251 ( .A(RoundFunction_STATE1[145]), .B(
        RoundFunction_T1_n366), .ZN(RoundFunction_TMP3_1[30]) );
  XNOR2_X1 RoundFunction_T1_U250 ( .A(RoundFunction_STATE1[144]), .B(
        RoundFunction_T1_n365), .ZN(RoundFunction_TMP3_1[29]) );
  XNOR2_X1 RoundFunction_T1_U249 ( .A(RoundFunction_STATE1[143]), .B(
        RoundFunction_T1_n364), .ZN(RoundFunction_TMP3_1[150]) );
  XNOR2_X1 RoundFunction_T1_U248 ( .A(RoundFunction_STATE1[142]), .B(
        RoundFunction_T1_n363), .ZN(RoundFunction_TMP3_1[149]) );
  XNOR2_X1 RoundFunction_T1_U247 ( .A(RoundFunction_STATE1[141]), .B(
        RoundFunction_T1_n362), .ZN(RoundFunction_TMP3_1[148]) );
  XNOR2_X1 RoundFunction_T1_U246 ( .A(RoundFunction_STATE1[140]), .B(
        RoundFunction_T1_n361), .ZN(RoundFunction_TMP3_1[147]) );
  XNOR2_X1 RoundFunction_T1_U245 ( .A(RoundFunction_STATE1[13]), .B(
        RoundFunction_T1_n393), .ZN(RoundFunction_TMP3_1[86]) );
  XNOR2_X1 RoundFunction_T1_U244 ( .A(RoundFunction_STATE1[139]), .B(
        RoundFunction_T1_n399), .ZN(RoundFunction_TMP3_1[146]) );
  XNOR2_X1 RoundFunction_T1_U243 ( .A(RoundFunction_T1_n360), .B(
        RoundFunction_T1_n359), .ZN(RoundFunction_T1_n399) );
  XNOR2_X1 RoundFunction_T1_U242 ( .A(RoundFunction_STATE1[138]), .B(
        RoundFunction_T1_n398), .ZN(RoundFunction_TMP3_1[145]) );
  XNOR2_X1 RoundFunction_T1_U241 ( .A(RoundFunction_T1_n358), .B(
        RoundFunction_T1_n357), .ZN(RoundFunction_T1_n398) );
  XNOR2_X1 RoundFunction_T1_U240 ( .A(RoundFunction_STATE1[137]), .B(
        RoundFunction_T1_n397), .ZN(RoundFunction_TMP3_1[144]) );
  XNOR2_X1 RoundFunction_T1_U239 ( .A(RoundFunction_T1_n356), .B(
        RoundFunction_T1_n355), .ZN(RoundFunction_T1_n397) );
  XNOR2_X1 RoundFunction_T1_U238 ( .A(RoundFunction_STATE1[136]), .B(
        RoundFunction_T1_n396), .ZN(RoundFunction_TMP3_1[151]) );
  XNOR2_X1 RoundFunction_T1_U237 ( .A(RoundFunction_T1_n354), .B(
        RoundFunction_T1_n353), .ZN(RoundFunction_T1_n396) );
  XNOR2_X1 RoundFunction_T1_U236 ( .A(RoundFunction_STATE1[135]), .B(
        RoundFunction_T1_n395), .ZN(RoundFunction_TMP3_1[68]) );
  XNOR2_X1 RoundFunction_T1_U235 ( .A(RoundFunction_T1_n352), .B(
        RoundFunction_T1_n351), .ZN(RoundFunction_T1_n395) );
  XNOR2_X1 RoundFunction_T1_U234 ( .A(RoundFunction_STATE1[134]), .B(
        RoundFunction_T1_n394), .ZN(RoundFunction_TMP3_1[67]) );
  XNOR2_X1 RoundFunction_T1_U233 ( .A(RoundFunction_T1_n350), .B(
        RoundFunction_T1_n349), .ZN(RoundFunction_T1_n394) );
  XNOR2_X1 RoundFunction_T1_U232 ( .A(RoundFunction_STATE1[133]), .B(
        RoundFunction_T1_n393), .ZN(RoundFunction_TMP3_1[66]) );
  XNOR2_X1 RoundFunction_T1_U231 ( .A(RoundFunction_T1_n348), .B(
        RoundFunction_T1_n347), .ZN(RoundFunction_T1_n393) );
  XNOR2_X1 RoundFunction_T1_U230 ( .A(RoundFunction_STATE1[132]), .B(
        RoundFunction_T1_n392), .ZN(RoundFunction_TMP3_1[65]) );
  XNOR2_X1 RoundFunction_T1_U229 ( .A(RoundFunction_STATE1[131]), .B(
        RoundFunction_T1_n391), .ZN(RoundFunction_TMP3_1[64]) );
  XNOR2_X1 RoundFunction_T1_U228 ( .A(RoundFunction_STATE1[130]), .B(
        RoundFunction_T1_n390), .ZN(RoundFunction_TMP3_1[71]) );
  XNOR2_X1 RoundFunction_T1_U227 ( .A(RoundFunction_STATE1[12]), .B(
        RoundFunction_T1_n392), .ZN(RoundFunction_TMP3_1[85]) );
  XNOR2_X1 RoundFunction_T1_U226 ( .A(RoundFunction_T1_n346), .B(
        RoundFunction_T1_n345), .ZN(RoundFunction_T1_n392) );
  XNOR2_X1 RoundFunction_T1_U225 ( .A(RoundFunction_STATE1[129]), .B(
        RoundFunction_T1_n400), .ZN(RoundFunction_TMP3_1[70]) );
  XNOR2_X1 RoundFunction_T1_U224 ( .A(RoundFunction_T1_n344), .B(
        RoundFunction_T1_n343), .ZN(RoundFunction_T1_n400) );
  XNOR2_X1 RoundFunction_T1_U223 ( .A(RoundFunction_STATE1[128]), .B(
        RoundFunction_T1_n389), .ZN(RoundFunction_TMP3_1[69]) );
  XNOR2_X1 RoundFunction_T1_U222 ( .A(RoundFunction_T1_n342), .B(
        RoundFunction_T1_n341), .ZN(RoundFunction_T1_n389) );
  XNOR2_X1 RoundFunction_T1_U221 ( .A(RoundFunction_STATE1[127]), .B(
        RoundFunction_T1_n388), .ZN(RoundFunction_TMP3_1[184]) );
  XNOR2_X1 RoundFunction_T1_U220 ( .A(RoundFunction_T1_n340), .B(
        RoundFunction_T1_n339), .ZN(RoundFunction_T1_n388) );
  XNOR2_X1 RoundFunction_T1_U219 ( .A(RoundFunction_STATE1[126]), .B(
        RoundFunction_T1_n387), .ZN(RoundFunction_TMP3_1[191]) );
  XNOR2_X1 RoundFunction_T1_U218 ( .A(RoundFunction_T1_n338), .B(
        RoundFunction_T1_n337), .ZN(RoundFunction_T1_n387) );
  XNOR2_X1 RoundFunction_T1_U217 ( .A(RoundFunction_STATE1[125]), .B(
        RoundFunction_T1_n386), .ZN(RoundFunction_TMP3_1[190]) );
  XNOR2_X1 RoundFunction_T1_U216 ( .A(RoundFunction_T1_n336), .B(
        RoundFunction_T1_n335), .ZN(RoundFunction_T1_n386) );
  XNOR2_X1 RoundFunction_T1_U215 ( .A(RoundFunction_STATE1[124]), .B(
        RoundFunction_T1_n385), .ZN(RoundFunction_TMP3_1[189]) );
  XNOR2_X1 RoundFunction_T1_U214 ( .A(RoundFunction_T1_n334), .B(
        RoundFunction_T1_n359), .ZN(RoundFunction_T1_n385) );
  XOR2_X1 RoundFunction_T1_U213 ( .A(RoundFunction_STATE1[11]), .B(
        RoundFunction_T1_n333), .Z(RoundFunction_T1_n359) );
  XNOR2_X1 RoundFunction_T1_U212 ( .A(RoundFunction_T1_n332), .B(
        RoundFunction_T1_n331), .ZN(RoundFunction_T1_n333) );
  XNOR2_X1 RoundFunction_T1_U211 ( .A(RoundFunction_STATE1[51]), .B(
        RoundFunction_STATE1[91]), .ZN(RoundFunction_T1_n331) );
  XOR2_X1 RoundFunction_T1_U210 ( .A(RoundFunction_STATE1[131]), .B(
        RoundFunction_STATE1[171]), .Z(RoundFunction_T1_n332) );
  XNOR2_X1 RoundFunction_T1_U209 ( .A(RoundFunction_STATE1[123]), .B(
        RoundFunction_T1_n384), .ZN(RoundFunction_TMP3_1[188]) );
  XNOR2_X1 RoundFunction_T1_U208 ( .A(RoundFunction_T1_n330), .B(
        RoundFunction_T1_n357), .ZN(RoundFunction_T1_n384) );
  XOR2_X1 RoundFunction_T1_U207 ( .A(RoundFunction_STATE1[10]), .B(
        RoundFunction_T1_n329), .Z(RoundFunction_T1_n357) );
  XNOR2_X1 RoundFunction_T1_U206 ( .A(RoundFunction_T1_n328), .B(
        RoundFunction_T1_n327), .ZN(RoundFunction_T1_n329) );
  XNOR2_X1 RoundFunction_T1_U205 ( .A(RoundFunction_STATE1[50]), .B(
        RoundFunction_STATE1[90]), .ZN(RoundFunction_T1_n327) );
  XOR2_X1 RoundFunction_T1_U204 ( .A(RoundFunction_STATE1[130]), .B(
        RoundFunction_STATE1[170]), .Z(RoundFunction_T1_n328) );
  XNOR2_X1 RoundFunction_T1_U203 ( .A(RoundFunction_STATE1[122]), .B(
        RoundFunction_T1_n383), .ZN(RoundFunction_TMP3_1[187]) );
  XNOR2_X1 RoundFunction_T1_U202 ( .A(RoundFunction_T1_n326), .B(
        RoundFunction_T1_n355), .ZN(RoundFunction_T1_n383) );
  XOR2_X1 RoundFunction_T1_U201 ( .A(RoundFunction_STATE1[89]), .B(
        RoundFunction_T1_n325), .Z(RoundFunction_T1_n355) );
  XNOR2_X1 RoundFunction_T1_U200 ( .A(RoundFunction_T1_n324), .B(
        RoundFunction_T1_n323), .ZN(RoundFunction_T1_n325) );
  XNOR2_X1 RoundFunction_T1_U199 ( .A(RoundFunction_STATE1[129]), .B(
        RoundFunction_STATE1[49]), .ZN(RoundFunction_T1_n323) );
  XOR2_X1 RoundFunction_T1_U198 ( .A(RoundFunction_STATE1[169]), .B(
        RoundFunction_STATE1[9]), .Z(RoundFunction_T1_n324) );
  XNOR2_X1 RoundFunction_T1_U197 ( .A(RoundFunction_STATE1[121]), .B(
        RoundFunction_T1_n382), .ZN(RoundFunction_TMP3_1[186]) );
  XNOR2_X1 RoundFunction_T1_U196 ( .A(RoundFunction_T1_n322), .B(
        RoundFunction_T1_n353), .ZN(RoundFunction_T1_n382) );
  XOR2_X1 RoundFunction_T1_U195 ( .A(RoundFunction_STATE1[128]), .B(
        RoundFunction_T1_n321), .Z(RoundFunction_T1_n353) );
  XNOR2_X1 RoundFunction_T1_U194 ( .A(RoundFunction_T1_n320), .B(
        RoundFunction_T1_n319), .ZN(RoundFunction_T1_n321) );
  XNOR2_X1 RoundFunction_T1_U193 ( .A(RoundFunction_STATE1[48]), .B(
        RoundFunction_STATE1[8]), .ZN(RoundFunction_T1_n319) );
  XOR2_X1 RoundFunction_T1_U192 ( .A(RoundFunction_STATE1[88]), .B(
        RoundFunction_STATE1[168]), .Z(RoundFunction_T1_n320) );
  XNOR2_X1 RoundFunction_T1_U191 ( .A(RoundFunction_STATE1[120]), .B(
        RoundFunction_T1_n381), .ZN(RoundFunction_TMP3_1[185]) );
  XNOR2_X1 RoundFunction_T1_U190 ( .A(RoundFunction_STATE1[11]), .B(
        RoundFunction_T1_n391), .ZN(RoundFunction_TMP3_1[84]) );
  XNOR2_X1 RoundFunction_T1_U189 ( .A(RoundFunction_T1_n318), .B(
        RoundFunction_T1_n317), .ZN(RoundFunction_T1_n391) );
  XNOR2_X1 RoundFunction_T1_U188 ( .A(RoundFunction_STATE1[119]), .B(
        RoundFunction_T1_n380), .ZN(RoundFunction_TMP3_1[182]) );
  XNOR2_X1 RoundFunction_T1_U187 ( .A(RoundFunction_T1_n354), .B(
        RoundFunction_T1_n349), .ZN(RoundFunction_T1_n380) );
  XOR2_X1 RoundFunction_T1_U186 ( .A(RoundFunction_STATE1[126]), .B(
        RoundFunction_T1_n316), .Z(RoundFunction_T1_n349) );
  XNOR2_X1 RoundFunction_T1_U185 ( .A(RoundFunction_T1_n315), .B(
        RoundFunction_T1_n314), .ZN(RoundFunction_T1_n316) );
  XNOR2_X1 RoundFunction_T1_U184 ( .A(RoundFunction_STATE1[46]), .B(
        RoundFunction_STATE1[86]), .ZN(RoundFunction_T1_n314) );
  XOR2_X1 RoundFunction_T1_U183 ( .A(RoundFunction_STATE1[6]), .B(
        RoundFunction_STATE1[166]), .Z(RoundFunction_T1_n315) );
  XOR2_X1 RoundFunction_T1_U182 ( .A(RoundFunction_STATE1[111]), .B(
        RoundFunction_T1_n313), .Z(RoundFunction_T1_n354) );
  XNOR2_X1 RoundFunction_T1_U181 ( .A(RoundFunction_T1_n312), .B(
        RoundFunction_T1_n311), .ZN(RoundFunction_T1_n313) );
  XNOR2_X1 RoundFunction_T1_U180 ( .A(RoundFunction_STATE1[31]), .B(
        RoundFunction_STATE1[71]), .ZN(RoundFunction_T1_n311) );
  XOR2_X1 RoundFunction_T1_U179 ( .A(RoundFunction_STATE1[151]), .B(
        RoundFunction_STATE1[191]), .Z(RoundFunction_T1_n312) );
  XNOR2_X1 RoundFunction_T1_U178 ( .A(RoundFunction_STATE1[118]), .B(
        RoundFunction_T1_n379), .ZN(RoundFunction_TMP3_1[181]) );
  XNOR2_X1 RoundFunction_T1_U177 ( .A(RoundFunction_T1_n310), .B(
        RoundFunction_T1_n347), .ZN(RoundFunction_T1_n379) );
  XOR2_X1 RoundFunction_T1_U176 ( .A(RoundFunction_STATE1[125]), .B(
        RoundFunction_T1_n309), .Z(RoundFunction_T1_n347) );
  XNOR2_X1 RoundFunction_T1_U175 ( .A(RoundFunction_T1_n308), .B(
        RoundFunction_T1_n307), .ZN(RoundFunction_T1_n309) );
  XNOR2_X1 RoundFunction_T1_U174 ( .A(RoundFunction_STATE1[45]), .B(
        RoundFunction_STATE1[85]), .ZN(RoundFunction_T1_n307) );
  XOR2_X1 RoundFunction_T1_U173 ( .A(RoundFunction_STATE1[5]), .B(
        RoundFunction_STATE1[165]), .Z(RoundFunction_T1_n308) );
  XNOR2_X1 RoundFunction_T1_U172 ( .A(RoundFunction_STATE1[117]), .B(
        RoundFunction_T1_n378), .ZN(RoundFunction_TMP3_1[180]) );
  XNOR2_X1 RoundFunction_T1_U171 ( .A(RoundFunction_T1_n306), .B(
        RoundFunction_T1_n345), .ZN(RoundFunction_T1_n378) );
  XOR2_X1 RoundFunction_T1_U170 ( .A(RoundFunction_STATE1[124]), .B(
        RoundFunction_T1_n305), .Z(RoundFunction_T1_n345) );
  XNOR2_X1 RoundFunction_T1_U169 ( .A(RoundFunction_T1_n304), .B(
        RoundFunction_T1_n303), .ZN(RoundFunction_T1_n305) );
  XNOR2_X1 RoundFunction_T1_U168 ( .A(RoundFunction_STATE1[44]), .B(
        RoundFunction_STATE1[84]), .ZN(RoundFunction_T1_n303) );
  XOR2_X1 RoundFunction_T1_U167 ( .A(RoundFunction_STATE1[4]), .B(
        RoundFunction_STATE1[164]), .Z(RoundFunction_T1_n304) );
  XNOR2_X1 RoundFunction_T1_U166 ( .A(RoundFunction_STATE1[116]), .B(
        RoundFunction_T1_n377), .ZN(RoundFunction_TMP3_1[179]) );
  XNOR2_X1 RoundFunction_T1_U165 ( .A(RoundFunction_T1_n302), .B(
        RoundFunction_T1_n317), .ZN(RoundFunction_T1_n377) );
  XOR2_X1 RoundFunction_T1_U164 ( .A(RoundFunction_STATE1[123]), .B(
        RoundFunction_T1_n301), .Z(RoundFunction_T1_n317) );
  XNOR2_X1 RoundFunction_T1_U163 ( .A(RoundFunction_T1_n300), .B(
        RoundFunction_T1_n299), .ZN(RoundFunction_T1_n301) );
  XNOR2_X1 RoundFunction_T1_U162 ( .A(RoundFunction_STATE1[3]), .B(
        RoundFunction_STATE1[83]), .ZN(RoundFunction_T1_n299) );
  XOR2_X1 RoundFunction_T1_U161 ( .A(RoundFunction_STATE1[43]), .B(
        RoundFunction_STATE1[163]), .Z(RoundFunction_T1_n300) );
  XNOR2_X1 RoundFunction_T1_U160 ( .A(RoundFunction_STATE1[115]), .B(
        RoundFunction_T1_n376), .ZN(RoundFunction_TMP3_1[178]) );
  XNOR2_X1 RoundFunction_T1_U159 ( .A(RoundFunction_T1_n298), .B(
        RoundFunction_T1_n297), .ZN(RoundFunction_T1_n376) );
  XNOR2_X1 RoundFunction_T1_U158 ( .A(RoundFunction_STATE1[114]), .B(
        RoundFunction_T1_n375), .ZN(RoundFunction_TMP3_1[177]) );
  XNOR2_X1 RoundFunction_T1_U157 ( .A(RoundFunction_T1_n343), .B(
        RoundFunction_T1_n360), .ZN(RoundFunction_T1_n375) );
  XOR2_X1 RoundFunction_T1_U156 ( .A(RoundFunction_STATE1[106]), .B(
        RoundFunction_T1_n296), .Z(RoundFunction_T1_n360) );
  XNOR2_X1 RoundFunction_T1_U155 ( .A(RoundFunction_T1_n295), .B(
        RoundFunction_T1_n294), .ZN(RoundFunction_T1_n296) );
  XNOR2_X1 RoundFunction_T1_U154 ( .A(RoundFunction_STATE1[26]), .B(
        RoundFunction_STATE1[66]), .ZN(RoundFunction_T1_n294) );
  XOR2_X1 RoundFunction_T1_U153 ( .A(RoundFunction_STATE1[146]), .B(
        RoundFunction_STATE1[186]), .Z(RoundFunction_T1_n295) );
  XOR2_X1 RoundFunction_T1_U152 ( .A(RoundFunction_STATE1[121]), .B(
        RoundFunction_T1_n293), .Z(RoundFunction_T1_n343) );
  XNOR2_X1 RoundFunction_T1_U151 ( .A(RoundFunction_T1_n292), .B(
        RoundFunction_T1_n291), .ZN(RoundFunction_T1_n293) );
  XNOR2_X1 RoundFunction_T1_U150 ( .A(RoundFunction_STATE1[1]), .B(
        RoundFunction_STATE1[81]), .ZN(RoundFunction_T1_n291) );
  XOR2_X1 RoundFunction_T1_U149 ( .A(RoundFunction_STATE1[41]), .B(
        RoundFunction_STATE1[161]), .Z(RoundFunction_T1_n292) );
  XNOR2_X1 RoundFunction_T1_U148 ( .A(RoundFunction_STATE1[113]), .B(
        RoundFunction_T1_n374), .ZN(RoundFunction_TMP3_1[176]) );
  XNOR2_X1 RoundFunction_T1_U147 ( .A(RoundFunction_T1_n358), .B(
        RoundFunction_T1_n341), .ZN(RoundFunction_T1_n374) );
  XOR2_X1 RoundFunction_T1_U146 ( .A(RoundFunction_STATE1[0]), .B(
        RoundFunction_T1_n290), .Z(RoundFunction_T1_n341) );
  XNOR2_X1 RoundFunction_T1_U145 ( .A(RoundFunction_T1_n289), .B(
        RoundFunction_T1_n288), .ZN(RoundFunction_T1_n290) );
  XNOR2_X1 RoundFunction_T1_U144 ( .A(RoundFunction_STATE1[40]), .B(
        RoundFunction_STATE1[80]), .ZN(RoundFunction_T1_n288) );
  XOR2_X1 RoundFunction_T1_U143 ( .A(RoundFunction_STATE1[120]), .B(
        RoundFunction_STATE1[160]), .Z(RoundFunction_T1_n289) );
  XOR2_X1 RoundFunction_T1_U142 ( .A(RoundFunction_STATE1[105]), .B(
        RoundFunction_T1_n287), .Z(RoundFunction_T1_n358) );
  XNOR2_X1 RoundFunction_T1_U141 ( .A(RoundFunction_T1_n286), .B(
        RoundFunction_T1_n285), .ZN(RoundFunction_T1_n287) );
  XNOR2_X1 RoundFunction_T1_U140 ( .A(RoundFunction_STATE1[25]), .B(
        RoundFunction_STATE1[65]), .ZN(RoundFunction_T1_n285) );
  XOR2_X1 RoundFunction_T1_U139 ( .A(RoundFunction_STATE1[145]), .B(
        RoundFunction_STATE1[185]), .Z(RoundFunction_T1_n286) );
  XNOR2_X1 RoundFunction_T1_U138 ( .A(RoundFunction_STATE1[112]), .B(
        RoundFunction_T1_n373), .ZN(RoundFunction_TMP3_1[183]) );
  XNOR2_X1 RoundFunction_T1_U137 ( .A(RoundFunction_T1_n356), .B(
        RoundFunction_T1_n351), .ZN(RoundFunction_T1_n373) );
  XOR2_X1 RoundFunction_T1_U136 ( .A(RoundFunction_STATE1[127]), .B(
        RoundFunction_T1_n284), .Z(RoundFunction_T1_n351) );
  XNOR2_X1 RoundFunction_T1_U135 ( .A(RoundFunction_T1_n283), .B(
        RoundFunction_T1_n282), .ZN(RoundFunction_T1_n284) );
  XNOR2_X1 RoundFunction_T1_U134 ( .A(RoundFunction_STATE1[47]), .B(
        RoundFunction_STATE1[87]), .ZN(RoundFunction_T1_n282) );
  XOR2_X1 RoundFunction_T1_U133 ( .A(RoundFunction_STATE1[7]), .B(
        RoundFunction_STATE1[167]), .Z(RoundFunction_T1_n283) );
  XOR2_X1 RoundFunction_T1_U132 ( .A(RoundFunction_STATE1[104]), .B(
        RoundFunction_T1_n281), .Z(RoundFunction_T1_n356) );
  XNOR2_X1 RoundFunction_T1_U131 ( .A(RoundFunction_T1_n280), .B(
        RoundFunction_T1_n279), .ZN(RoundFunction_T1_n281) );
  XNOR2_X1 RoundFunction_T1_U130 ( .A(RoundFunction_STATE1[24]), .B(
        RoundFunction_STATE1[64]), .ZN(RoundFunction_T1_n279) );
  XOR2_X1 RoundFunction_T1_U129 ( .A(RoundFunction_STATE1[144]), .B(
        RoundFunction_STATE1[184]), .Z(RoundFunction_T1_n280) );
  XNOR2_X1 RoundFunction_T1_U128 ( .A(RoundFunction_STATE1[111]), .B(
        RoundFunction_T1_n372), .ZN(RoundFunction_TMP3_1[96]) );
  XNOR2_X1 RoundFunction_T1_U127 ( .A(RoundFunction_T1_n342), .B(
        RoundFunction_T1_n337), .ZN(RoundFunction_T1_n372) );
  XOR2_X1 RoundFunction_T1_U126 ( .A(RoundFunction_STATE1[118]), .B(
        RoundFunction_T1_n278), .Z(RoundFunction_T1_n337) );
  XNOR2_X1 RoundFunction_T1_U125 ( .A(RoundFunction_T1_n277), .B(
        RoundFunction_T1_n276), .ZN(RoundFunction_T1_n278) );
  XNOR2_X1 RoundFunction_T1_U124 ( .A(RoundFunction_STATE1[198]), .B(
        RoundFunction_STATE1[78]), .ZN(RoundFunction_T1_n276) );
  XOR2_X1 RoundFunction_T1_U123 ( .A(RoundFunction_STATE1[38]), .B(
        RoundFunction_STATE1[158]), .Z(RoundFunction_T1_n277) );
  XOR2_X1 RoundFunction_T1_U122 ( .A(RoundFunction_STATE1[103]), .B(
        RoundFunction_T1_n275), .Z(RoundFunction_T1_n342) );
  XNOR2_X1 RoundFunction_T1_U121 ( .A(RoundFunction_T1_n274), .B(
        RoundFunction_T1_n273), .ZN(RoundFunction_T1_n275) );
  XNOR2_X1 RoundFunction_T1_U120 ( .A(RoundFunction_STATE1[23]), .B(
        RoundFunction_STATE1[63]), .ZN(RoundFunction_T1_n273) );
  XOR2_X1 RoundFunction_T1_U119 ( .A(RoundFunction_STATE1[143]), .B(
        RoundFunction_STATE1[183]), .Z(RoundFunction_T1_n274) );
  XNOR2_X1 RoundFunction_T1_U118 ( .A(RoundFunction_STATE1[110]), .B(
        RoundFunction_T1_n371), .ZN(RoundFunction_TMP3_1[103]) );
  XNOR2_X1 RoundFunction_T1_U117 ( .A(RoundFunction_T1_n352), .B(
        RoundFunction_T1_n335), .ZN(RoundFunction_T1_n371) );
  XOR2_X1 RoundFunction_T1_U116 ( .A(RoundFunction_STATE1[117]), .B(
        RoundFunction_T1_n272), .Z(RoundFunction_T1_n335) );
  XNOR2_X1 RoundFunction_T1_U115 ( .A(RoundFunction_T1_n271), .B(
        RoundFunction_T1_n270), .ZN(RoundFunction_T1_n272) );
  XNOR2_X1 RoundFunction_T1_U114 ( .A(RoundFunction_STATE1[197]), .B(
        RoundFunction_STATE1[77]), .ZN(RoundFunction_T1_n270) );
  XOR2_X1 RoundFunction_T1_U113 ( .A(RoundFunction_STATE1[37]), .B(
        RoundFunction_STATE1[157]), .Z(RoundFunction_T1_n271) );
  XOR2_X1 RoundFunction_T1_U112 ( .A(RoundFunction_STATE1[102]), .B(
        RoundFunction_T1_n269), .Z(RoundFunction_T1_n352) );
  XNOR2_X1 RoundFunction_T1_U111 ( .A(RoundFunction_T1_n268), .B(
        RoundFunction_T1_n267), .ZN(RoundFunction_T1_n269) );
  XNOR2_X1 RoundFunction_T1_U110 ( .A(RoundFunction_STATE1[22]), .B(
        RoundFunction_STATE1[62]), .ZN(RoundFunction_T1_n267) );
  XOR2_X1 RoundFunction_T1_U109 ( .A(RoundFunction_STATE1[142]), .B(
        RoundFunction_STATE1[182]), .Z(RoundFunction_T1_n268) );
  XNOR2_X1 RoundFunction_T1_U108 ( .A(RoundFunction_STATE1[10]), .B(
        RoundFunction_T1_n390), .ZN(RoundFunction_TMP3_1[83]) );
  XNOR2_X1 RoundFunction_T1_U107 ( .A(RoundFunction_T1_n266), .B(
        RoundFunction_T1_n297), .ZN(RoundFunction_T1_n390) );
  XOR2_X1 RoundFunction_T1_U106 ( .A(RoundFunction_STATE1[122]), .B(
        RoundFunction_T1_n265), .Z(RoundFunction_T1_n297) );
  XNOR2_X1 RoundFunction_T1_U105 ( .A(RoundFunction_T1_n264), .B(
        RoundFunction_T1_n263), .ZN(RoundFunction_T1_n265) );
  XNOR2_X1 RoundFunction_T1_U104 ( .A(RoundFunction_STATE1[2]), .B(
        RoundFunction_STATE1[82]), .ZN(RoundFunction_T1_n263) );
  XOR2_X1 RoundFunction_T1_U103 ( .A(RoundFunction_STATE1[42]), .B(
        RoundFunction_STATE1[162]), .Z(RoundFunction_T1_n264) );
  XNOR2_X1 RoundFunction_T1_U102 ( .A(RoundFunction_STATE1[109]), .B(
        RoundFunction_T1_n370), .ZN(RoundFunction_TMP3_1[102]) );
  XNOR2_X1 RoundFunction_T1_U101 ( .A(RoundFunction_T1_n350), .B(
        RoundFunction_T1_n334), .ZN(RoundFunction_T1_n370) );
  XOR2_X1 RoundFunction_T1_U100 ( .A(RoundFunction_STATE1[116]), .B(
        RoundFunction_T1_n262), .Z(RoundFunction_T1_n334) );
  XNOR2_X1 RoundFunction_T1_U99 ( .A(RoundFunction_T1_n261), .B(
        RoundFunction_T1_n260), .ZN(RoundFunction_T1_n262) );
  XNOR2_X1 RoundFunction_T1_U98 ( .A(RoundFunction_STATE1[196]), .B(
        RoundFunction_STATE1[76]), .ZN(RoundFunction_T1_n260) );
  XOR2_X1 RoundFunction_T1_U97 ( .A(RoundFunction_STATE1[36]), .B(
        RoundFunction_STATE1[156]), .Z(RoundFunction_T1_n261) );
  XOR2_X1 RoundFunction_T1_U96 ( .A(RoundFunction_STATE1[101]), .B(
        RoundFunction_T1_n259), .Z(RoundFunction_T1_n350) );
  XNOR2_X1 RoundFunction_T1_U95 ( .A(RoundFunction_T1_n258), .B(
        RoundFunction_T1_n257), .ZN(RoundFunction_T1_n259) );
  XNOR2_X1 RoundFunction_T1_U94 ( .A(RoundFunction_STATE1[21]), .B(
        RoundFunction_STATE1[61]), .ZN(RoundFunction_T1_n257) );
  XOR2_X1 RoundFunction_T1_U93 ( .A(RoundFunction_STATE1[141]), .B(
        RoundFunction_STATE1[181]), .Z(RoundFunction_T1_n258) );
  XNOR2_X1 RoundFunction_T1_U92 ( .A(RoundFunction_STATE1[108]), .B(
        RoundFunction_T1_n369), .ZN(RoundFunction_TMP3_1[101]) );
  XNOR2_X1 RoundFunction_T1_U91 ( .A(RoundFunction_T1_n348), .B(
        RoundFunction_T1_n330), .ZN(RoundFunction_T1_n369) );
  XOR2_X1 RoundFunction_T1_U90 ( .A(RoundFunction_STATE1[115]), .B(
        RoundFunction_T1_n256), .Z(RoundFunction_T1_n330) );
  XNOR2_X1 RoundFunction_T1_U89 ( .A(RoundFunction_T1_n255), .B(
        RoundFunction_T1_n254), .ZN(RoundFunction_T1_n256) );
  XNOR2_X1 RoundFunction_T1_U88 ( .A(RoundFunction_STATE1[195]), .B(
        RoundFunction_STATE1[75]), .ZN(RoundFunction_T1_n254) );
  XOR2_X1 RoundFunction_T1_U87 ( .A(RoundFunction_STATE1[35]), .B(
        RoundFunction_STATE1[155]), .Z(RoundFunction_T1_n255) );
  XOR2_X1 RoundFunction_T1_U86 ( .A(RoundFunction_STATE1[100]), .B(
        RoundFunction_T1_n253), .Z(RoundFunction_T1_n348) );
  XNOR2_X1 RoundFunction_T1_U85 ( .A(RoundFunction_T1_n252), .B(
        RoundFunction_T1_n251), .ZN(RoundFunction_T1_n253) );
  XNOR2_X1 RoundFunction_T1_U84 ( .A(RoundFunction_STATE1[20]), .B(
        RoundFunction_STATE1[60]), .ZN(RoundFunction_T1_n251) );
  XOR2_X1 RoundFunction_T1_U83 ( .A(RoundFunction_STATE1[140]), .B(
        RoundFunction_STATE1[180]), .Z(RoundFunction_T1_n252) );
  XNOR2_X1 RoundFunction_T1_U82 ( .A(RoundFunction_STATE1[107]), .B(
        RoundFunction_T1_n368), .ZN(RoundFunction_TMP3_1[100]) );
  XNOR2_X1 RoundFunction_T1_U81 ( .A(RoundFunction_T1_n346), .B(
        RoundFunction_T1_n326), .ZN(RoundFunction_T1_n368) );
  XOR2_X1 RoundFunction_T1_U80 ( .A(RoundFunction_STATE1[114]), .B(
        RoundFunction_T1_n250), .Z(RoundFunction_T1_n326) );
  XNOR2_X1 RoundFunction_T1_U79 ( .A(RoundFunction_T1_n249), .B(
        RoundFunction_T1_n248), .ZN(RoundFunction_T1_n250) );
  XNOR2_X1 RoundFunction_T1_U78 ( .A(RoundFunction_STATE1[194]), .B(
        RoundFunction_STATE1[74]), .ZN(RoundFunction_T1_n248) );
  XOR2_X1 RoundFunction_T1_U77 ( .A(RoundFunction_STATE1[34]), .B(
        RoundFunction_STATE1[154]), .Z(RoundFunction_T1_n249) );
  XOR2_X1 RoundFunction_T1_U76 ( .A(RoundFunction_STATE1[59]), .B(
        RoundFunction_T1_n247), .Z(RoundFunction_T1_n346) );
  XNOR2_X1 RoundFunction_T1_U75 ( .A(RoundFunction_T1_n246), .B(
        RoundFunction_T1_n245), .ZN(RoundFunction_T1_n247) );
  XNOR2_X1 RoundFunction_T1_U74 ( .A(RoundFunction_STATE1[139]), .B(
        RoundFunction_STATE1[19]), .ZN(RoundFunction_T1_n245) );
  XOR2_X1 RoundFunction_T1_U73 ( .A(RoundFunction_STATE1[179]), .B(
        RoundFunction_STATE1[99]), .Z(RoundFunction_T1_n246) );
  XNOR2_X1 RoundFunction_T1_U72 ( .A(RoundFunction_STATE1[106]), .B(
        RoundFunction_T1_n367), .ZN(RoundFunction_TMP3_1[99]) );
  XNOR2_X1 RoundFunction_T1_U71 ( .A(RoundFunction_T1_n318), .B(
        RoundFunction_T1_n322), .ZN(RoundFunction_T1_n367) );
  XOR2_X1 RoundFunction_T1_U70 ( .A(RoundFunction_STATE1[113]), .B(
        RoundFunction_T1_n244), .Z(RoundFunction_T1_n322) );
  XNOR2_X1 RoundFunction_T1_U69 ( .A(RoundFunction_T1_n243), .B(
        RoundFunction_T1_n242), .ZN(RoundFunction_T1_n244) );
  XNOR2_X1 RoundFunction_T1_U68 ( .A(RoundFunction_STATE1[193]), .B(
        RoundFunction_STATE1[73]), .ZN(RoundFunction_T1_n242) );
  XOR2_X1 RoundFunction_T1_U67 ( .A(RoundFunction_STATE1[33]), .B(
        RoundFunction_STATE1[153]), .Z(RoundFunction_T1_n243) );
  XOR2_X1 RoundFunction_T1_U66 ( .A(RoundFunction_STATE1[58]), .B(
        RoundFunction_T1_n241), .Z(RoundFunction_T1_n318) );
  XNOR2_X1 RoundFunction_T1_U65 ( .A(RoundFunction_T1_n240), .B(
        RoundFunction_T1_n239), .ZN(RoundFunction_T1_n241) );
  XNOR2_X1 RoundFunction_T1_U64 ( .A(RoundFunction_STATE1[138]), .B(
        RoundFunction_STATE1[18]), .ZN(RoundFunction_T1_n239) );
  XOR2_X1 RoundFunction_T1_U63 ( .A(RoundFunction_STATE1[178]), .B(
        RoundFunction_STATE1[98]), .Z(RoundFunction_T1_n240) );
  XNOR2_X1 RoundFunction_T1_U62 ( .A(RoundFunction_STATE1[105]), .B(
        RoundFunction_T1_n366), .ZN(RoundFunction_TMP3_1[98]) );
  XNOR2_X1 RoundFunction_T1_U61 ( .A(RoundFunction_T1_n238), .B(
        RoundFunction_T1_n266), .ZN(RoundFunction_T1_n366) );
  XOR2_X1 RoundFunction_T1_U60 ( .A(RoundFunction_STATE1[57]), .B(
        RoundFunction_T1_n237), .Z(RoundFunction_T1_n266) );
  XNOR2_X1 RoundFunction_T1_U59 ( .A(RoundFunction_T1_n236), .B(
        RoundFunction_T1_n235), .ZN(RoundFunction_T1_n237) );
  XNOR2_X1 RoundFunction_T1_U58 ( .A(RoundFunction_STATE1[137]), .B(
        RoundFunction_STATE1[17]), .ZN(RoundFunction_T1_n235) );
  XOR2_X1 RoundFunction_T1_U57 ( .A(RoundFunction_STATE1[177]), .B(
        RoundFunction_STATE1[97]), .Z(RoundFunction_T1_n236) );
  XNOR2_X1 RoundFunction_T1_U56 ( .A(RoundFunction_STATE1[104]), .B(
        RoundFunction_T1_n365), .ZN(RoundFunction_TMP3_1[97]) );
  XNOR2_X1 RoundFunction_T1_U55 ( .A(RoundFunction_T1_n344), .B(
        RoundFunction_T1_n339), .ZN(RoundFunction_T1_n365) );
  XOR2_X1 RoundFunction_T1_U54 ( .A(RoundFunction_STATE1[119]), .B(
        RoundFunction_T1_n234), .Z(RoundFunction_T1_n339) );
  XNOR2_X1 RoundFunction_T1_U53 ( .A(RoundFunction_T1_n233), .B(
        RoundFunction_T1_n232), .ZN(RoundFunction_T1_n234) );
  XNOR2_X1 RoundFunction_T1_U52 ( .A(RoundFunction_STATE1[199]), .B(
        RoundFunction_STATE1[79]), .ZN(RoundFunction_T1_n232) );
  XOR2_X1 RoundFunction_T1_U51 ( .A(RoundFunction_STATE1[39]), .B(
        RoundFunction_STATE1[159]), .Z(RoundFunction_T1_n233) );
  XOR2_X1 RoundFunction_T1_U50 ( .A(RoundFunction_STATE1[136]), .B(
        RoundFunction_T1_n231), .Z(RoundFunction_T1_n344) );
  XNOR2_X1 RoundFunction_T1_U49 ( .A(RoundFunction_T1_n230), .B(
        RoundFunction_T1_n229), .ZN(RoundFunction_T1_n231) );
  XNOR2_X1 RoundFunction_T1_U48 ( .A(RoundFunction_STATE1[176]), .B(
        RoundFunction_STATE1[96]), .ZN(RoundFunction_T1_n229) );
  XOR2_X1 RoundFunction_T1_U47 ( .A(RoundFunction_STATE1[56]), .B(
        RoundFunction_STATE1[16]), .Z(RoundFunction_T1_n230) );
  XNOR2_X1 RoundFunction_T1_U46 ( .A(RoundFunction_STATE1[103]), .B(
        RoundFunction_T1_n364), .ZN(RoundFunction_TMP3_1[18]) );
  XNOR2_X1 RoundFunction_T1_U45 ( .A(RoundFunction_T1_n228), .B(
        RoundFunction_T1_n310), .ZN(RoundFunction_T1_n364) );
  XOR2_X1 RoundFunction_T1_U44 ( .A(RoundFunction_STATE1[110]), .B(
        RoundFunction_T1_n227), .Z(RoundFunction_T1_n310) );
  XNOR2_X1 RoundFunction_T1_U43 ( .A(RoundFunction_T1_n226), .B(
        RoundFunction_T1_n225), .ZN(RoundFunction_T1_n227) );
  XNOR2_X1 RoundFunction_T1_U42 ( .A(RoundFunction_STATE1[190]), .B(
        RoundFunction_STATE1[70]), .ZN(RoundFunction_T1_n225) );
  XOR2_X1 RoundFunction_T1_U41 ( .A(RoundFunction_STATE1[30]), .B(
        RoundFunction_STATE1[150]), .Z(RoundFunction_T1_n226) );
  XNOR2_X1 RoundFunction_T1_U40 ( .A(RoundFunction_STATE1[102]), .B(
        RoundFunction_T1_n363), .ZN(RoundFunction_TMP3_1[17]) );
  XNOR2_X1 RoundFunction_T1_U39 ( .A(RoundFunction_T1_n340), .B(
        RoundFunction_T1_n306), .ZN(RoundFunction_T1_n363) );
  XOR2_X1 RoundFunction_T1_U38 ( .A(RoundFunction_STATE1[109]), .B(
        RoundFunction_T1_n224), .Z(RoundFunction_T1_n306) );
  XNOR2_X1 RoundFunction_T1_U37 ( .A(RoundFunction_T1_n223), .B(
        RoundFunction_T1_n222), .ZN(RoundFunction_T1_n224) );
  XNOR2_X1 RoundFunction_T1_U36 ( .A(RoundFunction_STATE1[189]), .B(
        RoundFunction_STATE1[69]), .ZN(RoundFunction_T1_n222) );
  XOR2_X1 RoundFunction_T1_U35 ( .A(RoundFunction_STATE1[29]), .B(
        RoundFunction_STATE1[149]), .Z(RoundFunction_T1_n223) );
  XOR2_X1 RoundFunction_T1_U34 ( .A(RoundFunction_STATE1[54]), .B(
        RoundFunction_T1_n221), .Z(RoundFunction_T1_n340) );
  XNOR2_X1 RoundFunction_T1_U33 ( .A(RoundFunction_T1_n220), .B(
        RoundFunction_T1_n219), .ZN(RoundFunction_T1_n221) );
  XNOR2_X1 RoundFunction_T1_U32 ( .A(RoundFunction_STATE1[134]), .B(
        RoundFunction_STATE1[174]), .ZN(RoundFunction_T1_n219) );
  XOR2_X1 RoundFunction_T1_U31 ( .A(RoundFunction_STATE1[14]), .B(
        RoundFunction_STATE1[94]), .Z(RoundFunction_T1_n220) );
  XNOR2_X1 RoundFunction_T1_U30 ( .A(RoundFunction_STATE1[101]), .B(
        RoundFunction_T1_n362), .ZN(RoundFunction_TMP3_1[16]) );
  XNOR2_X1 RoundFunction_T1_U29 ( .A(RoundFunction_T1_n338), .B(
        RoundFunction_T1_n302), .ZN(RoundFunction_T1_n362) );
  XOR2_X1 RoundFunction_T1_U28 ( .A(RoundFunction_STATE1[108]), .B(
        RoundFunction_T1_n218), .Z(RoundFunction_T1_n302) );
  XNOR2_X1 RoundFunction_T1_U27 ( .A(RoundFunction_T1_n217), .B(
        RoundFunction_T1_n216), .ZN(RoundFunction_T1_n218) );
  XNOR2_X1 RoundFunction_T1_U26 ( .A(RoundFunction_STATE1[188]), .B(
        RoundFunction_STATE1[68]), .ZN(RoundFunction_T1_n216) );
  XOR2_X1 RoundFunction_T1_U25 ( .A(RoundFunction_STATE1[28]), .B(
        RoundFunction_STATE1[148]), .Z(RoundFunction_T1_n217) );
  XOR2_X1 RoundFunction_T1_U24 ( .A(RoundFunction_STATE1[53]), .B(
        RoundFunction_T1_n215), .Z(RoundFunction_T1_n338) );
  XNOR2_X1 RoundFunction_T1_U23 ( .A(RoundFunction_T1_n214), .B(
        RoundFunction_T1_n213), .ZN(RoundFunction_T1_n215) );
  XNOR2_X1 RoundFunction_T1_U22 ( .A(RoundFunction_STATE1[133]), .B(
        RoundFunction_STATE1[173]), .ZN(RoundFunction_T1_n213) );
  XOR2_X1 RoundFunction_T1_U21 ( .A(RoundFunction_STATE1[13]), .B(
        RoundFunction_STATE1[93]), .Z(RoundFunction_T1_n214) );
  XNOR2_X1 RoundFunction_T1_U20 ( .A(RoundFunction_STATE1[100]), .B(
        RoundFunction_T1_n361), .ZN(RoundFunction_TMP3_1[23]) );
  XNOR2_X1 RoundFunction_T1_U19 ( .A(RoundFunction_T1_n336), .B(
        RoundFunction_T1_n298), .ZN(RoundFunction_T1_n361) );
  XOR2_X1 RoundFunction_T1_U18 ( .A(RoundFunction_STATE1[107]), .B(
        RoundFunction_T1_n212), .Z(RoundFunction_T1_n298) );
  XNOR2_X1 RoundFunction_T1_U17 ( .A(RoundFunction_T1_n211), .B(
        RoundFunction_T1_n210), .ZN(RoundFunction_T1_n212) );
  XNOR2_X1 RoundFunction_T1_U16 ( .A(RoundFunction_STATE1[187]), .B(
        RoundFunction_STATE1[67]), .ZN(RoundFunction_T1_n210) );
  XOR2_X1 RoundFunction_T1_U15 ( .A(RoundFunction_STATE1[27]), .B(
        RoundFunction_STATE1[147]), .Z(RoundFunction_T1_n211) );
  XOR2_X1 RoundFunction_T1_U14 ( .A(RoundFunction_STATE1[52]), .B(
        RoundFunction_T1_n209), .Z(RoundFunction_T1_n336) );
  XNOR2_X1 RoundFunction_T1_U13 ( .A(RoundFunction_T1_n208), .B(
        RoundFunction_T1_n207), .ZN(RoundFunction_T1_n209) );
  XNOR2_X1 RoundFunction_T1_U12 ( .A(RoundFunction_STATE1[12]), .B(
        RoundFunction_STATE1[172]), .ZN(RoundFunction_T1_n207) );
  XOR2_X1 RoundFunction_T1_U11 ( .A(RoundFunction_STATE1[132]), .B(
        RoundFunction_STATE1[92]), .Z(RoundFunction_T1_n208) );
  XNOR2_X1 RoundFunction_T1_U10 ( .A(RoundFunction_STATE1[0]), .B(
        RoundFunction_T1_n381), .ZN(RoundFunction_TMP3_1[0]) );
  XNOR2_X1 RoundFunction_T1_U9 ( .A(RoundFunction_T1_n238), .B(
        RoundFunction_T1_n228), .ZN(RoundFunction_T1_n381) );
  XOR2_X1 RoundFunction_T1_U8 ( .A(RoundFunction_STATE1[55]), .B(
        RoundFunction_T1_n206), .Z(RoundFunction_T1_n228) );
  XNOR2_X1 RoundFunction_T1_U7 ( .A(RoundFunction_T1_n205), .B(
        RoundFunction_T1_n204), .ZN(RoundFunction_T1_n206) );
  XNOR2_X1 RoundFunction_T1_U6 ( .A(RoundFunction_STATE1[135]), .B(
        RoundFunction_STATE1[175]), .ZN(RoundFunction_T1_n204) );
  XOR2_X1 RoundFunction_T1_U5 ( .A(RoundFunction_STATE1[15]), .B(
        RoundFunction_STATE1[95]), .Z(RoundFunction_T1_n205) );
  XOR2_X1 RoundFunction_T1_U4 ( .A(RoundFunction_STATE1[112]), .B(
        RoundFunction_T1_n203), .Z(RoundFunction_T1_n238) );
  XNOR2_X1 RoundFunction_T1_U3 ( .A(RoundFunction_T1_n202), .B(
        RoundFunction_T1_n201), .ZN(RoundFunction_T1_n203) );
  XNOR2_X1 RoundFunction_T1_U2 ( .A(RoundFunction_STATE1[192]), .B(
        RoundFunction_STATE1[72]), .ZN(RoundFunction_T1_n201) );
  XOR2_X1 RoundFunction_T1_U1 ( .A(RoundFunction_STATE1[32]), .B(
        RoundFunction_STATE1[152]), .Z(RoundFunction_T1_n202) );
  XOR2_X1 RoundFunction_I1_U8 ( .A(CONST[7]), .B(RoundFunction_TMP4_1[7]), .Z(
        RESULT1[199]) );
  XOR2_X1 RoundFunction_I1_U7 ( .A(1'b0), .B(RoundFunction_TMP4_1[6]), .Z(
        RESULT1[198]) );
  XOR2_X1 RoundFunction_I1_U6 ( .A(1'b0), .B(RoundFunction_TMP4_1[5]), .Z(
        RESULT1[197]) );
  XOR2_X1 RoundFunction_I1_U5 ( .A(1'b0), .B(RoundFunction_TMP4_1[4]), .Z(
        RESULT1[196]) );
  XOR2_X1 RoundFunction_I1_U4 ( .A(CONST[3]), .B(RoundFunction_TMP4_1[3]), .Z(
        RESULT1[195]) );
  XOR2_X1 RoundFunction_I1_U3 ( .A(1'b0), .B(RoundFunction_TMP4_1[2]), .Z(
        RESULT1[194]) );
  XOR2_X1 RoundFunction_I1_U2 ( .A(CONST[1]), .B(RoundFunction_TMP4_1[1]), .Z(
        RESULT1[193]) );
  XOR2_X1 RoundFunction_I1_U1 ( .A(CONST[0]), .B(RoundFunction_TMP4_1[0]), .Z(
        RESULT1[192]) );
  XNOR2_X1 RoundFunction_T2_U400 ( .A(RoundFunction_STATE2[9]), .B(
        RoundFunction_T2_n400), .ZN(RoundFunction_TMP3_2[82]) );
  XNOR2_X1 RoundFunction_T2_U399 ( .A(RoundFunction_STATE2[99]), .B(
        RoundFunction_T2_n399), .ZN(RoundFunction_TMP3_2[22]) );
  XNOR2_X1 RoundFunction_T2_U398 ( .A(RoundFunction_STATE2[98]), .B(
        RoundFunction_T2_n398), .ZN(RoundFunction_TMP3_2[21]) );
  XNOR2_X1 RoundFunction_T2_U397 ( .A(RoundFunction_STATE2[97]), .B(
        RoundFunction_T2_n397), .ZN(RoundFunction_TMP3_2[20]) );
  XNOR2_X1 RoundFunction_T2_U396 ( .A(RoundFunction_STATE2[96]), .B(
        RoundFunction_T2_n396), .ZN(RoundFunction_TMP3_2[19]) );
  XNOR2_X1 RoundFunction_T2_U395 ( .A(RoundFunction_STATE2[95]), .B(
        RoundFunction_T2_n395), .ZN(RoundFunction_TMP3_2[137]) );
  XNOR2_X1 RoundFunction_T2_U394 ( .A(RoundFunction_STATE2[94]), .B(
        RoundFunction_T2_n394), .ZN(RoundFunction_TMP3_2[136]) );
  XNOR2_X1 RoundFunction_T2_U393 ( .A(RoundFunction_STATE2[93]), .B(
        RoundFunction_T2_n393), .ZN(RoundFunction_TMP3_2[143]) );
  XNOR2_X1 RoundFunction_T2_U392 ( .A(RoundFunction_STATE2[92]), .B(
        RoundFunction_T2_n392), .ZN(RoundFunction_TMP3_2[142]) );
  XNOR2_X1 RoundFunction_T2_U391 ( .A(RoundFunction_STATE2[91]), .B(
        RoundFunction_T2_n391), .ZN(RoundFunction_TMP3_2[141]) );
  XNOR2_X1 RoundFunction_T2_U390 ( .A(RoundFunction_STATE2[90]), .B(
        RoundFunction_T2_n390), .ZN(RoundFunction_TMP3_2[140]) );
  XNOR2_X1 RoundFunction_T2_U389 ( .A(RoundFunction_STATE2[8]), .B(
        RoundFunction_T2_n389), .ZN(RoundFunction_TMP3_2[81]) );
  XNOR2_X1 RoundFunction_T2_U388 ( .A(RoundFunction_STATE2[89]), .B(
        RoundFunction_T2_n400), .ZN(RoundFunction_TMP3_2[139]) );
  XNOR2_X1 RoundFunction_T2_U387 ( .A(RoundFunction_STATE2[88]), .B(
        RoundFunction_T2_n389), .ZN(RoundFunction_TMP3_2[138]) );
  XNOR2_X1 RoundFunction_T2_U386 ( .A(RoundFunction_STATE2[87]), .B(
        RoundFunction_T2_n388), .ZN(RoundFunction_TMP3_2[58]) );
  XNOR2_X1 RoundFunction_T2_U385 ( .A(RoundFunction_STATE2[86]), .B(
        RoundFunction_T2_n387), .ZN(RoundFunction_TMP3_2[57]) );
  XNOR2_X1 RoundFunction_T2_U384 ( .A(RoundFunction_STATE2[85]), .B(
        RoundFunction_T2_n386), .ZN(RoundFunction_TMP3_2[56]) );
  XNOR2_X1 RoundFunction_T2_U383 ( .A(RoundFunction_STATE2[84]), .B(
        RoundFunction_T2_n385), .ZN(RoundFunction_TMP3_2[63]) );
  XNOR2_X1 RoundFunction_T2_U382 ( .A(RoundFunction_STATE2[83]), .B(
        RoundFunction_T2_n384), .ZN(RoundFunction_TMP3_2[62]) );
  XNOR2_X1 RoundFunction_T2_U381 ( .A(RoundFunction_STATE2[82]), .B(
        RoundFunction_T2_n383), .ZN(RoundFunction_TMP3_2[61]) );
  XNOR2_X1 RoundFunction_T2_U380 ( .A(RoundFunction_STATE2[81]), .B(
        RoundFunction_T2_n382), .ZN(RoundFunction_TMP3_2[60]) );
  XNOR2_X1 RoundFunction_T2_U379 ( .A(RoundFunction_STATE2[80]), .B(
        RoundFunction_T2_n381), .ZN(RoundFunction_TMP3_2[59]) );
  XNOR2_X1 RoundFunction_T2_U378 ( .A(RoundFunction_STATE2[7]), .B(
        RoundFunction_T2_n388), .ZN(RoundFunction_TMP3_2[7]) );
  XNOR2_X1 RoundFunction_T2_U377 ( .A(RoundFunction_STATE2[79]), .B(
        RoundFunction_T2_n380), .ZN(RoundFunction_TMP3_2[51]) );
  XNOR2_X1 RoundFunction_T2_U376 ( .A(RoundFunction_STATE2[78]), .B(
        RoundFunction_T2_n379), .ZN(RoundFunction_TMP3_2[50]) );
  XNOR2_X1 RoundFunction_T2_U375 ( .A(RoundFunction_STATE2[77]), .B(
        RoundFunction_T2_n378), .ZN(RoundFunction_TMP3_2[49]) );
  XNOR2_X1 RoundFunction_T2_U374 ( .A(RoundFunction_STATE2[76]), .B(
        RoundFunction_T2_n377), .ZN(RoundFunction_TMP3_2[48]) );
  XNOR2_X1 RoundFunction_T2_U373 ( .A(RoundFunction_STATE2[75]), .B(
        RoundFunction_T2_n376), .ZN(RoundFunction_TMP3_2[55]) );
  XNOR2_X1 RoundFunction_T2_U372 ( .A(RoundFunction_STATE2[74]), .B(
        RoundFunction_T2_n375), .ZN(RoundFunction_TMP3_2[54]) );
  XNOR2_X1 RoundFunction_T2_U371 ( .A(RoundFunction_STATE2[73]), .B(
        RoundFunction_T2_n374), .ZN(RoundFunction_TMP3_2[53]) );
  XNOR2_X1 RoundFunction_T2_U370 ( .A(RoundFunction_STATE2[72]), .B(
        RoundFunction_T2_n373), .ZN(RoundFunction_TMP3_2[52]) );
  XNOR2_X1 RoundFunction_T2_U369 ( .A(RoundFunction_STATE2[71]), .B(
        RoundFunction_T2_n372), .ZN(RoundFunction_TMP3_2[174]) );
  XNOR2_X1 RoundFunction_T2_U368 ( .A(RoundFunction_STATE2[70]), .B(
        RoundFunction_T2_n371), .ZN(RoundFunction_TMP3_2[173]) );
  XNOR2_X1 RoundFunction_T2_U367 ( .A(RoundFunction_STATE2[6]), .B(
        RoundFunction_T2_n387), .ZN(RoundFunction_TMP3_2[6]) );
  XNOR2_X1 RoundFunction_T2_U366 ( .A(RoundFunction_STATE2[69]), .B(
        RoundFunction_T2_n370), .ZN(RoundFunction_TMP3_2[172]) );
  XNOR2_X1 RoundFunction_T2_U365 ( .A(RoundFunction_STATE2[68]), .B(
        RoundFunction_T2_n369), .ZN(RoundFunction_TMP3_2[171]) );
  XNOR2_X1 RoundFunction_T2_U364 ( .A(RoundFunction_STATE2[67]), .B(
        RoundFunction_T2_n368), .ZN(RoundFunction_TMP3_2[170]) );
  XNOR2_X1 RoundFunction_T2_U363 ( .A(RoundFunction_STATE2[66]), .B(
        RoundFunction_T2_n367), .ZN(RoundFunction_TMP3_2[169]) );
  XNOR2_X1 RoundFunction_T2_U362 ( .A(RoundFunction_STATE2[65]), .B(
        RoundFunction_T2_n366), .ZN(RoundFunction_TMP3_2[168]) );
  XNOR2_X1 RoundFunction_T2_U361 ( .A(RoundFunction_STATE2[64]), .B(
        RoundFunction_T2_n365), .ZN(RoundFunction_TMP3_2[175]) );
  XNOR2_X1 RoundFunction_T2_U360 ( .A(RoundFunction_STATE2[63]), .B(
        RoundFunction_T2_n364), .ZN(RoundFunction_TMP3_2[93]) );
  XNOR2_X1 RoundFunction_T2_U359 ( .A(RoundFunction_STATE2[62]), .B(
        RoundFunction_T2_n363), .ZN(RoundFunction_TMP3_2[92]) );
  XNOR2_X1 RoundFunction_T2_U358 ( .A(RoundFunction_STATE2[61]), .B(
        RoundFunction_T2_n362), .ZN(RoundFunction_TMP3_2[91]) );
  XNOR2_X1 RoundFunction_T2_U357 ( .A(RoundFunction_STATE2[60]), .B(
        RoundFunction_T2_n361), .ZN(RoundFunction_TMP3_2[90]) );
  XNOR2_X1 RoundFunction_T2_U356 ( .A(RoundFunction_STATE2[5]), .B(
        RoundFunction_T2_n386), .ZN(RoundFunction_TMP3_2[5]) );
  XNOR2_X1 RoundFunction_T2_U355 ( .A(RoundFunction_STATE2[59]), .B(
        RoundFunction_T2_n399), .ZN(RoundFunction_TMP3_2[89]) );
  XNOR2_X1 RoundFunction_T2_U354 ( .A(RoundFunction_STATE2[58]), .B(
        RoundFunction_T2_n398), .ZN(RoundFunction_TMP3_2[88]) );
  XNOR2_X1 RoundFunction_T2_U353 ( .A(RoundFunction_STATE2[57]), .B(
        RoundFunction_T2_n397), .ZN(RoundFunction_TMP3_2[95]) );
  XNOR2_X1 RoundFunction_T2_U352 ( .A(RoundFunction_STATE2[56]), .B(
        RoundFunction_T2_n396), .ZN(RoundFunction_TMP3_2[94]) );
  XNOR2_X1 RoundFunction_T2_U351 ( .A(RoundFunction_STATE2[55]), .B(
        RoundFunction_T2_n395), .ZN(RoundFunction_TMP3_2[11]) );
  XNOR2_X1 RoundFunction_T2_U350 ( .A(RoundFunction_STATE2[54]), .B(
        RoundFunction_T2_n394), .ZN(RoundFunction_TMP3_2[10]) );
  XNOR2_X1 RoundFunction_T2_U349 ( .A(RoundFunction_STATE2[53]), .B(
        RoundFunction_T2_n393), .ZN(RoundFunction_TMP3_2[9]) );
  XNOR2_X1 RoundFunction_T2_U348 ( .A(RoundFunction_STATE2[52]), .B(
        RoundFunction_T2_n392), .ZN(RoundFunction_TMP3_2[8]) );
  XNOR2_X1 RoundFunction_T2_U347 ( .A(RoundFunction_STATE2[51]), .B(
        RoundFunction_T2_n391), .ZN(RoundFunction_TMP3_2[15]) );
  XNOR2_X1 RoundFunction_T2_U346 ( .A(RoundFunction_STATE2[50]), .B(
        RoundFunction_T2_n390), .ZN(RoundFunction_TMP3_2[14]) );
  XNOR2_X1 RoundFunction_T2_U345 ( .A(RoundFunction_STATE2[4]), .B(
        RoundFunction_T2_n385), .ZN(RoundFunction_TMP3_2[4]) );
  XNOR2_X1 RoundFunction_T2_U344 ( .A(RoundFunction_STATE2[49]), .B(
        RoundFunction_T2_n400), .ZN(RoundFunction_TMP3_2[13]) );
  XNOR2_X1 RoundFunction_T2_U343 ( .A(RoundFunction_STATE2[48]), .B(
        RoundFunction_T2_n389), .ZN(RoundFunction_TMP3_2[12]) );
  XNOR2_X1 RoundFunction_T2_U342 ( .A(RoundFunction_STATE2[47]), .B(
        RoundFunction_T2_n388), .ZN(RoundFunction_TMP3_2[131]) );
  XNOR2_X1 RoundFunction_T2_U341 ( .A(RoundFunction_STATE2[46]), .B(
        RoundFunction_T2_n387), .ZN(RoundFunction_TMP3_2[130]) );
  XNOR2_X1 RoundFunction_T2_U340 ( .A(RoundFunction_STATE2[45]), .B(
        RoundFunction_T2_n386), .ZN(RoundFunction_TMP3_2[129]) );
  XNOR2_X1 RoundFunction_T2_U339 ( .A(RoundFunction_STATE2[44]), .B(
        RoundFunction_T2_n385), .ZN(RoundFunction_TMP3_2[128]) );
  XNOR2_X1 RoundFunction_T2_U338 ( .A(RoundFunction_STATE2[43]), .B(
        RoundFunction_T2_n384), .ZN(RoundFunction_TMP3_2[135]) );
  XNOR2_X1 RoundFunction_T2_U337 ( .A(RoundFunction_STATE2[42]), .B(
        RoundFunction_T2_n383), .ZN(RoundFunction_TMP3_2[134]) );
  XNOR2_X1 RoundFunction_T2_U336 ( .A(RoundFunction_STATE2[41]), .B(
        RoundFunction_T2_n382), .ZN(RoundFunction_TMP3_2[133]) );
  XNOR2_X1 RoundFunction_T2_U335 ( .A(RoundFunction_STATE2[40]), .B(
        RoundFunction_T2_n381), .ZN(RoundFunction_TMP3_2[132]) );
  XNOR2_X1 RoundFunction_T2_U334 ( .A(RoundFunction_STATE2[3]), .B(
        RoundFunction_T2_n384), .ZN(RoundFunction_TMP3_2[3]) );
  XNOR2_X1 RoundFunction_T2_U333 ( .A(RoundFunction_STATE2[39]), .B(
        RoundFunction_T2_n380), .ZN(RoundFunction_TMP3_2[122]) );
  XNOR2_X1 RoundFunction_T2_U332 ( .A(RoundFunction_STATE2[38]), .B(
        RoundFunction_T2_n379), .ZN(RoundFunction_TMP3_2[121]) );
  XNOR2_X1 RoundFunction_T2_U331 ( .A(RoundFunction_STATE2[37]), .B(
        RoundFunction_T2_n378), .ZN(RoundFunction_TMP3_2[120]) );
  XNOR2_X1 RoundFunction_T2_U330 ( .A(RoundFunction_STATE2[36]), .B(
        RoundFunction_T2_n377), .ZN(RoundFunction_TMP3_2[127]) );
  XNOR2_X1 RoundFunction_T2_U329 ( .A(RoundFunction_STATE2[35]), .B(
        RoundFunction_T2_n376), .ZN(RoundFunction_TMP3_2[126]) );
  XNOR2_X1 RoundFunction_T2_U328 ( .A(RoundFunction_STATE2[34]), .B(
        RoundFunction_T2_n375), .ZN(RoundFunction_TMP3_2[125]) );
  XNOR2_X1 RoundFunction_T2_U327 ( .A(RoundFunction_STATE2[33]), .B(
        RoundFunction_T2_n374), .ZN(RoundFunction_TMP3_2[124]) );
  XNOR2_X1 RoundFunction_T2_U326 ( .A(RoundFunction_STATE2[32]), .B(
        RoundFunction_T2_n373), .ZN(RoundFunction_TMP3_2[123]) );
  XNOR2_X1 RoundFunction_T2_U325 ( .A(RoundFunction_STATE2[31]), .B(
        RoundFunction_T2_n372), .ZN(RoundFunction_TMP3_2[43]) );
  XNOR2_X1 RoundFunction_T2_U324 ( .A(RoundFunction_STATE2[30]), .B(
        RoundFunction_T2_n371), .ZN(RoundFunction_TMP3_2[42]) );
  XNOR2_X1 RoundFunction_T2_U323 ( .A(RoundFunction_STATE2[2]), .B(
        RoundFunction_T2_n383), .ZN(RoundFunction_TMP3_2[2]) );
  XNOR2_X1 RoundFunction_T2_U322 ( .A(RoundFunction_STATE2[29]), .B(
        RoundFunction_T2_n370), .ZN(RoundFunction_TMP3_2[41]) );
  XNOR2_X1 RoundFunction_T2_U321 ( .A(RoundFunction_STATE2[28]), .B(
        RoundFunction_T2_n369), .ZN(RoundFunction_TMP3_2[40]) );
  XNOR2_X1 RoundFunction_T2_U320 ( .A(RoundFunction_STATE2[27]), .B(
        RoundFunction_T2_n368), .ZN(RoundFunction_TMP3_2[47]) );
  XNOR2_X1 RoundFunction_T2_U319 ( .A(RoundFunction_STATE2[26]), .B(
        RoundFunction_T2_n367), .ZN(RoundFunction_TMP3_2[46]) );
  XNOR2_X1 RoundFunction_T2_U318 ( .A(RoundFunction_STATE2[25]), .B(
        RoundFunction_T2_n366), .ZN(RoundFunction_TMP3_2[45]) );
  XNOR2_X1 RoundFunction_T2_U317 ( .A(RoundFunction_STATE2[24]), .B(
        RoundFunction_T2_n365), .ZN(RoundFunction_TMP3_2[44]) );
  XNOR2_X1 RoundFunction_T2_U316 ( .A(RoundFunction_STATE2[23]), .B(
        RoundFunction_T2_n364), .ZN(RoundFunction_TMP3_2[165]) );
  XNOR2_X1 RoundFunction_T2_U315 ( .A(RoundFunction_STATE2[22]), .B(
        RoundFunction_T2_n363), .ZN(RoundFunction_TMP3_2[164]) );
  XNOR2_X1 RoundFunction_T2_U314 ( .A(RoundFunction_STATE2[21]), .B(
        RoundFunction_T2_n362), .ZN(RoundFunction_TMP3_2[163]) );
  XNOR2_X1 RoundFunction_T2_U313 ( .A(RoundFunction_STATE2[20]), .B(
        RoundFunction_T2_n361), .ZN(RoundFunction_TMP3_2[162]) );
  XNOR2_X1 RoundFunction_T2_U312 ( .A(RoundFunction_STATE2[1]), .B(
        RoundFunction_T2_n382), .ZN(RoundFunction_TMP3_2[1]) );
  XNOR2_X1 RoundFunction_T2_U311 ( .A(RoundFunction_STATE2[19]), .B(
        RoundFunction_T2_n399), .ZN(RoundFunction_TMP3_2[161]) );
  XNOR2_X1 RoundFunction_T2_U310 ( .A(RoundFunction_STATE2[199]), .B(
        RoundFunction_T2_n380), .ZN(RoundFunction_TMP3_2[37]) );
  XNOR2_X1 RoundFunction_T2_U309 ( .A(RoundFunction_STATE2[198]), .B(
        RoundFunction_T2_n379), .ZN(RoundFunction_TMP3_2[36]) );
  XNOR2_X1 RoundFunction_T2_U308 ( .A(RoundFunction_STATE2[197]), .B(
        RoundFunction_T2_n378), .ZN(RoundFunction_TMP3_2[35]) );
  XNOR2_X1 RoundFunction_T2_U307 ( .A(RoundFunction_STATE2[196]), .B(
        RoundFunction_T2_n377), .ZN(RoundFunction_TMP3_2[34]) );
  XNOR2_X1 RoundFunction_T2_U306 ( .A(RoundFunction_STATE2[195]), .B(
        RoundFunction_T2_n376), .ZN(RoundFunction_TMP3_2[33]) );
  XNOR2_X1 RoundFunction_T2_U305 ( .A(RoundFunction_STATE2[194]), .B(
        RoundFunction_T2_n375), .ZN(RoundFunction_TMP3_2[32]) );
  XNOR2_X1 RoundFunction_T2_U304 ( .A(RoundFunction_STATE2[193]), .B(
        RoundFunction_T2_n374), .ZN(RoundFunction_TMP3_2[39]) );
  XNOR2_X1 RoundFunction_T2_U303 ( .A(RoundFunction_STATE2[192]), .B(
        RoundFunction_T2_n373), .ZN(RoundFunction_TMP3_2[38]) );
  XNOR2_X1 RoundFunction_T2_U302 ( .A(RoundFunction_STATE2[191]), .B(
        RoundFunction_T2_n372), .ZN(RoundFunction_TMP3_2[159]) );
  XNOR2_X1 RoundFunction_T2_U301 ( .A(RoundFunction_STATE2[190]), .B(
        RoundFunction_T2_n371), .ZN(RoundFunction_TMP3_2[158]) );
  XNOR2_X1 RoundFunction_T2_U300 ( .A(RoundFunction_STATE2[18]), .B(
        RoundFunction_T2_n398), .ZN(RoundFunction_TMP3_2[160]) );
  XNOR2_X1 RoundFunction_T2_U299 ( .A(RoundFunction_STATE2[189]), .B(
        RoundFunction_T2_n370), .ZN(RoundFunction_TMP3_2[157]) );
  XNOR2_X1 RoundFunction_T2_U298 ( .A(RoundFunction_STATE2[188]), .B(
        RoundFunction_T2_n369), .ZN(RoundFunction_TMP3_2[156]) );
  XNOR2_X1 RoundFunction_T2_U297 ( .A(RoundFunction_STATE2[187]), .B(
        RoundFunction_T2_n368), .ZN(RoundFunction_TMP3_2[155]) );
  XNOR2_X1 RoundFunction_T2_U296 ( .A(RoundFunction_STATE2[186]), .B(
        RoundFunction_T2_n367), .ZN(RoundFunction_TMP3_2[154]) );
  XNOR2_X1 RoundFunction_T2_U295 ( .A(RoundFunction_STATE2[185]), .B(
        RoundFunction_T2_n366), .ZN(RoundFunction_TMP3_2[153]) );
  XNOR2_X1 RoundFunction_T2_U294 ( .A(RoundFunction_STATE2[184]), .B(
        RoundFunction_T2_n365), .ZN(RoundFunction_TMP3_2[152]) );
  XNOR2_X1 RoundFunction_T2_U293 ( .A(RoundFunction_STATE2[183]), .B(
        RoundFunction_T2_n364), .ZN(RoundFunction_TMP3_2[76]) );
  XNOR2_X1 RoundFunction_T2_U292 ( .A(RoundFunction_STATE2[182]), .B(
        RoundFunction_T2_n363), .ZN(RoundFunction_TMP3_2[75]) );
  XNOR2_X1 RoundFunction_T2_U291 ( .A(RoundFunction_STATE2[181]), .B(
        RoundFunction_T2_n362), .ZN(RoundFunction_TMP3_2[74]) );
  XNOR2_X1 RoundFunction_T2_U290 ( .A(RoundFunction_STATE2[180]), .B(
        RoundFunction_T2_n361), .ZN(RoundFunction_TMP3_2[73]) );
  XNOR2_X1 RoundFunction_T2_U289 ( .A(RoundFunction_STATE2[17]), .B(
        RoundFunction_T2_n397), .ZN(RoundFunction_TMP3_2[167]) );
  XNOR2_X1 RoundFunction_T2_U288 ( .A(RoundFunction_STATE2[179]), .B(
        RoundFunction_T2_n399), .ZN(RoundFunction_TMP3_2[72]) );
  XNOR2_X1 RoundFunction_T2_U287 ( .A(RoundFunction_STATE2[178]), .B(
        RoundFunction_T2_n398), .ZN(RoundFunction_TMP3_2[79]) );
  XNOR2_X1 RoundFunction_T2_U286 ( .A(RoundFunction_STATE2[177]), .B(
        RoundFunction_T2_n397), .ZN(RoundFunction_TMP3_2[78]) );
  XNOR2_X1 RoundFunction_T2_U285 ( .A(RoundFunction_STATE2[176]), .B(
        RoundFunction_T2_n396), .ZN(RoundFunction_TMP3_2[77]) );
  XNOR2_X1 RoundFunction_T2_U284 ( .A(RoundFunction_STATE2[175]), .B(
        RoundFunction_T2_n395), .ZN(RoundFunction_TMP3_2[193]) );
  XNOR2_X1 RoundFunction_T2_U283 ( .A(RoundFunction_STATE2[174]), .B(
        RoundFunction_T2_n394), .ZN(RoundFunction_TMP3_2[192]) );
  XNOR2_X1 RoundFunction_T2_U282 ( .A(RoundFunction_STATE2[173]), .B(
        RoundFunction_T2_n393), .ZN(RoundFunction_TMP3_2[199]) );
  XNOR2_X1 RoundFunction_T2_U281 ( .A(RoundFunction_STATE2[172]), .B(
        RoundFunction_T2_n392), .ZN(RoundFunction_TMP3_2[198]) );
  XNOR2_X1 RoundFunction_T2_U280 ( .A(RoundFunction_STATE2[171]), .B(
        RoundFunction_T2_n391), .ZN(RoundFunction_TMP3_2[197]) );
  XNOR2_X1 RoundFunction_T2_U279 ( .A(RoundFunction_STATE2[170]), .B(
        RoundFunction_T2_n390), .ZN(RoundFunction_TMP3_2[196]) );
  XNOR2_X1 RoundFunction_T2_U278 ( .A(RoundFunction_STATE2[16]), .B(
        RoundFunction_T2_n396), .ZN(RoundFunction_TMP3_2[166]) );
  XNOR2_X1 RoundFunction_T2_U277 ( .A(RoundFunction_STATE2[169]), .B(
        RoundFunction_T2_n400), .ZN(RoundFunction_TMP3_2[195]) );
  XNOR2_X1 RoundFunction_T2_U276 ( .A(RoundFunction_STATE2[168]), .B(
        RoundFunction_T2_n389), .ZN(RoundFunction_TMP3_2[194]) );
  XNOR2_X1 RoundFunction_T2_U275 ( .A(RoundFunction_STATE2[167]), .B(
        RoundFunction_T2_n388), .ZN(RoundFunction_TMP3_2[113]) );
  XNOR2_X1 RoundFunction_T2_U274 ( .A(RoundFunction_STATE2[166]), .B(
        RoundFunction_T2_n387), .ZN(RoundFunction_TMP3_2[112]) );
  XNOR2_X1 RoundFunction_T2_U273 ( .A(RoundFunction_STATE2[165]), .B(
        RoundFunction_T2_n386), .ZN(RoundFunction_TMP3_2[119]) );
  XNOR2_X1 RoundFunction_T2_U272 ( .A(RoundFunction_STATE2[164]), .B(
        RoundFunction_T2_n385), .ZN(RoundFunction_TMP3_2[118]) );
  XNOR2_X1 RoundFunction_T2_U271 ( .A(RoundFunction_STATE2[163]), .B(
        RoundFunction_T2_n384), .ZN(RoundFunction_TMP3_2[117]) );
  XNOR2_X1 RoundFunction_T2_U270 ( .A(RoundFunction_STATE2[162]), .B(
        RoundFunction_T2_n383), .ZN(RoundFunction_TMP3_2[116]) );
  XNOR2_X1 RoundFunction_T2_U269 ( .A(RoundFunction_STATE2[161]), .B(
        RoundFunction_T2_n382), .ZN(RoundFunction_TMP3_2[115]) );
  XNOR2_X1 RoundFunction_T2_U268 ( .A(RoundFunction_STATE2[160]), .B(
        RoundFunction_T2_n381), .ZN(RoundFunction_TMP3_2[114]) );
  XNOR2_X1 RoundFunction_T2_U267 ( .A(RoundFunction_STATE2[15]), .B(
        RoundFunction_T2_n395), .ZN(RoundFunction_TMP3_2[80]) );
  XNOR2_X1 RoundFunction_T2_U266 ( .A(RoundFunction_STATE2[159]), .B(
        RoundFunction_T2_n380), .ZN(RoundFunction_TMP3_2[111]) );
  XNOR2_X1 RoundFunction_T2_U265 ( .A(RoundFunction_STATE2[158]), .B(
        RoundFunction_T2_n379), .ZN(RoundFunction_TMP3_2[110]) );
  XNOR2_X1 RoundFunction_T2_U264 ( .A(RoundFunction_STATE2[157]), .B(
        RoundFunction_T2_n378), .ZN(RoundFunction_TMP3_2[109]) );
  XNOR2_X1 RoundFunction_T2_U263 ( .A(RoundFunction_STATE2[156]), .B(
        RoundFunction_T2_n377), .ZN(RoundFunction_TMP3_2[108]) );
  XNOR2_X1 RoundFunction_T2_U262 ( .A(RoundFunction_STATE2[155]), .B(
        RoundFunction_T2_n376), .ZN(RoundFunction_TMP3_2[107]) );
  XNOR2_X1 RoundFunction_T2_U261 ( .A(RoundFunction_STATE2[154]), .B(
        RoundFunction_T2_n375), .ZN(RoundFunction_TMP3_2[106]) );
  XNOR2_X1 RoundFunction_T2_U260 ( .A(RoundFunction_STATE2[153]), .B(
        RoundFunction_T2_n374), .ZN(RoundFunction_TMP3_2[105]) );
  XNOR2_X1 RoundFunction_T2_U259 ( .A(RoundFunction_STATE2[152]), .B(
        RoundFunction_T2_n373), .ZN(RoundFunction_TMP3_2[104]) );
  XNOR2_X1 RoundFunction_T2_U258 ( .A(RoundFunction_STATE2[151]), .B(
        RoundFunction_T2_n372), .ZN(RoundFunction_TMP3_2[28]) );
  XNOR2_X1 RoundFunction_T2_U257 ( .A(RoundFunction_STATE2[150]), .B(
        RoundFunction_T2_n371), .ZN(RoundFunction_TMP3_2[27]) );
  XNOR2_X1 RoundFunction_T2_U256 ( .A(RoundFunction_STATE2[14]), .B(
        RoundFunction_T2_n394), .ZN(RoundFunction_TMP3_2[87]) );
  XNOR2_X1 RoundFunction_T2_U255 ( .A(RoundFunction_STATE2[149]), .B(
        RoundFunction_T2_n370), .ZN(RoundFunction_TMP3_2[26]) );
  XNOR2_X1 RoundFunction_T2_U254 ( .A(RoundFunction_STATE2[148]), .B(
        RoundFunction_T2_n369), .ZN(RoundFunction_TMP3_2[25]) );
  XNOR2_X1 RoundFunction_T2_U253 ( .A(RoundFunction_STATE2[147]), .B(
        RoundFunction_T2_n368), .ZN(RoundFunction_TMP3_2[24]) );
  XNOR2_X1 RoundFunction_T2_U252 ( .A(RoundFunction_STATE2[146]), .B(
        RoundFunction_T2_n367), .ZN(RoundFunction_TMP3_2[31]) );
  XNOR2_X1 RoundFunction_T2_U251 ( .A(RoundFunction_STATE2[145]), .B(
        RoundFunction_T2_n366), .ZN(RoundFunction_TMP3_2[30]) );
  XNOR2_X1 RoundFunction_T2_U250 ( .A(RoundFunction_STATE2[144]), .B(
        RoundFunction_T2_n365), .ZN(RoundFunction_TMP3_2[29]) );
  XNOR2_X1 RoundFunction_T2_U249 ( .A(RoundFunction_STATE2[143]), .B(
        RoundFunction_T2_n364), .ZN(RoundFunction_TMP3_2[150]) );
  XNOR2_X1 RoundFunction_T2_U248 ( .A(RoundFunction_STATE2[142]), .B(
        RoundFunction_T2_n363), .ZN(RoundFunction_TMP3_2[149]) );
  XNOR2_X1 RoundFunction_T2_U247 ( .A(RoundFunction_STATE2[141]), .B(
        RoundFunction_T2_n362), .ZN(RoundFunction_TMP3_2[148]) );
  XNOR2_X1 RoundFunction_T2_U246 ( .A(RoundFunction_STATE2[140]), .B(
        RoundFunction_T2_n361), .ZN(RoundFunction_TMP3_2[147]) );
  XNOR2_X1 RoundFunction_T2_U245 ( .A(RoundFunction_STATE2[13]), .B(
        RoundFunction_T2_n393), .ZN(RoundFunction_TMP3_2[86]) );
  XNOR2_X1 RoundFunction_T2_U244 ( .A(RoundFunction_STATE2[139]), .B(
        RoundFunction_T2_n399), .ZN(RoundFunction_TMP3_2[146]) );
  XNOR2_X1 RoundFunction_T2_U243 ( .A(RoundFunction_T2_n360), .B(
        RoundFunction_T2_n359), .ZN(RoundFunction_T2_n399) );
  XNOR2_X1 RoundFunction_T2_U242 ( .A(RoundFunction_STATE2[138]), .B(
        RoundFunction_T2_n398), .ZN(RoundFunction_TMP3_2[145]) );
  XNOR2_X1 RoundFunction_T2_U241 ( .A(RoundFunction_T2_n358), .B(
        RoundFunction_T2_n357), .ZN(RoundFunction_T2_n398) );
  XNOR2_X1 RoundFunction_T2_U240 ( .A(RoundFunction_STATE2[137]), .B(
        RoundFunction_T2_n397), .ZN(RoundFunction_TMP3_2[144]) );
  XNOR2_X1 RoundFunction_T2_U239 ( .A(RoundFunction_T2_n356), .B(
        RoundFunction_T2_n355), .ZN(RoundFunction_T2_n397) );
  XNOR2_X1 RoundFunction_T2_U238 ( .A(RoundFunction_STATE2[136]), .B(
        RoundFunction_T2_n396), .ZN(RoundFunction_TMP3_2[151]) );
  XNOR2_X1 RoundFunction_T2_U237 ( .A(RoundFunction_T2_n354), .B(
        RoundFunction_T2_n353), .ZN(RoundFunction_T2_n396) );
  XNOR2_X1 RoundFunction_T2_U236 ( .A(RoundFunction_STATE2[135]), .B(
        RoundFunction_T2_n395), .ZN(RoundFunction_TMP3_2[68]) );
  XNOR2_X1 RoundFunction_T2_U235 ( .A(RoundFunction_T2_n352), .B(
        RoundFunction_T2_n351), .ZN(RoundFunction_T2_n395) );
  XNOR2_X1 RoundFunction_T2_U234 ( .A(RoundFunction_STATE2[134]), .B(
        RoundFunction_T2_n394), .ZN(RoundFunction_TMP3_2[67]) );
  XNOR2_X1 RoundFunction_T2_U233 ( .A(RoundFunction_T2_n350), .B(
        RoundFunction_T2_n349), .ZN(RoundFunction_T2_n394) );
  XNOR2_X1 RoundFunction_T2_U232 ( .A(RoundFunction_STATE2[133]), .B(
        RoundFunction_T2_n393), .ZN(RoundFunction_TMP3_2[66]) );
  XNOR2_X1 RoundFunction_T2_U231 ( .A(RoundFunction_T2_n348), .B(
        RoundFunction_T2_n347), .ZN(RoundFunction_T2_n393) );
  XNOR2_X1 RoundFunction_T2_U230 ( .A(RoundFunction_STATE2[132]), .B(
        RoundFunction_T2_n392), .ZN(RoundFunction_TMP3_2[65]) );
  XNOR2_X1 RoundFunction_T2_U229 ( .A(RoundFunction_STATE2[131]), .B(
        RoundFunction_T2_n391), .ZN(RoundFunction_TMP3_2[64]) );
  XNOR2_X1 RoundFunction_T2_U228 ( .A(RoundFunction_STATE2[130]), .B(
        RoundFunction_T2_n390), .ZN(RoundFunction_TMP3_2[71]) );
  XNOR2_X1 RoundFunction_T2_U227 ( .A(RoundFunction_STATE2[12]), .B(
        RoundFunction_T2_n392), .ZN(RoundFunction_TMP3_2[85]) );
  XNOR2_X1 RoundFunction_T2_U226 ( .A(RoundFunction_T2_n346), .B(
        RoundFunction_T2_n345), .ZN(RoundFunction_T2_n392) );
  XNOR2_X1 RoundFunction_T2_U225 ( .A(RoundFunction_STATE2[129]), .B(
        RoundFunction_T2_n400), .ZN(RoundFunction_TMP3_2[70]) );
  XNOR2_X1 RoundFunction_T2_U224 ( .A(RoundFunction_T2_n344), .B(
        RoundFunction_T2_n343), .ZN(RoundFunction_T2_n400) );
  XNOR2_X1 RoundFunction_T2_U223 ( .A(RoundFunction_STATE2[128]), .B(
        RoundFunction_T2_n389), .ZN(RoundFunction_TMP3_2[69]) );
  XNOR2_X1 RoundFunction_T2_U222 ( .A(RoundFunction_T2_n342), .B(
        RoundFunction_T2_n341), .ZN(RoundFunction_T2_n389) );
  XNOR2_X1 RoundFunction_T2_U221 ( .A(RoundFunction_STATE2[127]), .B(
        RoundFunction_T2_n388), .ZN(RoundFunction_TMP3_2[184]) );
  XNOR2_X1 RoundFunction_T2_U220 ( .A(RoundFunction_T2_n340), .B(
        RoundFunction_T2_n339), .ZN(RoundFunction_T2_n388) );
  XNOR2_X1 RoundFunction_T2_U219 ( .A(RoundFunction_STATE2[126]), .B(
        RoundFunction_T2_n387), .ZN(RoundFunction_TMP3_2[191]) );
  XNOR2_X1 RoundFunction_T2_U218 ( .A(RoundFunction_T2_n338), .B(
        RoundFunction_T2_n337), .ZN(RoundFunction_T2_n387) );
  XNOR2_X1 RoundFunction_T2_U217 ( .A(RoundFunction_STATE2[125]), .B(
        RoundFunction_T2_n386), .ZN(RoundFunction_TMP3_2[190]) );
  XNOR2_X1 RoundFunction_T2_U216 ( .A(RoundFunction_T2_n336), .B(
        RoundFunction_T2_n335), .ZN(RoundFunction_T2_n386) );
  XNOR2_X1 RoundFunction_T2_U215 ( .A(RoundFunction_STATE2[124]), .B(
        RoundFunction_T2_n385), .ZN(RoundFunction_TMP3_2[189]) );
  XNOR2_X1 RoundFunction_T2_U214 ( .A(RoundFunction_T2_n334), .B(
        RoundFunction_T2_n359), .ZN(RoundFunction_T2_n385) );
  XOR2_X1 RoundFunction_T2_U213 ( .A(RoundFunction_STATE2[11]), .B(
        RoundFunction_T2_n333), .Z(RoundFunction_T2_n359) );
  XNOR2_X1 RoundFunction_T2_U212 ( .A(RoundFunction_T2_n332), .B(
        RoundFunction_T2_n331), .ZN(RoundFunction_T2_n333) );
  XNOR2_X1 RoundFunction_T2_U211 ( .A(RoundFunction_STATE2[51]), .B(
        RoundFunction_STATE2[91]), .ZN(RoundFunction_T2_n331) );
  XOR2_X1 RoundFunction_T2_U210 ( .A(RoundFunction_STATE2[131]), .B(
        RoundFunction_STATE2[171]), .Z(RoundFunction_T2_n332) );
  XNOR2_X1 RoundFunction_T2_U209 ( .A(RoundFunction_STATE2[123]), .B(
        RoundFunction_T2_n384), .ZN(RoundFunction_TMP3_2[188]) );
  XNOR2_X1 RoundFunction_T2_U208 ( .A(RoundFunction_T2_n330), .B(
        RoundFunction_T2_n357), .ZN(RoundFunction_T2_n384) );
  XOR2_X1 RoundFunction_T2_U207 ( .A(RoundFunction_STATE2[10]), .B(
        RoundFunction_T2_n329), .Z(RoundFunction_T2_n357) );
  XNOR2_X1 RoundFunction_T2_U206 ( .A(RoundFunction_T2_n328), .B(
        RoundFunction_T2_n327), .ZN(RoundFunction_T2_n329) );
  XNOR2_X1 RoundFunction_T2_U205 ( .A(RoundFunction_STATE2[50]), .B(
        RoundFunction_STATE2[90]), .ZN(RoundFunction_T2_n327) );
  XOR2_X1 RoundFunction_T2_U204 ( .A(RoundFunction_STATE2[130]), .B(
        RoundFunction_STATE2[170]), .Z(RoundFunction_T2_n328) );
  XNOR2_X1 RoundFunction_T2_U203 ( .A(RoundFunction_STATE2[122]), .B(
        RoundFunction_T2_n383), .ZN(RoundFunction_TMP3_2[187]) );
  XNOR2_X1 RoundFunction_T2_U202 ( .A(RoundFunction_T2_n326), .B(
        RoundFunction_T2_n355), .ZN(RoundFunction_T2_n383) );
  XOR2_X1 RoundFunction_T2_U201 ( .A(RoundFunction_STATE2[89]), .B(
        RoundFunction_T2_n325), .Z(RoundFunction_T2_n355) );
  XNOR2_X1 RoundFunction_T2_U200 ( .A(RoundFunction_T2_n324), .B(
        RoundFunction_T2_n323), .ZN(RoundFunction_T2_n325) );
  XNOR2_X1 RoundFunction_T2_U199 ( .A(RoundFunction_STATE2[129]), .B(
        RoundFunction_STATE2[49]), .ZN(RoundFunction_T2_n323) );
  XOR2_X1 RoundFunction_T2_U198 ( .A(RoundFunction_STATE2[169]), .B(
        RoundFunction_STATE2[9]), .Z(RoundFunction_T2_n324) );
  XNOR2_X1 RoundFunction_T2_U197 ( .A(RoundFunction_STATE2[121]), .B(
        RoundFunction_T2_n382), .ZN(RoundFunction_TMP3_2[186]) );
  XNOR2_X1 RoundFunction_T2_U196 ( .A(RoundFunction_T2_n322), .B(
        RoundFunction_T2_n353), .ZN(RoundFunction_T2_n382) );
  XOR2_X1 RoundFunction_T2_U195 ( .A(RoundFunction_STATE2[128]), .B(
        RoundFunction_T2_n321), .Z(RoundFunction_T2_n353) );
  XNOR2_X1 RoundFunction_T2_U194 ( .A(RoundFunction_T2_n320), .B(
        RoundFunction_T2_n319), .ZN(RoundFunction_T2_n321) );
  XNOR2_X1 RoundFunction_T2_U193 ( .A(RoundFunction_STATE2[48]), .B(
        RoundFunction_STATE2[8]), .ZN(RoundFunction_T2_n319) );
  XOR2_X1 RoundFunction_T2_U192 ( .A(RoundFunction_STATE2[88]), .B(
        RoundFunction_STATE2[168]), .Z(RoundFunction_T2_n320) );
  XNOR2_X1 RoundFunction_T2_U191 ( .A(RoundFunction_STATE2[120]), .B(
        RoundFunction_T2_n381), .ZN(RoundFunction_TMP3_2[185]) );
  XNOR2_X1 RoundFunction_T2_U190 ( .A(RoundFunction_STATE2[11]), .B(
        RoundFunction_T2_n391), .ZN(RoundFunction_TMP3_2[84]) );
  XNOR2_X1 RoundFunction_T2_U189 ( .A(RoundFunction_T2_n318), .B(
        RoundFunction_T2_n317), .ZN(RoundFunction_T2_n391) );
  XNOR2_X1 RoundFunction_T2_U188 ( .A(RoundFunction_STATE2[119]), .B(
        RoundFunction_T2_n380), .ZN(RoundFunction_TMP3_2[182]) );
  XNOR2_X1 RoundFunction_T2_U187 ( .A(RoundFunction_T2_n354), .B(
        RoundFunction_T2_n349), .ZN(RoundFunction_T2_n380) );
  XOR2_X1 RoundFunction_T2_U186 ( .A(RoundFunction_STATE2[126]), .B(
        RoundFunction_T2_n316), .Z(RoundFunction_T2_n349) );
  XNOR2_X1 RoundFunction_T2_U185 ( .A(RoundFunction_T2_n315), .B(
        RoundFunction_T2_n314), .ZN(RoundFunction_T2_n316) );
  XNOR2_X1 RoundFunction_T2_U184 ( .A(RoundFunction_STATE2[46]), .B(
        RoundFunction_STATE2[86]), .ZN(RoundFunction_T2_n314) );
  XOR2_X1 RoundFunction_T2_U183 ( .A(RoundFunction_STATE2[6]), .B(
        RoundFunction_STATE2[166]), .Z(RoundFunction_T2_n315) );
  XOR2_X1 RoundFunction_T2_U182 ( .A(RoundFunction_STATE2[111]), .B(
        RoundFunction_T2_n313), .Z(RoundFunction_T2_n354) );
  XNOR2_X1 RoundFunction_T2_U181 ( .A(RoundFunction_T2_n312), .B(
        RoundFunction_T2_n311), .ZN(RoundFunction_T2_n313) );
  XNOR2_X1 RoundFunction_T2_U180 ( .A(RoundFunction_STATE2[31]), .B(
        RoundFunction_STATE2[71]), .ZN(RoundFunction_T2_n311) );
  XOR2_X1 RoundFunction_T2_U179 ( .A(RoundFunction_STATE2[151]), .B(
        RoundFunction_STATE2[191]), .Z(RoundFunction_T2_n312) );
  XNOR2_X1 RoundFunction_T2_U178 ( .A(RoundFunction_STATE2[118]), .B(
        RoundFunction_T2_n379), .ZN(RoundFunction_TMP3_2[181]) );
  XNOR2_X1 RoundFunction_T2_U177 ( .A(RoundFunction_T2_n310), .B(
        RoundFunction_T2_n347), .ZN(RoundFunction_T2_n379) );
  XOR2_X1 RoundFunction_T2_U176 ( .A(RoundFunction_STATE2[125]), .B(
        RoundFunction_T2_n309), .Z(RoundFunction_T2_n347) );
  XNOR2_X1 RoundFunction_T2_U175 ( .A(RoundFunction_T2_n308), .B(
        RoundFunction_T2_n307), .ZN(RoundFunction_T2_n309) );
  XNOR2_X1 RoundFunction_T2_U174 ( .A(RoundFunction_STATE2[45]), .B(
        RoundFunction_STATE2[85]), .ZN(RoundFunction_T2_n307) );
  XOR2_X1 RoundFunction_T2_U173 ( .A(RoundFunction_STATE2[5]), .B(
        RoundFunction_STATE2[165]), .Z(RoundFunction_T2_n308) );
  XNOR2_X1 RoundFunction_T2_U172 ( .A(RoundFunction_STATE2[117]), .B(
        RoundFunction_T2_n378), .ZN(RoundFunction_TMP3_2[180]) );
  XNOR2_X1 RoundFunction_T2_U171 ( .A(RoundFunction_T2_n306), .B(
        RoundFunction_T2_n345), .ZN(RoundFunction_T2_n378) );
  XOR2_X1 RoundFunction_T2_U170 ( .A(RoundFunction_STATE2[124]), .B(
        RoundFunction_T2_n305), .Z(RoundFunction_T2_n345) );
  XNOR2_X1 RoundFunction_T2_U169 ( .A(RoundFunction_T2_n304), .B(
        RoundFunction_T2_n303), .ZN(RoundFunction_T2_n305) );
  XNOR2_X1 RoundFunction_T2_U168 ( .A(RoundFunction_STATE2[44]), .B(
        RoundFunction_STATE2[84]), .ZN(RoundFunction_T2_n303) );
  XOR2_X1 RoundFunction_T2_U167 ( .A(RoundFunction_STATE2[4]), .B(
        RoundFunction_STATE2[164]), .Z(RoundFunction_T2_n304) );
  XNOR2_X1 RoundFunction_T2_U166 ( .A(RoundFunction_STATE2[116]), .B(
        RoundFunction_T2_n377), .ZN(RoundFunction_TMP3_2[179]) );
  XNOR2_X1 RoundFunction_T2_U165 ( .A(RoundFunction_T2_n302), .B(
        RoundFunction_T2_n317), .ZN(RoundFunction_T2_n377) );
  XOR2_X1 RoundFunction_T2_U164 ( .A(RoundFunction_STATE2[123]), .B(
        RoundFunction_T2_n301), .Z(RoundFunction_T2_n317) );
  XNOR2_X1 RoundFunction_T2_U163 ( .A(RoundFunction_T2_n300), .B(
        RoundFunction_T2_n299), .ZN(RoundFunction_T2_n301) );
  XNOR2_X1 RoundFunction_T2_U162 ( .A(RoundFunction_STATE2[3]), .B(
        RoundFunction_STATE2[83]), .ZN(RoundFunction_T2_n299) );
  XOR2_X1 RoundFunction_T2_U161 ( .A(RoundFunction_STATE2[43]), .B(
        RoundFunction_STATE2[163]), .Z(RoundFunction_T2_n300) );
  XNOR2_X1 RoundFunction_T2_U160 ( .A(RoundFunction_STATE2[115]), .B(
        RoundFunction_T2_n376), .ZN(RoundFunction_TMP3_2[178]) );
  XNOR2_X1 RoundFunction_T2_U159 ( .A(RoundFunction_T2_n298), .B(
        RoundFunction_T2_n297), .ZN(RoundFunction_T2_n376) );
  XNOR2_X1 RoundFunction_T2_U158 ( .A(RoundFunction_STATE2[114]), .B(
        RoundFunction_T2_n375), .ZN(RoundFunction_TMP3_2[177]) );
  XNOR2_X1 RoundFunction_T2_U157 ( .A(RoundFunction_T2_n343), .B(
        RoundFunction_T2_n360), .ZN(RoundFunction_T2_n375) );
  XOR2_X1 RoundFunction_T2_U156 ( .A(RoundFunction_STATE2[106]), .B(
        RoundFunction_T2_n296), .Z(RoundFunction_T2_n360) );
  XNOR2_X1 RoundFunction_T2_U155 ( .A(RoundFunction_T2_n295), .B(
        RoundFunction_T2_n294), .ZN(RoundFunction_T2_n296) );
  XNOR2_X1 RoundFunction_T2_U154 ( .A(RoundFunction_STATE2[26]), .B(
        RoundFunction_STATE2[66]), .ZN(RoundFunction_T2_n294) );
  XOR2_X1 RoundFunction_T2_U153 ( .A(RoundFunction_STATE2[146]), .B(
        RoundFunction_STATE2[186]), .Z(RoundFunction_T2_n295) );
  XOR2_X1 RoundFunction_T2_U152 ( .A(RoundFunction_STATE2[121]), .B(
        RoundFunction_T2_n293), .Z(RoundFunction_T2_n343) );
  XNOR2_X1 RoundFunction_T2_U151 ( .A(RoundFunction_T2_n292), .B(
        RoundFunction_T2_n291), .ZN(RoundFunction_T2_n293) );
  XNOR2_X1 RoundFunction_T2_U150 ( .A(RoundFunction_STATE2[1]), .B(
        RoundFunction_STATE2[81]), .ZN(RoundFunction_T2_n291) );
  XOR2_X1 RoundFunction_T2_U149 ( .A(RoundFunction_STATE2[41]), .B(
        RoundFunction_STATE2[161]), .Z(RoundFunction_T2_n292) );
  XNOR2_X1 RoundFunction_T2_U148 ( .A(RoundFunction_STATE2[113]), .B(
        RoundFunction_T2_n374), .ZN(RoundFunction_TMP3_2[176]) );
  XNOR2_X1 RoundFunction_T2_U147 ( .A(RoundFunction_T2_n358), .B(
        RoundFunction_T2_n341), .ZN(RoundFunction_T2_n374) );
  XOR2_X1 RoundFunction_T2_U146 ( .A(RoundFunction_STATE2[0]), .B(
        RoundFunction_T2_n290), .Z(RoundFunction_T2_n341) );
  XNOR2_X1 RoundFunction_T2_U145 ( .A(RoundFunction_T2_n289), .B(
        RoundFunction_T2_n288), .ZN(RoundFunction_T2_n290) );
  XNOR2_X1 RoundFunction_T2_U144 ( .A(RoundFunction_STATE2[40]), .B(
        RoundFunction_STATE2[80]), .ZN(RoundFunction_T2_n288) );
  XOR2_X1 RoundFunction_T2_U143 ( .A(RoundFunction_STATE2[120]), .B(
        RoundFunction_STATE2[160]), .Z(RoundFunction_T2_n289) );
  XOR2_X1 RoundFunction_T2_U142 ( .A(RoundFunction_STATE2[105]), .B(
        RoundFunction_T2_n287), .Z(RoundFunction_T2_n358) );
  XNOR2_X1 RoundFunction_T2_U141 ( .A(RoundFunction_T2_n286), .B(
        RoundFunction_T2_n285), .ZN(RoundFunction_T2_n287) );
  XNOR2_X1 RoundFunction_T2_U140 ( .A(RoundFunction_STATE2[25]), .B(
        RoundFunction_STATE2[65]), .ZN(RoundFunction_T2_n285) );
  XOR2_X1 RoundFunction_T2_U139 ( .A(RoundFunction_STATE2[145]), .B(
        RoundFunction_STATE2[185]), .Z(RoundFunction_T2_n286) );
  XNOR2_X1 RoundFunction_T2_U138 ( .A(RoundFunction_STATE2[112]), .B(
        RoundFunction_T2_n373), .ZN(RoundFunction_TMP3_2[183]) );
  XNOR2_X1 RoundFunction_T2_U137 ( .A(RoundFunction_T2_n356), .B(
        RoundFunction_T2_n351), .ZN(RoundFunction_T2_n373) );
  XOR2_X1 RoundFunction_T2_U136 ( .A(RoundFunction_STATE2[127]), .B(
        RoundFunction_T2_n284), .Z(RoundFunction_T2_n351) );
  XNOR2_X1 RoundFunction_T2_U135 ( .A(RoundFunction_T2_n283), .B(
        RoundFunction_T2_n282), .ZN(RoundFunction_T2_n284) );
  XNOR2_X1 RoundFunction_T2_U134 ( .A(RoundFunction_STATE2[47]), .B(
        RoundFunction_STATE2[87]), .ZN(RoundFunction_T2_n282) );
  XOR2_X1 RoundFunction_T2_U133 ( .A(RoundFunction_STATE2[7]), .B(
        RoundFunction_STATE2[167]), .Z(RoundFunction_T2_n283) );
  XOR2_X1 RoundFunction_T2_U132 ( .A(RoundFunction_STATE2[104]), .B(
        RoundFunction_T2_n281), .Z(RoundFunction_T2_n356) );
  XNOR2_X1 RoundFunction_T2_U131 ( .A(RoundFunction_T2_n280), .B(
        RoundFunction_T2_n279), .ZN(RoundFunction_T2_n281) );
  XNOR2_X1 RoundFunction_T2_U130 ( .A(RoundFunction_STATE2[24]), .B(
        RoundFunction_STATE2[64]), .ZN(RoundFunction_T2_n279) );
  XOR2_X1 RoundFunction_T2_U129 ( .A(RoundFunction_STATE2[144]), .B(
        RoundFunction_STATE2[184]), .Z(RoundFunction_T2_n280) );
  XNOR2_X1 RoundFunction_T2_U128 ( .A(RoundFunction_STATE2[111]), .B(
        RoundFunction_T2_n372), .ZN(RoundFunction_TMP3_2[96]) );
  XNOR2_X1 RoundFunction_T2_U127 ( .A(RoundFunction_T2_n342), .B(
        RoundFunction_T2_n337), .ZN(RoundFunction_T2_n372) );
  XOR2_X1 RoundFunction_T2_U126 ( .A(RoundFunction_STATE2[118]), .B(
        RoundFunction_T2_n278), .Z(RoundFunction_T2_n337) );
  XNOR2_X1 RoundFunction_T2_U125 ( .A(RoundFunction_T2_n277), .B(
        RoundFunction_T2_n276), .ZN(RoundFunction_T2_n278) );
  XNOR2_X1 RoundFunction_T2_U124 ( .A(RoundFunction_STATE2[198]), .B(
        RoundFunction_STATE2[78]), .ZN(RoundFunction_T2_n276) );
  XOR2_X1 RoundFunction_T2_U123 ( .A(RoundFunction_STATE2[38]), .B(
        RoundFunction_STATE2[158]), .Z(RoundFunction_T2_n277) );
  XOR2_X1 RoundFunction_T2_U122 ( .A(RoundFunction_STATE2[103]), .B(
        RoundFunction_T2_n275), .Z(RoundFunction_T2_n342) );
  XNOR2_X1 RoundFunction_T2_U121 ( .A(RoundFunction_T2_n274), .B(
        RoundFunction_T2_n273), .ZN(RoundFunction_T2_n275) );
  XNOR2_X1 RoundFunction_T2_U120 ( .A(RoundFunction_STATE2[23]), .B(
        RoundFunction_STATE2[63]), .ZN(RoundFunction_T2_n273) );
  XOR2_X1 RoundFunction_T2_U119 ( .A(RoundFunction_STATE2[143]), .B(
        RoundFunction_STATE2[183]), .Z(RoundFunction_T2_n274) );
  XNOR2_X1 RoundFunction_T2_U118 ( .A(RoundFunction_STATE2[110]), .B(
        RoundFunction_T2_n371), .ZN(RoundFunction_TMP3_2[103]) );
  XNOR2_X1 RoundFunction_T2_U117 ( .A(RoundFunction_T2_n352), .B(
        RoundFunction_T2_n335), .ZN(RoundFunction_T2_n371) );
  XOR2_X1 RoundFunction_T2_U116 ( .A(RoundFunction_STATE2[117]), .B(
        RoundFunction_T2_n272), .Z(RoundFunction_T2_n335) );
  XNOR2_X1 RoundFunction_T2_U115 ( .A(RoundFunction_T2_n271), .B(
        RoundFunction_T2_n270), .ZN(RoundFunction_T2_n272) );
  XNOR2_X1 RoundFunction_T2_U114 ( .A(RoundFunction_STATE2[197]), .B(
        RoundFunction_STATE2[77]), .ZN(RoundFunction_T2_n270) );
  XOR2_X1 RoundFunction_T2_U113 ( .A(RoundFunction_STATE2[37]), .B(
        RoundFunction_STATE2[157]), .Z(RoundFunction_T2_n271) );
  XOR2_X1 RoundFunction_T2_U112 ( .A(RoundFunction_STATE2[102]), .B(
        RoundFunction_T2_n269), .Z(RoundFunction_T2_n352) );
  XNOR2_X1 RoundFunction_T2_U111 ( .A(RoundFunction_T2_n268), .B(
        RoundFunction_T2_n267), .ZN(RoundFunction_T2_n269) );
  XNOR2_X1 RoundFunction_T2_U110 ( .A(RoundFunction_STATE2[22]), .B(
        RoundFunction_STATE2[62]), .ZN(RoundFunction_T2_n267) );
  XOR2_X1 RoundFunction_T2_U109 ( .A(RoundFunction_STATE2[142]), .B(
        RoundFunction_STATE2[182]), .Z(RoundFunction_T2_n268) );
  XNOR2_X1 RoundFunction_T2_U108 ( .A(RoundFunction_STATE2[10]), .B(
        RoundFunction_T2_n390), .ZN(RoundFunction_TMP3_2[83]) );
  XNOR2_X1 RoundFunction_T2_U107 ( .A(RoundFunction_T2_n266), .B(
        RoundFunction_T2_n297), .ZN(RoundFunction_T2_n390) );
  XOR2_X1 RoundFunction_T2_U106 ( .A(RoundFunction_STATE2[122]), .B(
        RoundFunction_T2_n265), .Z(RoundFunction_T2_n297) );
  XNOR2_X1 RoundFunction_T2_U105 ( .A(RoundFunction_T2_n264), .B(
        RoundFunction_T2_n263), .ZN(RoundFunction_T2_n265) );
  XNOR2_X1 RoundFunction_T2_U104 ( .A(RoundFunction_STATE2[2]), .B(
        RoundFunction_STATE2[82]), .ZN(RoundFunction_T2_n263) );
  XOR2_X1 RoundFunction_T2_U103 ( .A(RoundFunction_STATE2[42]), .B(
        RoundFunction_STATE2[162]), .Z(RoundFunction_T2_n264) );
  XNOR2_X1 RoundFunction_T2_U102 ( .A(RoundFunction_STATE2[109]), .B(
        RoundFunction_T2_n370), .ZN(RoundFunction_TMP3_2[102]) );
  XNOR2_X1 RoundFunction_T2_U101 ( .A(RoundFunction_T2_n350), .B(
        RoundFunction_T2_n334), .ZN(RoundFunction_T2_n370) );
  XOR2_X1 RoundFunction_T2_U100 ( .A(RoundFunction_STATE2[116]), .B(
        RoundFunction_T2_n262), .Z(RoundFunction_T2_n334) );
  XNOR2_X1 RoundFunction_T2_U99 ( .A(RoundFunction_T2_n261), .B(
        RoundFunction_T2_n260), .ZN(RoundFunction_T2_n262) );
  XNOR2_X1 RoundFunction_T2_U98 ( .A(RoundFunction_STATE2[196]), .B(
        RoundFunction_STATE2[76]), .ZN(RoundFunction_T2_n260) );
  XOR2_X1 RoundFunction_T2_U97 ( .A(RoundFunction_STATE2[36]), .B(
        RoundFunction_STATE2[156]), .Z(RoundFunction_T2_n261) );
  XOR2_X1 RoundFunction_T2_U96 ( .A(RoundFunction_STATE2[101]), .B(
        RoundFunction_T2_n259), .Z(RoundFunction_T2_n350) );
  XNOR2_X1 RoundFunction_T2_U95 ( .A(RoundFunction_T2_n258), .B(
        RoundFunction_T2_n257), .ZN(RoundFunction_T2_n259) );
  XNOR2_X1 RoundFunction_T2_U94 ( .A(RoundFunction_STATE2[21]), .B(
        RoundFunction_STATE2[61]), .ZN(RoundFunction_T2_n257) );
  XOR2_X1 RoundFunction_T2_U93 ( .A(RoundFunction_STATE2[141]), .B(
        RoundFunction_STATE2[181]), .Z(RoundFunction_T2_n258) );
  XNOR2_X1 RoundFunction_T2_U92 ( .A(RoundFunction_STATE2[108]), .B(
        RoundFunction_T2_n369), .ZN(RoundFunction_TMP3_2[101]) );
  XNOR2_X1 RoundFunction_T2_U91 ( .A(RoundFunction_T2_n348), .B(
        RoundFunction_T2_n330), .ZN(RoundFunction_T2_n369) );
  XOR2_X1 RoundFunction_T2_U90 ( .A(RoundFunction_STATE2[115]), .B(
        RoundFunction_T2_n256), .Z(RoundFunction_T2_n330) );
  XNOR2_X1 RoundFunction_T2_U89 ( .A(RoundFunction_T2_n255), .B(
        RoundFunction_T2_n254), .ZN(RoundFunction_T2_n256) );
  XNOR2_X1 RoundFunction_T2_U88 ( .A(RoundFunction_STATE2[195]), .B(
        RoundFunction_STATE2[75]), .ZN(RoundFunction_T2_n254) );
  XOR2_X1 RoundFunction_T2_U87 ( .A(RoundFunction_STATE2[35]), .B(
        RoundFunction_STATE2[155]), .Z(RoundFunction_T2_n255) );
  XOR2_X1 RoundFunction_T2_U86 ( .A(RoundFunction_STATE2[100]), .B(
        RoundFunction_T2_n253), .Z(RoundFunction_T2_n348) );
  XNOR2_X1 RoundFunction_T2_U85 ( .A(RoundFunction_T2_n252), .B(
        RoundFunction_T2_n251), .ZN(RoundFunction_T2_n253) );
  XNOR2_X1 RoundFunction_T2_U84 ( .A(RoundFunction_STATE2[20]), .B(
        RoundFunction_STATE2[60]), .ZN(RoundFunction_T2_n251) );
  XOR2_X1 RoundFunction_T2_U83 ( .A(RoundFunction_STATE2[140]), .B(
        RoundFunction_STATE2[180]), .Z(RoundFunction_T2_n252) );
  XNOR2_X1 RoundFunction_T2_U82 ( .A(RoundFunction_STATE2[107]), .B(
        RoundFunction_T2_n368), .ZN(RoundFunction_TMP3_2[100]) );
  XNOR2_X1 RoundFunction_T2_U81 ( .A(RoundFunction_T2_n346), .B(
        RoundFunction_T2_n326), .ZN(RoundFunction_T2_n368) );
  XOR2_X1 RoundFunction_T2_U80 ( .A(RoundFunction_STATE2[114]), .B(
        RoundFunction_T2_n250), .Z(RoundFunction_T2_n326) );
  XNOR2_X1 RoundFunction_T2_U79 ( .A(RoundFunction_T2_n249), .B(
        RoundFunction_T2_n248), .ZN(RoundFunction_T2_n250) );
  XNOR2_X1 RoundFunction_T2_U78 ( .A(RoundFunction_STATE2[194]), .B(
        RoundFunction_STATE2[74]), .ZN(RoundFunction_T2_n248) );
  XOR2_X1 RoundFunction_T2_U77 ( .A(RoundFunction_STATE2[34]), .B(
        RoundFunction_STATE2[154]), .Z(RoundFunction_T2_n249) );
  XOR2_X1 RoundFunction_T2_U76 ( .A(RoundFunction_STATE2[59]), .B(
        RoundFunction_T2_n247), .Z(RoundFunction_T2_n346) );
  XNOR2_X1 RoundFunction_T2_U75 ( .A(RoundFunction_T2_n246), .B(
        RoundFunction_T2_n245), .ZN(RoundFunction_T2_n247) );
  XNOR2_X1 RoundFunction_T2_U74 ( .A(RoundFunction_STATE2[139]), .B(
        RoundFunction_STATE2[19]), .ZN(RoundFunction_T2_n245) );
  XOR2_X1 RoundFunction_T2_U73 ( .A(RoundFunction_STATE2[179]), .B(
        RoundFunction_STATE2[99]), .Z(RoundFunction_T2_n246) );
  XNOR2_X1 RoundFunction_T2_U72 ( .A(RoundFunction_STATE2[106]), .B(
        RoundFunction_T2_n367), .ZN(RoundFunction_TMP3_2[99]) );
  XNOR2_X1 RoundFunction_T2_U71 ( .A(RoundFunction_T2_n318), .B(
        RoundFunction_T2_n322), .ZN(RoundFunction_T2_n367) );
  XOR2_X1 RoundFunction_T2_U70 ( .A(RoundFunction_STATE2[113]), .B(
        RoundFunction_T2_n244), .Z(RoundFunction_T2_n322) );
  XNOR2_X1 RoundFunction_T2_U69 ( .A(RoundFunction_T2_n243), .B(
        RoundFunction_T2_n242), .ZN(RoundFunction_T2_n244) );
  XNOR2_X1 RoundFunction_T2_U68 ( .A(RoundFunction_STATE2[193]), .B(
        RoundFunction_STATE2[73]), .ZN(RoundFunction_T2_n242) );
  XOR2_X1 RoundFunction_T2_U67 ( .A(RoundFunction_STATE2[33]), .B(
        RoundFunction_STATE2[153]), .Z(RoundFunction_T2_n243) );
  XOR2_X1 RoundFunction_T2_U66 ( .A(RoundFunction_STATE2[58]), .B(
        RoundFunction_T2_n241), .Z(RoundFunction_T2_n318) );
  XNOR2_X1 RoundFunction_T2_U65 ( .A(RoundFunction_T2_n240), .B(
        RoundFunction_T2_n239), .ZN(RoundFunction_T2_n241) );
  XNOR2_X1 RoundFunction_T2_U64 ( .A(RoundFunction_STATE2[138]), .B(
        RoundFunction_STATE2[18]), .ZN(RoundFunction_T2_n239) );
  XOR2_X1 RoundFunction_T2_U63 ( .A(RoundFunction_STATE2[178]), .B(
        RoundFunction_STATE2[98]), .Z(RoundFunction_T2_n240) );
  XNOR2_X1 RoundFunction_T2_U62 ( .A(RoundFunction_STATE2[105]), .B(
        RoundFunction_T2_n366), .ZN(RoundFunction_TMP3_2[98]) );
  XNOR2_X1 RoundFunction_T2_U61 ( .A(RoundFunction_T2_n238), .B(
        RoundFunction_T2_n266), .ZN(RoundFunction_T2_n366) );
  XOR2_X1 RoundFunction_T2_U60 ( .A(RoundFunction_STATE2[57]), .B(
        RoundFunction_T2_n237), .Z(RoundFunction_T2_n266) );
  XNOR2_X1 RoundFunction_T2_U59 ( .A(RoundFunction_T2_n236), .B(
        RoundFunction_T2_n235), .ZN(RoundFunction_T2_n237) );
  XNOR2_X1 RoundFunction_T2_U58 ( .A(RoundFunction_STATE2[137]), .B(
        RoundFunction_STATE2[17]), .ZN(RoundFunction_T2_n235) );
  XOR2_X1 RoundFunction_T2_U57 ( .A(RoundFunction_STATE2[177]), .B(
        RoundFunction_STATE2[97]), .Z(RoundFunction_T2_n236) );
  XNOR2_X1 RoundFunction_T2_U56 ( .A(RoundFunction_STATE2[104]), .B(
        RoundFunction_T2_n365), .ZN(RoundFunction_TMP3_2[97]) );
  XNOR2_X1 RoundFunction_T2_U55 ( .A(RoundFunction_T2_n344), .B(
        RoundFunction_T2_n339), .ZN(RoundFunction_T2_n365) );
  XOR2_X1 RoundFunction_T2_U54 ( .A(RoundFunction_STATE2[119]), .B(
        RoundFunction_T2_n234), .Z(RoundFunction_T2_n339) );
  XNOR2_X1 RoundFunction_T2_U53 ( .A(RoundFunction_T2_n233), .B(
        RoundFunction_T2_n232), .ZN(RoundFunction_T2_n234) );
  XNOR2_X1 RoundFunction_T2_U52 ( .A(RoundFunction_STATE2[199]), .B(
        RoundFunction_STATE2[79]), .ZN(RoundFunction_T2_n232) );
  XOR2_X1 RoundFunction_T2_U51 ( .A(RoundFunction_STATE2[39]), .B(
        RoundFunction_STATE2[159]), .Z(RoundFunction_T2_n233) );
  XOR2_X1 RoundFunction_T2_U50 ( .A(RoundFunction_STATE2[136]), .B(
        RoundFunction_T2_n231), .Z(RoundFunction_T2_n344) );
  XNOR2_X1 RoundFunction_T2_U49 ( .A(RoundFunction_T2_n230), .B(
        RoundFunction_T2_n229), .ZN(RoundFunction_T2_n231) );
  XNOR2_X1 RoundFunction_T2_U48 ( .A(RoundFunction_STATE2[176]), .B(
        RoundFunction_STATE2[96]), .ZN(RoundFunction_T2_n229) );
  XOR2_X1 RoundFunction_T2_U47 ( .A(RoundFunction_STATE2[56]), .B(
        RoundFunction_STATE2[16]), .Z(RoundFunction_T2_n230) );
  XNOR2_X1 RoundFunction_T2_U46 ( .A(RoundFunction_STATE2[103]), .B(
        RoundFunction_T2_n364), .ZN(RoundFunction_TMP3_2[18]) );
  XNOR2_X1 RoundFunction_T2_U45 ( .A(RoundFunction_T2_n228), .B(
        RoundFunction_T2_n310), .ZN(RoundFunction_T2_n364) );
  XOR2_X1 RoundFunction_T2_U44 ( .A(RoundFunction_STATE2[110]), .B(
        RoundFunction_T2_n227), .Z(RoundFunction_T2_n310) );
  XNOR2_X1 RoundFunction_T2_U43 ( .A(RoundFunction_T2_n226), .B(
        RoundFunction_T2_n225), .ZN(RoundFunction_T2_n227) );
  XNOR2_X1 RoundFunction_T2_U42 ( .A(RoundFunction_STATE2[190]), .B(
        RoundFunction_STATE2[70]), .ZN(RoundFunction_T2_n225) );
  XOR2_X1 RoundFunction_T2_U41 ( .A(RoundFunction_STATE2[30]), .B(
        RoundFunction_STATE2[150]), .Z(RoundFunction_T2_n226) );
  XNOR2_X1 RoundFunction_T2_U40 ( .A(RoundFunction_STATE2[102]), .B(
        RoundFunction_T2_n363), .ZN(RoundFunction_TMP3_2[17]) );
  XNOR2_X1 RoundFunction_T2_U39 ( .A(RoundFunction_T2_n340), .B(
        RoundFunction_T2_n306), .ZN(RoundFunction_T2_n363) );
  XOR2_X1 RoundFunction_T2_U38 ( .A(RoundFunction_STATE2[109]), .B(
        RoundFunction_T2_n224), .Z(RoundFunction_T2_n306) );
  XNOR2_X1 RoundFunction_T2_U37 ( .A(RoundFunction_T2_n223), .B(
        RoundFunction_T2_n222), .ZN(RoundFunction_T2_n224) );
  XNOR2_X1 RoundFunction_T2_U36 ( .A(RoundFunction_STATE2[189]), .B(
        RoundFunction_STATE2[69]), .ZN(RoundFunction_T2_n222) );
  XOR2_X1 RoundFunction_T2_U35 ( .A(RoundFunction_STATE2[29]), .B(
        RoundFunction_STATE2[149]), .Z(RoundFunction_T2_n223) );
  XOR2_X1 RoundFunction_T2_U34 ( .A(RoundFunction_STATE2[54]), .B(
        RoundFunction_T2_n221), .Z(RoundFunction_T2_n340) );
  XNOR2_X1 RoundFunction_T2_U33 ( .A(RoundFunction_T2_n220), .B(
        RoundFunction_T2_n219), .ZN(RoundFunction_T2_n221) );
  XNOR2_X1 RoundFunction_T2_U32 ( .A(RoundFunction_STATE2[134]), .B(
        RoundFunction_STATE2[174]), .ZN(RoundFunction_T2_n219) );
  XOR2_X1 RoundFunction_T2_U31 ( .A(RoundFunction_STATE2[14]), .B(
        RoundFunction_STATE2[94]), .Z(RoundFunction_T2_n220) );
  XNOR2_X1 RoundFunction_T2_U30 ( .A(RoundFunction_STATE2[101]), .B(
        RoundFunction_T2_n362), .ZN(RoundFunction_TMP3_2[16]) );
  XNOR2_X1 RoundFunction_T2_U29 ( .A(RoundFunction_T2_n338), .B(
        RoundFunction_T2_n302), .ZN(RoundFunction_T2_n362) );
  XOR2_X1 RoundFunction_T2_U28 ( .A(RoundFunction_STATE2[108]), .B(
        RoundFunction_T2_n218), .Z(RoundFunction_T2_n302) );
  XNOR2_X1 RoundFunction_T2_U27 ( .A(RoundFunction_T2_n217), .B(
        RoundFunction_T2_n216), .ZN(RoundFunction_T2_n218) );
  XNOR2_X1 RoundFunction_T2_U26 ( .A(RoundFunction_STATE2[188]), .B(
        RoundFunction_STATE2[68]), .ZN(RoundFunction_T2_n216) );
  XOR2_X1 RoundFunction_T2_U25 ( .A(RoundFunction_STATE2[28]), .B(
        RoundFunction_STATE2[148]), .Z(RoundFunction_T2_n217) );
  XOR2_X1 RoundFunction_T2_U24 ( .A(RoundFunction_STATE2[53]), .B(
        RoundFunction_T2_n215), .Z(RoundFunction_T2_n338) );
  XNOR2_X1 RoundFunction_T2_U23 ( .A(RoundFunction_T2_n214), .B(
        RoundFunction_T2_n213), .ZN(RoundFunction_T2_n215) );
  XNOR2_X1 RoundFunction_T2_U22 ( .A(RoundFunction_STATE2[133]), .B(
        RoundFunction_STATE2[173]), .ZN(RoundFunction_T2_n213) );
  XOR2_X1 RoundFunction_T2_U21 ( .A(RoundFunction_STATE2[13]), .B(
        RoundFunction_STATE2[93]), .Z(RoundFunction_T2_n214) );
  XNOR2_X1 RoundFunction_T2_U20 ( .A(RoundFunction_STATE2[100]), .B(
        RoundFunction_T2_n361), .ZN(RoundFunction_TMP3_2[23]) );
  XNOR2_X1 RoundFunction_T2_U19 ( .A(RoundFunction_T2_n336), .B(
        RoundFunction_T2_n298), .ZN(RoundFunction_T2_n361) );
  XOR2_X1 RoundFunction_T2_U18 ( .A(RoundFunction_STATE2[107]), .B(
        RoundFunction_T2_n212), .Z(RoundFunction_T2_n298) );
  XNOR2_X1 RoundFunction_T2_U17 ( .A(RoundFunction_T2_n211), .B(
        RoundFunction_T2_n210), .ZN(RoundFunction_T2_n212) );
  XNOR2_X1 RoundFunction_T2_U16 ( .A(RoundFunction_STATE2[187]), .B(
        RoundFunction_STATE2[67]), .ZN(RoundFunction_T2_n210) );
  XOR2_X1 RoundFunction_T2_U15 ( .A(RoundFunction_STATE2[27]), .B(
        RoundFunction_STATE2[147]), .Z(RoundFunction_T2_n211) );
  XOR2_X1 RoundFunction_T2_U14 ( .A(RoundFunction_STATE2[52]), .B(
        RoundFunction_T2_n209), .Z(RoundFunction_T2_n336) );
  XNOR2_X1 RoundFunction_T2_U13 ( .A(RoundFunction_T2_n208), .B(
        RoundFunction_T2_n207), .ZN(RoundFunction_T2_n209) );
  XNOR2_X1 RoundFunction_T2_U12 ( .A(RoundFunction_STATE2[12]), .B(
        RoundFunction_STATE2[172]), .ZN(RoundFunction_T2_n207) );
  XOR2_X1 RoundFunction_T2_U11 ( .A(RoundFunction_STATE2[132]), .B(
        RoundFunction_STATE2[92]), .Z(RoundFunction_T2_n208) );
  XNOR2_X1 RoundFunction_T2_U10 ( .A(RoundFunction_STATE2[0]), .B(
        RoundFunction_T2_n381), .ZN(RoundFunction_TMP3_2[0]) );
  XNOR2_X1 RoundFunction_T2_U9 ( .A(RoundFunction_T2_n238), .B(
        RoundFunction_T2_n228), .ZN(RoundFunction_T2_n381) );
  XOR2_X1 RoundFunction_T2_U8 ( .A(RoundFunction_STATE2[55]), .B(
        RoundFunction_T2_n206), .Z(RoundFunction_T2_n228) );
  XNOR2_X1 RoundFunction_T2_U7 ( .A(RoundFunction_T2_n205), .B(
        RoundFunction_T2_n204), .ZN(RoundFunction_T2_n206) );
  XNOR2_X1 RoundFunction_T2_U6 ( .A(RoundFunction_STATE2[135]), .B(
        RoundFunction_STATE2[175]), .ZN(RoundFunction_T2_n204) );
  XOR2_X1 RoundFunction_T2_U5 ( .A(RoundFunction_STATE2[15]), .B(
        RoundFunction_STATE2[95]), .Z(RoundFunction_T2_n205) );
  XOR2_X1 RoundFunction_T2_U4 ( .A(RoundFunction_STATE2[112]), .B(
        RoundFunction_T2_n203), .Z(RoundFunction_T2_n238) );
  XNOR2_X1 RoundFunction_T2_U3 ( .A(RoundFunction_T2_n202), .B(
        RoundFunction_T2_n201), .ZN(RoundFunction_T2_n203) );
  XNOR2_X1 RoundFunction_T2_U2 ( .A(RoundFunction_STATE2[192]), .B(
        RoundFunction_STATE2[72]), .ZN(RoundFunction_T2_n201) );
  XOR2_X1 RoundFunction_T2_U1 ( .A(RoundFunction_STATE2[32]), .B(
        RoundFunction_STATE2[152]), .Z(RoundFunction_T2_n202) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_0_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[16]), .CK(RoundFunction_C_Inst_Chi_NoFresh_0_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[16]), .CK(RoundFunction_C_Inst_Chi_NoFresh_0_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[24]), .CK(RoundFunction_C_Inst_Chi_NoFresh_0_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[24]), .CK(RoundFunction_C_Inst_Chi_NoFresh_0_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[32]), .CK(RoundFunction_C_Inst_Chi_NoFresh_0_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[32]), .CK(RoundFunction_C_Inst_Chi_NoFresh_0_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[0]), .CK(RoundFunction_C_Inst_Chi_NoFresh_0_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[0]), .CK(RoundFunction_C_Inst_Chi_NoFresh_0_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[8]), .CK(RoundFunction_C_Inst_Chi_NoFresh_0_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[8]), .CK(RoundFunction_C_Inst_Chi_NoFresh_0_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[1]), .Z(RESULT1[160]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[3]), .Z(RESULT2[160]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[5]), .Z(RESULT1[168]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[7]), .Z(RESULT2[168]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[9]), .Z(RESULT1[176]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[11]), .Z(RESULT2[176]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[13]), .Z(RESULT1[184]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[15]), .Z(RESULT2[184]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[17]), .Z(
        RoundFunction_TMP4_1[0]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[19]), .Z(RESULT2[192]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_1_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[17]), .CK(RoundFunction_C_Inst_Chi_NoFresh_1_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[17]), .CK(RoundFunction_C_Inst_Chi_NoFresh_1_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[25]), .CK(RoundFunction_C_Inst_Chi_NoFresh_1_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[33]), .CK(RoundFunction_C_Inst_Chi_NoFresh_1_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[33]), .CK(RoundFunction_C_Inst_Chi_NoFresh_1_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[1]), .CK(RoundFunction_C_Inst_Chi_NoFresh_1_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[1]), .CK(RoundFunction_C_Inst_Chi_NoFresh_1_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[9]), .CK(RoundFunction_C_Inst_Chi_NoFresh_1_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[9]), .CK(RoundFunction_C_Inst_Chi_NoFresh_1_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[1]), .Z(RESULT1[161]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[3]), .Z(RESULT2[161]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[5]), .Z(RESULT1[169]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[7]), .Z(RESULT2[169]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[9]), .Z(RESULT1[177]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[11]), .Z(RESULT2[177]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[13]), .Z(RESULT1[185]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[15]), .Z(RESULT2[185]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[17]), .Z(
        RoundFunction_TMP4_1[1]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[19]), .Z(RESULT2[193]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_2_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[18]), .CK(RoundFunction_C_Inst_Chi_NoFresh_2_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[18]), .CK(RoundFunction_C_Inst_Chi_NoFresh_2_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[26]), .CK(RoundFunction_C_Inst_Chi_NoFresh_2_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[26]), .CK(RoundFunction_C_Inst_Chi_NoFresh_2_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[34]), .CK(RoundFunction_C_Inst_Chi_NoFresh_2_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[34]), .CK(RoundFunction_C_Inst_Chi_NoFresh_2_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[2]), .CK(RoundFunction_C_Inst_Chi_NoFresh_2_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[2]), .CK(RoundFunction_C_Inst_Chi_NoFresh_2_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[10]), .CK(RoundFunction_C_Inst_Chi_NoFresh_2_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[10]), .CK(RoundFunction_C_Inst_Chi_NoFresh_2_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[1]), .Z(RESULT1[162]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[3]), .Z(RESULT2[162]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[5]), .Z(RESULT1[170]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[7]), .Z(RESULT2[170]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[9]), .Z(RESULT1[178]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[11]), .Z(RESULT2[178]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[13]), .Z(RESULT1[186]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[15]), .Z(RESULT2[186]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[17]), .Z(
        RoundFunction_TMP4_1[2]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[19]), .Z(RESULT2[194]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_3_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[19]), .CK(RoundFunction_C_Inst_Chi_NoFresh_3_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[27]), .CK(RoundFunction_C_Inst_Chi_NoFresh_3_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[27]), .CK(RoundFunction_C_Inst_Chi_NoFresh_3_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[35]), .CK(RoundFunction_C_Inst_Chi_NoFresh_3_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[35]), .CK(RoundFunction_C_Inst_Chi_NoFresh_3_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[3]), .CK(RoundFunction_C_Inst_Chi_NoFresh_3_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[3]), .CK(RoundFunction_C_Inst_Chi_NoFresh_3_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[11]), .CK(RoundFunction_C_Inst_Chi_NoFresh_3_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[11]), .CK(RoundFunction_C_Inst_Chi_NoFresh_3_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[1]), .Z(RESULT1[163]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[3]), .Z(RESULT2[163]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[5]), .Z(RESULT1[171]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[7]), .Z(RESULT2[171]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[9]), .Z(RESULT1[179]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[11]), .Z(RESULT2[179]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[13]), .Z(RESULT1[187]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[15]), .Z(RESULT2[187]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[17]), .Z(
        RoundFunction_TMP4_1[3]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[19]), .Z(RESULT2[195]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_4_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[20]), .CK(RoundFunction_C_Inst_Chi_NoFresh_4_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[28]), .CK(RoundFunction_C_Inst_Chi_NoFresh_4_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[28]), .CK(RoundFunction_C_Inst_Chi_NoFresh_4_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[4]), .CK(RoundFunction_C_Inst_Chi_NoFresh_4_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[4]), .CK(RoundFunction_C_Inst_Chi_NoFresh_4_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[12]), .CK(RoundFunction_C_Inst_Chi_NoFresh_4_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[1]), .Z(RESULT1[164]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[3]), .Z(RESULT2[164]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[5]), .Z(RESULT1[172]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[7]), .Z(RESULT2[172]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[9]), .Z(RESULT1[180]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[11]), .Z(RESULT2[180]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[13]), .Z(RESULT1[188]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[15]), .Z(RESULT2[188]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[17]), .Z(
        RoundFunction_TMP4_1[4]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[19]), .Z(RESULT2[196]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_5_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[21]), .CK(RoundFunction_C_Inst_Chi_NoFresh_5_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[29]), .CK(RoundFunction_C_Inst_Chi_NoFresh_5_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[29]), .CK(RoundFunction_C_Inst_Chi_NoFresh_5_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[37]), .CK(RoundFunction_C_Inst_Chi_NoFresh_5_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[37]), .CK(RoundFunction_C_Inst_Chi_NoFresh_5_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[5]), .CK(RoundFunction_C_Inst_Chi_NoFresh_5_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[5]), .CK(RoundFunction_C_Inst_Chi_NoFresh_5_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[13]), .CK(RoundFunction_C_Inst_Chi_NoFresh_5_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[13]), .CK(RoundFunction_C_Inst_Chi_NoFresh_5_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[1]), .Z(RESULT1[165]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[3]), .Z(RESULT2[165]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[5]), .Z(RESULT1[173]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[7]), .Z(RESULT2[173]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[9]), .Z(RESULT1[181]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[11]), .Z(RESULT2[181]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[13]), .Z(RESULT1[189]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[15]), .Z(RESULT2[189]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[17]), .Z(
        RoundFunction_TMP4_1[5]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[19]), .Z(RESULT2[197]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_6_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[22]), .CK(RoundFunction_C_Inst_Chi_NoFresh_6_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[22]), .CK(RoundFunction_C_Inst_Chi_NoFresh_6_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[30]), .CK(RoundFunction_C_Inst_Chi_NoFresh_6_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[30]), .CK(RoundFunction_C_Inst_Chi_NoFresh_6_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[38]), .CK(RoundFunction_C_Inst_Chi_NoFresh_6_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[38]), .CK(RoundFunction_C_Inst_Chi_NoFresh_6_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[6]), .CK(RoundFunction_C_Inst_Chi_NoFresh_6_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[6]), .CK(RoundFunction_C_Inst_Chi_NoFresh_6_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[14]), .CK(RoundFunction_C_Inst_Chi_NoFresh_6_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[1]), .Z(RESULT1[166]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[3]), .Z(RESULT2[166]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[5]), .Z(RESULT1[174]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[7]), .Z(RESULT2[174]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[9]), .Z(RESULT1[182]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[11]), .Z(RESULT2[182]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[13]), .Z(RESULT1[190]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[15]), .Z(RESULT2[190]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[17]), .Z(
        RoundFunction_TMP4_1[6]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[19]), .Z(RESULT2[198]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_7_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[23]), .CK(RoundFunction_C_Inst_Chi_NoFresh_7_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[23]), .CK(RoundFunction_C_Inst_Chi_NoFresh_7_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[31]), .CK(RoundFunction_C_Inst_Chi_NoFresh_7_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[31]), .CK(RoundFunction_C_Inst_Chi_NoFresh_7_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[39]), .CK(RoundFunction_C_Inst_Chi_NoFresh_7_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[39]), .CK(RoundFunction_C_Inst_Chi_NoFresh_7_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[7]), .CK(RoundFunction_C_Inst_Chi_NoFresh_7_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[15]), .CK(RoundFunction_C_Inst_Chi_NoFresh_7_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[15]), .CK(RoundFunction_C_Inst_Chi_NoFresh_7_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[1]), .Z(RESULT1[167]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[3]), .Z(RESULT2[167]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[5]), .Z(RESULT1[175]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[7]), .Z(RESULT2[175]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[9]), .Z(RESULT1[183]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[11]), .Z(RESULT2[183]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[13]), .Z(RESULT1[191]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[15]), .Z(RESULT2[191]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[17]), .Z(
        RoundFunction_TMP4_1[7]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[19]), .Z(RESULT2[199]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_8_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[56]), .CK(RoundFunction_C_Inst_Chi_NoFresh_8_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[56]), .CK(RoundFunction_C_Inst_Chi_NoFresh_8_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[64]), .CK(RoundFunction_C_Inst_Chi_NoFresh_8_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[64]), .CK(RoundFunction_C_Inst_Chi_NoFresh_8_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[72]), .CK(RoundFunction_C_Inst_Chi_NoFresh_8_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[72]), .CK(RoundFunction_C_Inst_Chi_NoFresh_8_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[40]), .CK(RoundFunction_C_Inst_Chi_NoFresh_8_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[40]), .CK(RoundFunction_C_Inst_Chi_NoFresh_8_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[48]), .CK(RoundFunction_C_Inst_Chi_NoFresh_8_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[48]), .CK(RoundFunction_C_Inst_Chi_NoFresh_8_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[1]), .Z(RESULT1[120]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[3]), .Z(RESULT2[120]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[5]), .Z(RESULT1[128]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[7]), .Z(RESULT2[128]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[9]), .Z(RESULT1[136]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[11]), .Z(RESULT2[136]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[13]), .Z(RESULT1[144]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[15]), .Z(RESULT2[144]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[17]), .Z(RESULT1[152]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[19]), .Z(RESULT2[152]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_9_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[57]), .CK(RoundFunction_C_Inst_Chi_NoFresh_9_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[57]), .CK(RoundFunction_C_Inst_Chi_NoFresh_9_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[65]), .CK(RoundFunction_C_Inst_Chi_NoFresh_9_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[65]), .CK(RoundFunction_C_Inst_Chi_NoFresh_9_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[73]), .CK(RoundFunction_C_Inst_Chi_NoFresh_9_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[73]), .CK(RoundFunction_C_Inst_Chi_NoFresh_9_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[41]), .CK(RoundFunction_C_Inst_Chi_NoFresh_9_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[41]), .CK(RoundFunction_C_Inst_Chi_NoFresh_9_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[49]), .CK(RoundFunction_C_Inst_Chi_NoFresh_9_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[49]), .CK(RoundFunction_C_Inst_Chi_NoFresh_9_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[1]), .Z(RESULT1[121]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[3]), .Z(RESULT2[121]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[5]), .Z(RESULT1[129]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[7]), .Z(RESULT2[129]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[9]), .Z(RESULT1[137]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[11]), .Z(RESULT2[137]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[13]), .Z(RESULT1[145]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[15]), .Z(RESULT2[145]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[17]), .Z(RESULT1[153]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[19]), .Z(RESULT2[153]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_10_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[58]), .CK(RoundFunction_C_Inst_Chi_NoFresh_10_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[58]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[66]), .CK(RoundFunction_C_Inst_Chi_NoFresh_10_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[66]), .CK(RoundFunction_C_Inst_Chi_NoFresh_10_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[74]), .CK(RoundFunction_C_Inst_Chi_NoFresh_10_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[74]), .CK(RoundFunction_C_Inst_Chi_NoFresh_10_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[42]), .CK(RoundFunction_C_Inst_Chi_NoFresh_10_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[42]), .CK(RoundFunction_C_Inst_Chi_NoFresh_10_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[50]), .CK(RoundFunction_C_Inst_Chi_NoFresh_10_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[50]), .CK(RoundFunction_C_Inst_Chi_NoFresh_10_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[1]), .Z(RESULT1[122]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[3]), .Z(RESULT2[122]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[5]), .Z(RESULT1[130]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[7]), .Z(RESULT2[130]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[9]), .Z(RESULT1[138]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[11]), .Z(RESULT2[138]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[13]), .Z(RESULT1[146]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[15]), .Z(RESULT2[146]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[17]), .Z(RESULT1[154]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[19]), .Z(RESULT2[154]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_11_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[59]), .CK(RoundFunction_C_Inst_Chi_NoFresh_11_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[59]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[67]), .CK(RoundFunction_C_Inst_Chi_NoFresh_11_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[67]), .CK(RoundFunction_C_Inst_Chi_NoFresh_11_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[75]), .CK(RoundFunction_C_Inst_Chi_NoFresh_11_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[75]), .CK(RoundFunction_C_Inst_Chi_NoFresh_11_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[43]), .CK(RoundFunction_C_Inst_Chi_NoFresh_11_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[43]), .CK(RoundFunction_C_Inst_Chi_NoFresh_11_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[51]), .CK(RoundFunction_C_Inst_Chi_NoFresh_11_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[51]), .CK(RoundFunction_C_Inst_Chi_NoFresh_11_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[1]), .Z(RESULT1[123]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[3]), .Z(RESULT2[123]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[5]), .Z(RESULT1[131]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[7]), .Z(RESULT2[131]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[9]), .Z(RESULT1[139]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[11]), .Z(RESULT2[139]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[13]), .Z(RESULT1[147]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[15]), .Z(RESULT2[147]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[17]), .Z(RESULT1[155]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[19]), .Z(RESULT2[155]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_12_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[60]), .CK(RoundFunction_C_Inst_Chi_NoFresh_12_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[60]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[68]), .CK(RoundFunction_C_Inst_Chi_NoFresh_12_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[68]), .CK(RoundFunction_C_Inst_Chi_NoFresh_12_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[76]), .CK(RoundFunction_C_Inst_Chi_NoFresh_12_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[76]), .CK(RoundFunction_C_Inst_Chi_NoFresh_12_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[44]), .CK(RoundFunction_C_Inst_Chi_NoFresh_12_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[44]), .CK(RoundFunction_C_Inst_Chi_NoFresh_12_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[52]), .CK(RoundFunction_C_Inst_Chi_NoFresh_12_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[52]), .CK(RoundFunction_C_Inst_Chi_NoFresh_12_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[1]), .Z(RESULT1[124]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[3]), .Z(RESULT2[124]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[5]), .Z(RESULT1[132]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[7]), .Z(RESULT2[132]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[9]), .Z(RESULT1[140]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[11]), .Z(RESULT2[140]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[13]), .Z(RESULT1[148]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[15]), .Z(RESULT2[148]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[17]), .Z(RESULT1[156]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[19]), .Z(RESULT2[156]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_13_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[61]), .CK(RoundFunction_C_Inst_Chi_NoFresh_13_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[61]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[69]), .CK(RoundFunction_C_Inst_Chi_NoFresh_13_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[69]), .CK(RoundFunction_C_Inst_Chi_NoFresh_13_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[77]), .CK(RoundFunction_C_Inst_Chi_NoFresh_13_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[77]), .CK(RoundFunction_C_Inst_Chi_NoFresh_13_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[45]), .CK(RoundFunction_C_Inst_Chi_NoFresh_13_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[45]), .CK(RoundFunction_C_Inst_Chi_NoFresh_13_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[53]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[53]), .CK(RoundFunction_C_Inst_Chi_NoFresh_13_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[1]), .Z(RESULT1[125]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[3]), .Z(RESULT2[125]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[5]), .Z(RESULT1[133]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[7]), .Z(RESULT2[133]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[9]), .Z(RESULT1[141]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[11]), .Z(RESULT2[141]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[13]), .Z(RESULT1[149]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[15]), .Z(RESULT2[149]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[17]), .Z(RESULT1[157]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[19]), .Z(RESULT2[157]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_14_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[62]), .CK(RoundFunction_C_Inst_Chi_NoFresh_14_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[62]), .CK(RoundFunction_C_Inst_Chi_NoFresh_14_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[70]), .CK(RoundFunction_C_Inst_Chi_NoFresh_14_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[70]), .CK(RoundFunction_C_Inst_Chi_NoFresh_14_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[78]), .CK(RoundFunction_C_Inst_Chi_NoFresh_14_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[78]), .CK(RoundFunction_C_Inst_Chi_NoFresh_14_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[46]), .CK(RoundFunction_C_Inst_Chi_NoFresh_14_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[46]), .CK(RoundFunction_C_Inst_Chi_NoFresh_14_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[54]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[54]), .CK(RoundFunction_C_Inst_Chi_NoFresh_14_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[1]), .Z(RESULT1[126]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[3]), .Z(RESULT2[126]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[5]), .Z(RESULT1[134]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[7]), .Z(RESULT2[134]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[9]), .Z(RESULT1[142]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[11]), .Z(RESULT2[142]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[13]), .Z(RESULT1[150]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[15]), .Z(RESULT2[150]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[17]), .Z(RESULT1[158]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[19]), .Z(RESULT2[158]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_15_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[63]), .CK(RoundFunction_C_Inst_Chi_NoFresh_15_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[63]), .CK(RoundFunction_C_Inst_Chi_NoFresh_15_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[71]), .CK(RoundFunction_C_Inst_Chi_NoFresh_15_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[71]), .CK(RoundFunction_C_Inst_Chi_NoFresh_15_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[79]), .CK(RoundFunction_C_Inst_Chi_NoFresh_15_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[79]), .CK(RoundFunction_C_Inst_Chi_NoFresh_15_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[47]), .CK(RoundFunction_C_Inst_Chi_NoFresh_15_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[47]), .CK(RoundFunction_C_Inst_Chi_NoFresh_15_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[55]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[55]), .CK(RoundFunction_C_Inst_Chi_NoFresh_15_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[1]), .Z(RESULT1[127]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[3]), .Z(RESULT2[127]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[5]), .Z(RESULT1[135]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[7]), .Z(RESULT2[135]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[9]), .Z(RESULT1[143]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[11]), .Z(RESULT2[143]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[13]), .Z(RESULT1[151]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[15]), .Z(RESULT2[151]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[17]), .Z(RESULT1[159]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[19]), .Z(RESULT2[159]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[96]), .CK(RoundFunction_C_Inst_Chi_NoFresh_16_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[96]), .CK(RoundFunction_C_Inst_Chi_NoFresh_16_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[104]), .CK(RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[104]), .CK(RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[112]), .CK(RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[112]), .CK(RoundFunction_C_Inst_Chi_NoFresh_16_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[80]), .CK(RoundFunction_C_Inst_Chi_NoFresh_16_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[80]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[88]), .CK(RoundFunction_C_Inst_Chi_NoFresh_16_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[88]), .CK(RoundFunction_C_Inst_Chi_NoFresh_16_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[1]), .Z(RESULT1[80]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[3]), .Z(RESULT2[80]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[5]), .Z(RESULT1[88]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[7]), .Z(RESULT2[88]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[9]), .Z(RESULT1[96]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[11]), .Z(RESULT2[96]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[13]), .Z(RESULT1[104]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[15]), .Z(RESULT2[104]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[17]), .Z(RESULT1[112]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[19]), .Z(RESULT2[112]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[97]), .CK(RoundFunction_C_Inst_Chi_NoFresh_17_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[97]), .CK(RoundFunction_C_Inst_Chi_NoFresh_17_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[105]), .CK(RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[105]), .CK(RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[113]), .CK(RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[113]), .CK(RoundFunction_C_Inst_Chi_NoFresh_17_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[81]), .CK(RoundFunction_C_Inst_Chi_NoFresh_17_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[81]), .CK(RoundFunction_C_Inst_Chi_NoFresh_17_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[89]), .CK(RoundFunction_C_Inst_Chi_NoFresh_17_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[89]), .CK(RoundFunction_C_Inst_Chi_NoFresh_17_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[1]), .Z(RESULT1[81]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[3]), .Z(RESULT2[81]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[5]), .Z(RESULT1[89]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[7]), .Z(RESULT2[89]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[9]), .Z(RESULT1[97]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[11]), .Z(RESULT2[97]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[13]), .Z(RESULT1[105]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[15]), .Z(RESULT2[105]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[17]), .Z(RESULT1[113]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[19]), .Z(RESULT2[113]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[98]), .CK(RoundFunction_C_Inst_Chi_NoFresh_18_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[98]), .CK(RoundFunction_C_Inst_Chi_NoFresh_18_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[106]), .CK(RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[106]), .CK(RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[114]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[114]), .CK(RoundFunction_C_Inst_Chi_NoFresh_18_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[82]), .CK(RoundFunction_C_Inst_Chi_NoFresh_18_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[82]), .CK(RoundFunction_C_Inst_Chi_NoFresh_18_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[90]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[90]), .CK(RoundFunction_C_Inst_Chi_NoFresh_18_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[1]), .Z(RESULT1[82]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[3]), .Z(RESULT2[82]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[5]), .Z(RESULT1[90]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[7]), .Z(RESULT2[90]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[9]), .Z(RESULT1[98]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[11]), .Z(RESULT2[98]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[13]), .Z(RESULT1[106]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[15]), .Z(RESULT2[106]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[17]), .Z(RESULT1[114]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[19]), .Z(RESULT2[114]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[99]), .CK(RoundFunction_C_Inst_Chi_NoFresh_19_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[99]), .CK(RoundFunction_C_Inst_Chi_NoFresh_19_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[107]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[107]), .CK(RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[115]), .CK(RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[115]), .CK(RoundFunction_C_Inst_Chi_NoFresh_19_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[83]), .CK(RoundFunction_C_Inst_Chi_NoFresh_19_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[83]), .CK(RoundFunction_C_Inst_Chi_NoFresh_19_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[91]), .CK(RoundFunction_C_Inst_Chi_NoFresh_19_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[91]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[1]), .Z(RESULT1[83]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[3]), .Z(RESULT2[83]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[5]), .Z(RESULT1[91]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[7]), .Z(RESULT2[91]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[9]), .Z(RESULT1[99]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[11]), .Z(RESULT2[99]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[13]), .Z(RESULT1[107]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[15]), .Z(RESULT2[107]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[17]), .Z(RESULT1[115]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[19]), .Z(RESULT2[115]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[100]), .CK(RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[100]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[108]), .CK(RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[108]), .CK(RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[116]), .CK(RoundFunction_C_Inst_Chi_NoFresh_20_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[116]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[84]), .CK(RoundFunction_C_Inst_Chi_NoFresh_20_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[84]), .CK(RoundFunction_C_Inst_Chi_NoFresh_20_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[92]), .CK(RoundFunction_C_Inst_Chi_NoFresh_20_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[92]), .CK(RoundFunction_C_Inst_Chi_NoFresh_20_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[1]), .Z(RESULT1[84]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[3]), .Z(RESULT2[84]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[5]), .Z(RESULT1[92]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[7]), .Z(RESULT2[92]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[9]), .Z(RESULT1[100]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[11]), .Z(RESULT2[100]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[13]), .Z(RESULT1[108]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[15]), .Z(RESULT2[108]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[17]), .Z(RESULT1[116]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[19]), .Z(RESULT2[116]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[101]), .CK(RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[101]), .CK(RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[109]), .CK(RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[109]), .CK(RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[117]), .CK(RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[117]), .CK(RoundFunction_C_Inst_Chi_NoFresh_21_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[85]), .CK(RoundFunction_C_Inst_Chi_NoFresh_21_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[85]), .CK(RoundFunction_C_Inst_Chi_NoFresh_21_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[93]), .CK(RoundFunction_C_Inst_Chi_NoFresh_21_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[93]), .CK(RoundFunction_C_Inst_Chi_NoFresh_21_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[1]), .Z(RESULT1[85]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[3]), .Z(RESULT2[85]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[5]), .Z(RESULT1[93]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[7]), .Z(RESULT2[93]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[9]), .Z(RESULT1[101]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[11]), .Z(RESULT2[101]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[13]), .Z(RESULT1[109]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[15]), .Z(RESULT2[109]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[17]), .Z(RESULT1[117]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[19]), .Z(RESULT2[117]) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[102]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[102]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[110]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[110]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[118]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[118]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[86]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[86]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[94]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[94]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[1]), .Z(RESULT1[86]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[3]), .Z(RESULT2[86]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[5]), .Z(RESULT1[94]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[7]), .Z(RESULT2[94]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[9]), .Z(RESULT1[102]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[11]), .Z(RESULT2[102]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[13]), .Z(RESULT1[110]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[15]), .Z(RESULT2[110]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[17]), .Z(RESULT1[118]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[19]), .Z(RESULT2[118]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[103]), .CK(RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[103]), .CK(RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[111]), .CK(RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[111]), .CK(RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[119]), .CK(RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[119]), .CK(RoundFunction_C_Inst_Chi_NoFresh_23_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[87]), .CK(RoundFunction_C_Inst_Chi_NoFresh_23_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[87]), .CK(RoundFunction_C_Inst_Chi_NoFresh_23_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[95]), .CK(RoundFunction_C_Inst_Chi_NoFresh_23_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[95]), .CK(RoundFunction_C_Inst_Chi_NoFresh_23_n1), 
        .Q(RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[1]), .Z(RESULT1[87]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[3]), .Z(RESULT2[87]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[5]), .Z(RESULT1[95]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[7]), .Z(RESULT2[95]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[9]), .Z(RESULT1[103]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[11]), .Z(RESULT2[103]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[13]), .Z(RESULT1[111]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[15]), .Z(RESULT2[111]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[17]), .Z(RESULT1[119]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[19]), .Z(RESULT2[119]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[136]), .CK(RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[136]), .CK(RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[144]), .CK(RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[144]), .CK(RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[152]), .CK(RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[152]), .CK(RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[120]), .CK(RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[120]), .CK(RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[128]), .CK(RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[128]), .CK(RoundFunction_C_Inst_Chi_NoFresh_24_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[1]), .Z(RESULT1[40]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[3]), .Z(RESULT2[40]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[5]), .Z(RESULT1[48]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[7]), .Z(RESULT2[48]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[9]), .Z(RESULT1[56]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[11]), .Z(RESULT2[56]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[13]), .Z(RESULT1[64]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[15]), .Z(RESULT2[64]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[17]), .Z(RESULT1[72]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[19]), .Z(RESULT2[72]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[137]), .CK(RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[137]), .CK(RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[145]), .CK(RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[145]), .CK(RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[153]), .CK(RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[153]), .CK(RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[121]), .CK(RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[121]), .CK(RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[129]), .CK(RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[129]), .CK(RoundFunction_C_Inst_Chi_NoFresh_25_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[1]), .Z(RESULT1[41]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[3]), .Z(RESULT2[41]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[5]), .Z(RESULT1[49]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[7]), .Z(RESULT2[49]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[9]), .Z(RESULT1[57]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[11]), .Z(RESULT2[57]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[13]), .Z(RESULT1[65]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[15]), .Z(RESULT2[65]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[17]), .Z(RESULT1[73]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[19]), .Z(RESULT2[73]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[138]), .CK(RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[138]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[146]), .CK(RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[146]), .CK(RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[154]), .CK(RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[154]), .CK(RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[122]), .CK(RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[122]), .CK(RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[130]), .CK(RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[130]), .CK(RoundFunction_C_Inst_Chi_NoFresh_26_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[1]), .Z(RESULT1[42]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[3]), .Z(RESULT2[42]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[5]), .Z(RESULT1[50]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[7]), .Z(RESULT2[50]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[9]), .Z(RESULT1[58]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[11]), .Z(RESULT2[58]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[13]), .Z(RESULT1[66]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[15]), .Z(RESULT2[66]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[17]), .Z(RESULT1[74]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[19]), .Z(RESULT2[74]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[139]), .CK(RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[139]), .CK(RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[147]), .CK(RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[147]), .CK(RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[155]), .CK(RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[155]), .CK(RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[123]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[123]), .CK(RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[131]), .CK(RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[131]), .CK(RoundFunction_C_Inst_Chi_NoFresh_27_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[1]), .Z(RESULT1[43]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[3]), .Z(RESULT2[43]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[5]), .Z(RESULT1[51]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[7]), .Z(RESULT2[51]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[9]), .Z(RESULT1[59]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[11]), .Z(RESULT2[59]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[13]), .Z(RESULT1[67]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[15]), .Z(RESULT2[67]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[17]), .Z(RESULT1[75]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[19]), .Z(RESULT2[75]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[140]), .CK(RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[140]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[148]), .CK(RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[148]), .CK(RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[156]), .CK(RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[156]), .CK(RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[124]), .CK(RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[124]), .CK(RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[132]), .CK(RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[132]), .CK(RoundFunction_C_Inst_Chi_NoFresh_28_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[1]), .Z(RESULT1[44]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[3]), .Z(RESULT2[44]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[5]), .Z(RESULT1[52]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[7]), .Z(RESULT2[52]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[9]), .Z(RESULT1[60]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[11]), .Z(RESULT2[60]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[13]), .Z(RESULT1[68]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[15]), .Z(RESULT2[68]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[17]), .Z(RESULT1[76]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[19]), .Z(RESULT2[76]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[141]), .CK(RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[141]), .CK(RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[149]), .CK(RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[149]), .CK(RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[157]), .CK(RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[157]), .CK(RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[125]), .CK(RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[125]), .CK(RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[133]), .CK(RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[133]), .CK(RoundFunction_C_Inst_Chi_NoFresh_29_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[1]), .Z(RESULT1[45]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[3]), .Z(RESULT2[45]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[5]), .Z(RESULT1[53]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[7]), .Z(RESULT2[53]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[9]), .Z(RESULT1[61]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[11]), .Z(RESULT2[61]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[13]), .Z(RESULT1[69]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[15]), .Z(RESULT2[69]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[17]), .Z(RESULT1[77]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[19]), .Z(RESULT2[77]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[142]), .CK(RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[142]), .CK(RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[150]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[150]), .CK(RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[158]), .CK(RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[158]), .CK(RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[126]), .CK(RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[126]), .CK(RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[134]), .CK(RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[134]), .CK(RoundFunction_C_Inst_Chi_NoFresh_30_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[1]), .Z(RESULT1[46]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[3]), .Z(RESULT2[46]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[5]), .Z(RESULT1[54]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[7]), .Z(RESULT2[54]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[9]), .Z(RESULT1[62]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[11]), .Z(RESULT2[62]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[13]), .Z(RESULT1[70]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[15]), .Z(RESULT2[70]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[17]), .Z(RESULT1[78]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[19]), .Z(RESULT2[78]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[143]), .CK(RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[143]), .CK(RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[151]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[151]), .CK(RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[159]), .CK(RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[159]), .CK(RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[127]), .CK(RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[127]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[135]), .CK(RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[135]), .CK(RoundFunction_C_Inst_Chi_NoFresh_31_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[1]), .Z(RESULT1[47]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[3]), .Z(RESULT2[47]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[5]), .Z(RESULT1[55]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[7]), .Z(RESULT2[55]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[9]), .Z(RESULT1[63]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[11]), .Z(RESULT2[63]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[13]), .Z(RESULT1[71]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[15]), .Z(RESULT2[71]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[17]), .Z(RESULT1[79]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[19]), .Z(RESULT2[79]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[176]), .CK(RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[176]), .CK(RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[184]), .CK(RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[184]), .CK(RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[192]), .CK(RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[192]), .CK(RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[160]), .CK(RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[160]), .CK(RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[168]), .CK(RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[168]), .CK(RoundFunction_C_Inst_Chi_NoFresh_32_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[1]), .Z(RESULT1[0]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[3]), .Z(RESULT2[0]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[5]), .Z(RESULT1[8]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[7]), .Z(RESULT2[8]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[9]), .Z(RESULT1[16]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[11]), .Z(RESULT2[16]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[13]), .Z(RESULT1[24]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[15]), .Z(RESULT2[24]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[17]), .Z(RESULT1[32]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[19]), .Z(RESULT2[32]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[177]), .CK(RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[177]), .CK(RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[185]), .CK(RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[185]), .CK(RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[193]), .CK(RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[193]), .CK(RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[161]), .CK(RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[161]), .CK(RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[169]), .CK(RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[169]), .CK(RoundFunction_C_Inst_Chi_NoFresh_33_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[1]), .Z(RESULT1[1]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[3]), .Z(RESULT2[1]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[5]), .Z(RESULT1[9]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[7]), .Z(RESULT2[9]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[9]), .Z(RESULT1[17]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[11]), .Z(RESULT2[17]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[13]), .Z(RESULT1[25]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[15]), .Z(RESULT2[25]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[17]), .Z(RESULT1[33]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[19]), .Z(RESULT2[33]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[178]), .CK(RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[178]), .CK(RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[186]), .CK(RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[186]), .CK(RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[194]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[194]), .CK(RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[162]), .CK(RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[162]), .CK(RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[170]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[170]), .CK(RoundFunction_C_Inst_Chi_NoFresh_34_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[1]), .Z(RESULT1[2]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[3]), .Z(RESULT2[2]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[5]), .Z(RESULT1[10]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[7]), .Z(RESULT2[10]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[9]), .Z(RESULT1[18]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[11]), .Z(RESULT2[18]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[13]), .Z(RESULT1[26]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[15]), .Z(RESULT2[26]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[17]), .Z(RESULT1[34]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[19]), .Z(RESULT2[34]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[179]), .CK(RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[179]), .CK(RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[187]), .CK(RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[187]), .CK(RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[195]), .CK(RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[195]), .CK(RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[163]), .CK(RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[163]), .CK(RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[171]), .CK(RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[171]), .CK(RoundFunction_C_Inst_Chi_NoFresh_35_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[1]), .Z(RESULT1[3]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[3]), .Z(RESULT2[3]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[5]), .Z(RESULT1[11]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[7]), .Z(RESULT2[11]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[9]), .Z(RESULT1[19]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[11]), .Z(RESULT2[19]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[13]), .Z(RESULT1[27]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[15]), .Z(RESULT2[27]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[17]), .Z(RESULT1[35]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[19]), .Z(RESULT2[35]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[180]), .CK(RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[180]), .CK(RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[188]), .CK(RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[188]), .CK(RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[196]), .CK(RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[196]), .CK(RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[164]), .CK(RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[164]), .CK(RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[172]), .CK(RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[172]), .CK(RoundFunction_C_Inst_Chi_NoFresh_36_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[1]), .Z(RESULT1[4]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[3]), .Z(RESULT2[4]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[5]), .Z(RESULT1[12]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[7]), .Z(RESULT2[12]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[9]), .Z(RESULT1[20]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[11]), .Z(RESULT2[20]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[13]), .Z(RESULT1[28]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[15]), .Z(RESULT2[28]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[17]), .Z(RESULT1[36]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[19]), .Z(RESULT2[36]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[4]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[13]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[14]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[181]), .CK(RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[181]), .CK(RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[189]), .CK(RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[189]), .CK(RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[197]), .CK(RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[197]), .CK(RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[165]), .CK(RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[165]), .CK(RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[173]), .CK(RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[173]), .CK(RoundFunction_C_Inst_Chi_NoFresh_37_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[1]), .Z(RESULT1[5]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[3]), .Z(RESULT2[5]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[5]), .Z(RESULT1[13]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[7]), .Z(RESULT2[13]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[9]), .Z(RESULT1[21]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[11]), .Z(RESULT2[21]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[13]), .Z(RESULT1[29]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[15]), .Z(RESULT2[29]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[17]), .Z(RESULT1[37]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[19]), .Z(RESULT2[37]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[182]), .CK(RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[182]), .CK(RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[190]), .CK(RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[190]), .CK(RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[198]), .CK(RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[198]), .CK(RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[166]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[166]), .CK(RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[174]), .CK(RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[174]), .CK(RoundFunction_C_Inst_Chi_NoFresh_38_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[1]), .Z(RESULT1[6]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[3]), .Z(RESULT2[6]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[5]), .Z(RESULT1[14]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[7]), .Z(RESULT2[14]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[9]), .Z(RESULT1[22]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[11]), .Z(RESULT2[22]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[13]), .Z(RESULT1[30]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[15]), .Z(RESULT2[30]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[17]), .Z(RESULT1[38]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[19]), .Z(RESULT2[38]) );
  BUF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_U3 ( .A(CLK), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[0]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[1]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[2]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[3]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[5]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[6]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[7]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[8]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[9]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[10]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[11]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[12]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[15]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[16]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[17]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[18]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[19]), .CK(
        RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[183]), .CK(RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[183]), .CK(RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[191]), .CK(RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[191]), .CK(RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[199]), .CK(RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[199]), .CK(RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[167]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[167]), .CK(RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[175]), .CK(RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[175]), .CK(RoundFunction_C_Inst_Chi_NoFresh_39_n1), .Q(RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_1__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_2__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_2__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[2]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_2__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_2__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_2__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_2__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_2__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_3__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[3]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_5__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_5__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_6__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_6__CF_Inst_n2) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_7__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_7__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[7]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_7__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_7__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_7__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_7__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_7__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_8__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[9]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[10]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_11__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[11]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_n4), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[12]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_n3) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_n4) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_13__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_13__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[13]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_13__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_13__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_13__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_13__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_13__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_14__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[14]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[15]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_n4) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_16__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_16__CF_Inst_n2), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[16]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_16__CF_Inst_n2) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_17__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_17__CF_Inst_n2), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[17]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_17__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_17__CF_Inst_n2) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n6), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[18]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n5), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n6) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_U4 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n6), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[19]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_U3 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n4), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n5) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n4) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .Z(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n6) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[1]), .Z(RESULT1[7]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[2]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[3]), .Z(RESULT2[7]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[4]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[5]), .Z(RESULT1[15]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[7]), .Z(RESULT2[15]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[8]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[9]), .Z(RESULT1[23]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[10]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[11]), .Z(RESULT2[23]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[13]), .Z(RESULT1[31]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[14]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[15]), .Z(RESULT2[31]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[16]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[17]), .Z(RESULT1[39]) );
  XOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[19]), .Z(RESULT2[39]) );
  OAI21_X1 FSM_U70 ( .B1(FSM_n152), .B2(FSM_n151), .A(FSM_n150), .ZN(FSM_n78)
         );
  OAI22_X1 FSM_U69 ( .A1(FSM_n7), .A2(FSM_n149), .B1(FSM_n8), .B2(FSM_n150), 
        .ZN(FSM_n77) );
  OAI221_X1 FSM_U68 ( .B1(FSM_n148), .B2(FSM_n98), .C1(FSM_n147), .C2(FSM_n146), .A(FSM_n103), .ZN(FSM_n76) );
  XNOR2_X1 FSM_U67 ( .A(FSM_n145), .B(FSM_n144), .ZN(FSM_n146) );
  AOI22_X1 FSM_U66 ( .A1(FSM_n87), .A2(FSM_n100), .B1(FSM_n7), .B2(FSM_n94), 
        .ZN(FSM_n144) );
  OAI22_X1 FSM_U65 ( .A1(FSM_n98), .A2(FSM_n150), .B1(FSM_n93), .B2(FSM_n149), 
        .ZN(FSM_n75) );
  OAI22_X1 FSM_U64 ( .A1(FSM_n97), .A2(FSM_n149), .B1(FSM_n93), .B2(FSM_n150), 
        .ZN(FSM_n74) );
  OAI22_X1 FSM_U63 ( .A1(FSM_n12), .A2(FSM_n149), .B1(FSM_n150), .B2(FSM_n97), 
        .ZN(FSM_n73) );
  OAI22_X1 FSM_U62 ( .A1(FSM_n12), .A2(FSM_n150), .B1(FSM_n149), .B2(FSM_n96), 
        .ZN(FSM_n72) );
  OAI22_X1 FSM_U61 ( .A1(FSM_n94), .A2(FSM_n149), .B1(FSM_n96), .B2(FSM_n150), 
        .ZN(FSM_n71) );
  OAI22_X1 FSM_U60 ( .A1(FSM_n8), .A2(FSM_n149), .B1(FSM_n94), .B2(FSM_n150), 
        .ZN(FSM_n70) );
  NAND2_X1 FSM_U59 ( .A1(FSM_n148), .A2(FSM_n103), .ZN(FSM_n150) );
  INV_X1 FSM_U58 ( .A(FSM_n147), .ZN(FSM_n148) );
  NAND2_X1 FSM_U57 ( .A1(FSM_n103), .A2(FSM_n147), .ZN(FSM_n149) );
  NAND3_X1 FSM_U56 ( .A1(FSM_n102), .A2(FSM_n86), .A3(FSM_n85), .ZN(FSM_n147)
         );
  OAI22_X1 FSM_U55 ( .A1(RESET), .A2(FSM_n143), .B1(FSM_n142), .B2(FSM_n151), 
        .ZN(FSM_n3) );
  NAND4_X1 FSM_U54 ( .A1(FSM_n19), .A2(FSM_n85), .A3(FSM_n103), .A4(FSM_n101), 
        .ZN(FSM_n151) );
  INV_X1 FSM_U53 ( .A(DONE), .ZN(FSM_n143) );
  NOR3_X1 FSM_U52 ( .A1(FSM_n19), .A2(FSM_n86), .A3(FSM_n85), .ZN(DONE) );
  NAND4_X1 FSM_U51 ( .A1(FSM_n141), .A2(FSM_n140), .A3(FSM_n139), .A4(FSM_n138), .ZN(FSM_CONST_internal_7) );
  AOI21_X1 FSM_U50 ( .B1(FSM_n137), .B2(FSM_n6), .A(FSM_n152), .ZN(FSM_n140)
         );
  NOR2_X1 FSM_U49 ( .A1(FSM_n136), .A2(FSM_n135), .ZN(FSM_n137) );
  NAND4_X1 FSM_U48 ( .A1(FSM_n134), .A2(FSM_n133), .A3(FSM_n132), .A4(FSM_n138), .ZN(FSM_CONST_internal_3) );
  NAND3_X1 FSM_U47 ( .A1(FSM_n8), .A2(FSM_n7), .A3(FSM_n131), .ZN(FSM_n138) );
  NOR4_X1 FSM_U46 ( .A1(FSM_n12), .A2(FSM_n96), .A3(FSM_n130), .A4(FSM_n129), 
        .ZN(FSM_n131) );
  INV_X1 FSM_U45 ( .A(FSM_n128), .ZN(FSM_n132) );
  OAI211_X1 FSM_U44 ( .C1(FSM_n127), .C2(FSM_n126), .A(FSM_n141), .B(FSM_n133), 
        .ZN(FSM_CONST_internal[1]) );
  NAND4_X1 FSM_U43 ( .A1(FSM_n125), .A2(FSM_n124), .A3(FSM_n95), .A4(FSM_n98), 
        .ZN(FSM_n133) );
  NOR4_X1 FSM_U42 ( .A1(FSM_n2), .A2(FSM_n7), .A3(FSM_n99), .A4(FSM_n93), .ZN(
        FSM_n124) );
  AOI211_X1 FSM_U41 ( .C1(FSM_n123), .C2(FSM_n96), .A(FSM_n128), .B(FSM_n122), 
        .ZN(FSM_n141) );
  NOR4_X1 FSM_U40 ( .A1(FSM_n97), .A2(FSM_n121), .A3(FSM_n145), .A4(FSM_n129), 
        .ZN(FSM_n128) );
  NAND2_X1 FSM_U39 ( .A1(FSM_n98), .A2(FSM_n93), .ZN(FSM_n129) );
  OAI21_X1 FSM_U38 ( .B1(FSM_n12), .B2(FSM_n2), .A(FSM_n136), .ZN(FSM_n145) );
  AOI22_X1 FSM_U37 ( .A1(FSM_n8), .A2(FSM_n120), .B1(FSM_n119), .B2(FSM_n95), 
        .ZN(FSM_n126) );
  NOR3_X1 FSM_U36 ( .A1(FSM_n87), .A2(FSM_n93), .A3(FSM_n118), .ZN(FSM_n119)
         );
  NOR3_X1 FSM_U35 ( .A1(FSM_n9), .A2(FSM_n94), .A3(FSM_n117), .ZN(FSM_n120) );
  NAND3_X1 FSM_U34 ( .A1(FSM_n134), .A2(FSM_n139), .A3(FSM_n116), .ZN(
        FSM_CONST_internal[0]) );
  INV_X1 FSM_U33 ( .A(FSM_n115), .ZN(FSM_n116) );
  AOI211_X1 FSM_U32 ( .C1(FSM_n94), .C2(FSM_n4), .A(FSM_n95), .B(FSM_n114), 
        .ZN(FSM_n115) );
  OAI221_X1 FSM_U31 ( .B1(FSM_n93), .B2(FSM_n125), .C1(FSM_n9), .C2(FSM_n130), 
        .A(FSM_n113), .ZN(FSM_n114) );
  INV_X1 FSM_U30 ( .A(FSM_n130), .ZN(FSM_n125) );
  NAND4_X1 FSM_U29 ( .A1(FSM_n113), .A2(FSM_n112), .A3(FSM_n94), .A4(FSM_n95), 
        .ZN(FSM_n139) );
  NOR2_X1 FSM_U28 ( .A1(FSM_n97), .A2(FSM_n93), .ZN(FSM_n112) );
  NOR2_X1 FSM_U27 ( .A1(FSM_n99), .A2(FSM_n127), .ZN(FSM_n113) );
  NAND3_X1 FSM_U26 ( .A1(FSM_n6), .A2(FSM_n7), .A3(FSM_n96), .ZN(FSM_n127) );
  NOR4_X1 FSM_U25 ( .A1(FSM_n152), .A2(FSM_n122), .A3(FSM_n111), .A4(FSM_n110), 
        .ZN(FSM_n134) );
  NOR4_X1 FSM_U24 ( .A1(FSM_n12), .A2(FSM_n6), .A3(FSM_n2), .A4(FSM_n135), 
        .ZN(FSM_n110) );
  NAND4_X1 FSM_U23 ( .A1(FSM_n4), .A2(FSM_n9), .A3(FSM_n109), .A4(FSM_n100), 
        .ZN(FSM_n135) );
  NOR2_X1 FSM_U22 ( .A1(FSM_n87), .A2(FSM_n95), .ZN(FSM_n109) );
  NOR3_X1 FSM_U21 ( .A1(FSM_n136), .A2(FSM_n130), .A3(FSM_n108), .ZN(FSM_n111)
         );
  NAND4_X1 FSM_U20 ( .A1(FSM_n7), .A2(FSM_n6), .A3(FSM_n95), .A4(FSM_n93), 
        .ZN(FSM_n108) );
  NAND2_X1 FSM_U19 ( .A1(FSM_n87), .A2(FSM_n97), .ZN(FSM_n130) );
  NAND2_X1 FSM_U18 ( .A1(FSM_n12), .A2(FSM_n2), .ZN(FSM_n136) );
  AOI21_X1 FSM_U17 ( .B1(FSM_n107), .B2(FSM_n106), .A(FSM_n9), .ZN(FSM_n122)
         );
  NAND3_X1 FSM_U16 ( .A1(FSM_n6), .A2(FSM_n2), .A3(FSM_n105), .ZN(FSM_n106) );
  NAND4_X1 FSM_U15 ( .A1(FSM_n94), .A2(FSM_n100), .A3(FSM_n96), .A4(FSM_n104), 
        .ZN(FSM_n107) );
  OAI33_X1 FSM_U14 ( .A1(FSM_n6), .A2(FSM_n8), .A3(FSM_n117), .B1(FSM_n98), 
        .B2(FSM_n118), .B3(FSM_n95), .ZN(FSM_n104) );
  NAND2_X1 FSM_U13 ( .A1(FSM_n99), .A2(FSM_n97), .ZN(FSM_n118) );
  NAND2_X1 FSM_U12 ( .A1(FSM_n12), .A2(FSM_n4), .ZN(FSM_n117) );
  INV_X1 FSM_U11 ( .A(FSM_n142), .ZN(FSM_n152) );
  NAND2_X1 FSM_U10 ( .A1(FSM_n2), .A2(FSM_n123), .ZN(FSM_n142) );
  AND3_X1 FSM_U9 ( .A1(FSM_n9), .A2(FSM_n105), .A3(FSM_n98), .ZN(FSM_n123) );
  NOR3_X1 FSM_U8 ( .A1(FSM_n4), .A2(FSM_n99), .A3(FSM_n121), .ZN(FSM_n105) );
  NAND3_X1 FSM_U7 ( .A1(FSM_n8), .A2(FSM_n7), .A3(FSM_n94), .ZN(FSM_n121) );
  INV_X1 FSM_U6 ( .A(RESET), .ZN(FSM_n103) );
  AOI21_X1 FSM_U5 ( .B1(FSM_n92), .B2(FSM_n152), .A(FSM_n91), .ZN(FSM_n79) );
  NOR2_X1 FSM_U4 ( .A1(FSM_n86), .A2(FSM_n102), .ZN(FSM_n92) );
  OAI211_X1 FSM_U3 ( .C1(FSM_n19), .C2(FSM_n101), .A(FSM_n85), .B(FSM_n103), 
        .ZN(FSM_n91) );
  DFF_X1 FSM_CONST_reg_0_ ( .D(FSM_CONST_internal[0]), .CK(CLK), .Q(CONST[0]), 
        .QN() );
  DFF_X1 FSM_CONST_reg_3_ ( .D(FSM_CONST_internal_3), .CK(CLK), .Q(CONST[3]), 
        .QN() );
  DFF_X1 FSM_CONST_reg_1_ ( .D(FSM_CONST_internal[1]), .CK(CLK), .Q(CONST[1]), 
        .QN() );
  DFF_X1 FSM_CONST_reg_7_ ( .D(FSM_CONST_internal_7), .CK(CLK), .Q(CONST[7]), 
        .QN() );
  DFF_X1 FSM_STATE_reg_1_ ( .D(FSM_n78), .CK(CLK), .Q(FSM_n19), .QN(FSM_n102)
         );
  DFF_X1 FSM_LFSR_reg_6_ ( .D(FSM_n70), .CK(CLK), .Q(FSM_n95), .QN(FSM_n8) );
  DFF_X1 FSM_LFSR_reg_5_ ( .D(FSM_n71), .CK(CLK), .Q(FSM_n87), .QN(FSM_n94) );
  DFF_X1 FSM_LFSR_reg_4_ ( .D(FSM_n72), .CK(CLK), .Q(FSM_n2), .QN(FSM_n96) );
  DFF_X1 FSM_LFSR_reg_3_ ( .D(FSM_n73), .CK(CLK), .Q(FSM_n99), .QN(FSM_n12) );
  DFF_X1 FSM_LFSR_reg_2_ ( .D(FSM_n74), .CK(CLK), .Q(FSM_n4), .QN(FSM_n97) );
  DFF_X1 FSM_LFSR_reg_1_ ( .D(FSM_n75), .CK(CLK), .Q(FSM_n9), .QN(FSM_n93) );
  DFF_X1 FSM_LFSR_reg_0_ ( .D(FSM_n76), .CK(CLK), .Q(FSM_n6), .QN(FSM_n98) );
  DFF_X1 FSM_LFSR_reg_7_ ( .D(FSM_n77), .CK(CLK), .Q(FSM_n100), .QN(FSM_n7) );
  DFF_X1 FSM_STATE_reg_2_ ( .D(FSM_n3), .CK(CLK), .Q(), .QN(FSM_n85) );
  DFF_X1 FSM_STATE_reg_0_ ( .D(FSM_n79), .CK(CLK), .Q(FSM_n86), .QN(FSM_n101)
         );
endmodule

