module circuit ( clk, rst, en, enc, p0, p1, p2, p3, b_guard, c_guard, d_guard, 
        k, c0, c1, c2, c3, done );
  input [63:0] p0;
  input [63:0] p1;
  input [63:0] p2;
  input [63:0] p3;
  input [3:0] b_guard;
  input [3:0] c_guard;
  input [3:0] d_guard;
  input [127:0] k;
  output [63:0] c0;
  output [63:0] c1;
  output [63:0] c2;
  output [63:0] c3;
  input clk, rst, en, enc;
  output done;
  wire   kext_64_, start_sig, en_sig, rc_63_, rc_62_, rc_61_, rc_60_, rc_59_,
         rc_58_, rc_57_, rc_56_, rc_55_, rc_54_, rc_53_, rc_52_, rc_51_,
         rc_50_, rc_49_, rc_48_, rc_47_, rc_46_, rc_45_, rc_44_, rc_43_,
         rc_42_, rc_41_, rc_40_, rc_39_, rc_38_, rc_37_, rc_36_, rc_35_,
         rc_34_, rc_33_, rc_32_, rc_31_, rc_30_, rc_29_, rc_28_, rc_27_,
         rc_26_, rc_25_, rc_24_, rc_23_, rc_22_, rc_21_, rc_20_, rc_19_,
         rc_18_, rc_17_, rc_16_, rc_14_, rc_13_, rc_12_, rc_11_, rc_10_, rc_9_,
         rc_8_, rc_7_, rc_6_, rc_5_, rc_4_, rc_3_, rc_2_, rc_1_, rc_0_,
         inv_sig, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, mux_w_n138,
         mux_w_n137, mux_w_n136, mux_w_n135, mux_x_n266, mux_x_n265,
         mux_x_n264, mux_x_n263, mux_y_n266, mux_y_n265, mux_y_n264,
         mux_y_n263, mux_z_n266, mux_z_n265, mux_z_n264, mux_z_n263,
         reg_w_n339, reg_w_n338, reg_w_n337, reg_w_n336, reg_w_n335,
         reg_w_n334, reg_w_n333, reg_w_n332, reg_w_n331, reg_w_n330,
         reg_w_n329, reg_w_n328, reg_w_n327, reg_w_n326, reg_w_n325,
         reg_w_n324, reg_w_n323, reg_w_n322, reg_w_n321, reg_w_n320,
         reg_w_n319, reg_w_n318, reg_w_n317, reg_w_n316, reg_w_n315,
         reg_w_n314, reg_w_n313, reg_w_n312, reg_w_n311, reg_w_n310,
         reg_w_n309, reg_w_n308, reg_w_n307, reg_w_n306, reg_w_n305,
         reg_w_n304, reg_w_n303, reg_w_n302, reg_w_n301, reg_w_n300,
         reg_w_n299, reg_w_n298, reg_w_n297, reg_w_n296, reg_w_n295,
         reg_w_n294, reg_w_n293, reg_w_n292, reg_w_n291, reg_w_n290,
         reg_w_n289, reg_w_n288, reg_w_n287, reg_w_n286, reg_w_n285,
         reg_w_n284, reg_w_n283, reg_w_n282, reg_w_n281, reg_w_n280,
         reg_w_n279, reg_w_n278, reg_w_n277, reg_w_n276, reg_w_n275,
         reg_w_n274, reg_w_n273, reg_w_n272, reg_w_n271, reg_w_n270,
         reg_w_n269, reg_w_n268, reg_w_n267, reg_w_n266, reg_w_n265,
         reg_w_n264, reg_w_n263, reg_w_n262, reg_w_n261, reg_w_n260,
         reg_w_n259, reg_w_n258, reg_w_n257, reg_w_n256, reg_w_n255,
         reg_w_n254, reg_w_n253, reg_w_n252, reg_w_n251, reg_w_n250,
         reg_w_n249, reg_w_n248, reg_w_n247, reg_w_n246, reg_w_n245,
         reg_w_n244, reg_w_n243, reg_w_n242, reg_w_n241, reg_w_n240,
         reg_w_n239, reg_w_n238, reg_w_n237, reg_w_n236, reg_w_n235,
         reg_w_n234, reg_w_n233, reg_w_n232, reg_w_n231, reg_w_n230,
         reg_w_n229, reg_w_n228, reg_w_n227, reg_w_n226, reg_w_n225,
         reg_w_n224, reg_w_n223, reg_w_n222, reg_w_n221, reg_w_n220,
         reg_w_n219, reg_w_n218, reg_w_n217, reg_w_n216, reg_w_n215,
         reg_w_n214, reg_w_n213, reg_w_n212, reg_w_n211, reg_w_n210,
         reg_w_n209, reg_w_n208, reg_w_n207, reg_w_n206, reg_w_n205,
         reg_w_n204, reg_w_n203, reg_w_n202, reg_w_n195, reg_w_n194,
         reg_w_n193, reg_w_n192, reg_w_n191, reg_w_n190, reg_w_n189,
         reg_w_n188, reg_w_n187, reg_w_n186, reg_w_n185, reg_w_n184,
         reg_w_n183, reg_w_n182, reg_w_n181, reg_w_n180, reg_w_n179,
         reg_w_n178, reg_w_n177, reg_w_n176, reg_w_n175, reg_w_n174,
         reg_w_n173, reg_w_n172, reg_w_n171, reg_w_n170, reg_w_n169,
         reg_w_n168, reg_w_n167, reg_w_n166, reg_w_n165, reg_w_n164,
         reg_w_n163, reg_w_n162, reg_w_n161, reg_w_n160, reg_w_n159,
         reg_w_n158, reg_w_n157, reg_w_n156, reg_w_n155, reg_w_n154,
         reg_w_n153, reg_w_n152, reg_w_n151, reg_w_n150, reg_w_n149,
         reg_w_n148, reg_w_n147, reg_w_n146, reg_w_n145, reg_w_n144,
         reg_w_n143, reg_w_n142, reg_w_n141, reg_w_n140, reg_w_n139,
         reg_w_n138, reg_w_n137, reg_w_n136, reg_w_n135, reg_w_n134,
         reg_w_n133, reg_w_n132, reg_x_n532, reg_x_n531, reg_x_n530,
         reg_x_n529, reg_x_n528, reg_x_n527, reg_x_n526, reg_x_n525,
         reg_x_n524, reg_x_n523, reg_x_n522, reg_x_n521, reg_x_n520,
         reg_x_n519, reg_x_n518, reg_x_n517, reg_x_n516, reg_x_n515,
         reg_x_n514, reg_x_n513, reg_x_n512, reg_x_n511, reg_x_n510,
         reg_x_n509, reg_x_n508, reg_x_n507, reg_x_n506, reg_x_n505,
         reg_x_n504, reg_x_n503, reg_x_n502, reg_x_n501, reg_x_n500,
         reg_x_n499, reg_x_n498, reg_x_n497, reg_x_n496, reg_x_n495,
         reg_x_n494, reg_x_n493, reg_x_n492, reg_x_n491, reg_x_n490,
         reg_x_n489, reg_x_n488, reg_x_n487, reg_x_n486, reg_x_n485,
         reg_x_n484, reg_x_n483, reg_x_n482, reg_x_n481, reg_x_n480,
         reg_x_n479, reg_x_n478, reg_x_n477, reg_x_n476, reg_x_n475,
         reg_x_n474, reg_x_n473, reg_x_n472, reg_x_n471, reg_x_n470,
         reg_x_n469, reg_x_n468, reg_x_n467, reg_x_n466, reg_x_n465,
         reg_x_n464, reg_x_n463, reg_x_n462, reg_x_n461, reg_x_n460,
         reg_x_n459, reg_x_n458, reg_x_n457, reg_x_n456, reg_x_n455,
         reg_x_n454, reg_x_n453, reg_x_n452, reg_x_n451, reg_x_n450,
         reg_x_n449, reg_x_n448, reg_x_n447, reg_x_n446, reg_x_n445,
         reg_x_n444, reg_x_n443, reg_x_n442, reg_x_n441, reg_x_n440,
         reg_x_n439, reg_x_n438, reg_x_n437, reg_x_n436, reg_x_n435,
         reg_x_n434, reg_x_n433, reg_x_n432, reg_x_n431, reg_x_n430,
         reg_x_n429, reg_x_n428, reg_x_n427, reg_x_n426, reg_x_n425,
         reg_x_n424, reg_x_n423, reg_x_n422, reg_x_n421, reg_x_n420,
         reg_x_n419, reg_x_n418, reg_x_n417, reg_x_n416, reg_x_n415,
         reg_x_n414, reg_x_n413, reg_x_n412, reg_x_n411, reg_x_n410,
         reg_x_n409, reg_x_n408, reg_x_n407, reg_x_n406, reg_x_n405,
         reg_x_n404, reg_x_n403, reg_x_n402, reg_x_n401, reg_x_n400,
         reg_x_n399, reg_x_n398, reg_x_n397, reg_x_n396, reg_x_n395,
         reg_x_n394, reg_x_n265, reg_x_n264, reg_x_n263, reg_x_n262,
         reg_x_n261, reg_x_n260, reg_x_n259, reg_x_n258, reg_x_n257,
         reg_x_n256, reg_x_n255, reg_x_n254, reg_x_n253, reg_x_n252,
         reg_x_n251, reg_x_n250, reg_x_n249, reg_x_n248, reg_x_n247,
         reg_x_n246, reg_x_n245, reg_x_n244, reg_x_n243, reg_x_n242,
         reg_x_n241, reg_x_n240, reg_x_n239, reg_x_n238, reg_x_n237,
         reg_x_n236, reg_x_n235, reg_x_n234, reg_x_n233, reg_x_n232,
         reg_x_n231, reg_x_n230, reg_x_n229, reg_x_n228, reg_x_n227,
         reg_x_n226, reg_x_n225, reg_x_n224, reg_x_n223, reg_x_n222,
         reg_x_n221, reg_x_n220, reg_x_n219, reg_x_n218, reg_x_n217,
         reg_x_n216, reg_x_n215, reg_x_n214, reg_x_n213, reg_x_n212,
         reg_x_n211, reg_x_n210, reg_x_n209, reg_x_n208, reg_x_n207,
         reg_x_n206, reg_x_n205, reg_x_n204, reg_x_n203, reg_x_n202,
         reg_y_n532, reg_y_n531, reg_y_n530, reg_y_n529, reg_y_n528,
         reg_y_n527, reg_y_n526, reg_y_n525, reg_y_n524, reg_y_n523,
         reg_y_n522, reg_y_n521, reg_y_n520, reg_y_n519, reg_y_n518,
         reg_y_n517, reg_y_n516, reg_y_n515, reg_y_n514, reg_y_n513,
         reg_y_n512, reg_y_n511, reg_y_n510, reg_y_n509, reg_y_n508,
         reg_y_n507, reg_y_n506, reg_y_n505, reg_y_n504, reg_y_n503,
         reg_y_n502, reg_y_n501, reg_y_n500, reg_y_n499, reg_y_n498,
         reg_y_n497, reg_y_n496, reg_y_n495, reg_y_n494, reg_y_n493,
         reg_y_n492, reg_y_n491, reg_y_n490, reg_y_n489, reg_y_n488,
         reg_y_n487, reg_y_n486, reg_y_n485, reg_y_n484, reg_y_n483,
         reg_y_n482, reg_y_n481, reg_y_n480, reg_y_n479, reg_y_n478,
         reg_y_n477, reg_y_n476, reg_y_n475, reg_y_n474, reg_y_n473,
         reg_y_n472, reg_y_n471, reg_y_n470, reg_y_n469, reg_y_n468,
         reg_y_n467, reg_y_n466, reg_y_n465, reg_y_n464, reg_y_n463,
         reg_y_n462, reg_y_n461, reg_y_n460, reg_y_n459, reg_y_n458,
         reg_y_n457, reg_y_n456, reg_y_n455, reg_y_n454, reg_y_n453,
         reg_y_n452, reg_y_n451, reg_y_n450, reg_y_n449, reg_y_n448,
         reg_y_n447, reg_y_n446, reg_y_n445, reg_y_n444, reg_y_n443,
         reg_y_n442, reg_y_n441, reg_y_n440, reg_y_n439, reg_y_n438,
         reg_y_n437, reg_y_n436, reg_y_n435, reg_y_n434, reg_y_n433,
         reg_y_n432, reg_y_n431, reg_y_n430, reg_y_n429, reg_y_n428,
         reg_y_n427, reg_y_n426, reg_y_n425, reg_y_n424, reg_y_n423,
         reg_y_n422, reg_y_n421, reg_y_n420, reg_y_n419, reg_y_n418,
         reg_y_n417, reg_y_n416, reg_y_n415, reg_y_n414, reg_y_n413,
         reg_y_n412, reg_y_n411, reg_y_n410, reg_y_n409, reg_y_n408,
         reg_y_n407, reg_y_n406, reg_y_n405, reg_y_n404, reg_y_n403,
         reg_y_n402, reg_y_n401, reg_y_n400, reg_y_n399, reg_y_n398,
         reg_y_n397, reg_y_n396, reg_y_n395, reg_y_n394, reg_y_n265,
         reg_y_n264, reg_y_n263, reg_y_n262, reg_y_n261, reg_y_n260,
         reg_y_n259, reg_y_n258, reg_y_n257, reg_y_n256, reg_y_n255,
         reg_y_n254, reg_y_n253, reg_y_n252, reg_y_n251, reg_y_n250,
         reg_y_n249, reg_y_n248, reg_y_n247, reg_y_n246, reg_y_n245,
         reg_y_n244, reg_y_n243, reg_y_n242, reg_y_n241, reg_y_n240,
         reg_y_n239, reg_y_n238, reg_y_n237, reg_y_n236, reg_y_n235,
         reg_y_n234, reg_y_n233, reg_y_n232, reg_y_n231, reg_y_n230,
         reg_y_n229, reg_y_n228, reg_y_n227, reg_y_n226, reg_y_n225,
         reg_y_n224, reg_y_n223, reg_y_n222, reg_y_n221, reg_y_n220,
         reg_y_n219, reg_y_n218, reg_y_n217, reg_y_n216, reg_y_n215,
         reg_y_n214, reg_y_n213, reg_y_n212, reg_y_n211, reg_y_n210,
         reg_y_n209, reg_y_n208, reg_y_n207, reg_y_n206, reg_y_n205,
         reg_y_n204, reg_y_n203, reg_y_n202, reg_z_n532, reg_z_n531,
         reg_z_n530, reg_z_n529, reg_z_n528, reg_z_n527, reg_z_n526,
         reg_z_n525, reg_z_n524, reg_z_n523, reg_z_n522, reg_z_n521,
         reg_z_n520, reg_z_n519, reg_z_n518, reg_z_n517, reg_z_n516,
         reg_z_n515, reg_z_n514, reg_z_n513, reg_z_n512, reg_z_n511,
         reg_z_n510, reg_z_n509, reg_z_n508, reg_z_n507, reg_z_n506,
         reg_z_n505, reg_z_n504, reg_z_n503, reg_z_n502, reg_z_n501,
         reg_z_n500, reg_z_n499, reg_z_n498, reg_z_n497, reg_z_n496,
         reg_z_n495, reg_z_n494, reg_z_n493, reg_z_n492, reg_z_n491,
         reg_z_n490, reg_z_n489, reg_z_n488, reg_z_n487, reg_z_n486,
         reg_z_n485, reg_z_n484, reg_z_n483, reg_z_n482, reg_z_n481,
         reg_z_n480, reg_z_n479, reg_z_n478, reg_z_n477, reg_z_n476,
         reg_z_n475, reg_z_n474, reg_z_n473, reg_z_n472, reg_z_n471,
         reg_z_n470, reg_z_n469, reg_z_n468, reg_z_n467, reg_z_n466,
         reg_z_n465, reg_z_n464, reg_z_n463, reg_z_n462, reg_z_n461,
         reg_z_n460, reg_z_n459, reg_z_n458, reg_z_n457, reg_z_n456,
         reg_z_n455, reg_z_n454, reg_z_n453, reg_z_n452, reg_z_n451,
         reg_z_n450, reg_z_n449, reg_z_n448, reg_z_n447, reg_z_n446,
         reg_z_n445, reg_z_n444, reg_z_n443, reg_z_n442, reg_z_n441,
         reg_z_n440, reg_z_n439, reg_z_n438, reg_z_n437, reg_z_n436,
         reg_z_n435, reg_z_n434, reg_z_n433, reg_z_n432, reg_z_n431,
         reg_z_n430, reg_z_n429, reg_z_n428, reg_z_n427, reg_z_n426,
         reg_z_n425, reg_z_n424, reg_z_n423, reg_z_n422, reg_z_n421,
         reg_z_n420, reg_z_n419, reg_z_n418, reg_z_n417, reg_z_n416,
         reg_z_n415, reg_z_n414, reg_z_n413, reg_z_n412, reg_z_n411,
         reg_z_n410, reg_z_n409, reg_z_n408, reg_z_n407, reg_z_n406,
         reg_z_n405, reg_z_n404, reg_z_n403, reg_z_n402, reg_z_n401,
         reg_z_n400, reg_z_n399, reg_z_n398, reg_z_n397, reg_z_n396,
         reg_z_n395, reg_z_n394, reg_z_n265, reg_z_n264, reg_z_n263,
         reg_z_n262, reg_z_n261, reg_z_n260, reg_z_n259, reg_z_n258,
         reg_z_n257, reg_z_n256, reg_z_n255, reg_z_n254, reg_z_n253,
         reg_z_n252, reg_z_n251, reg_z_n250, reg_z_n249, reg_z_n248,
         reg_z_n247, reg_z_n246, reg_z_n245, reg_z_n244, reg_z_n243,
         reg_z_n242, reg_z_n241, reg_z_n240, reg_z_n239, reg_z_n238,
         reg_z_n237, reg_z_n236, reg_z_n235, reg_z_n234, reg_z_n233,
         reg_z_n232, reg_z_n231, reg_z_n230, reg_z_n229, reg_z_n228,
         reg_z_n227, reg_z_n226, reg_z_n225, reg_z_n224, reg_z_n223,
         reg_z_n222, reg_z_n221, reg_z_n220, reg_z_n219, reg_z_n218,
         reg_z_n217, reg_z_n216, reg_z_n215, reg_z_n214, reg_z_n213,
         reg_z_n212, reg_z_n211, reg_z_n210, reg_z_n209, reg_z_n208,
         reg_z_n207, reg_z_n206, reg_z_n205, reg_z_n204, reg_z_n203,
         reg_z_n202, reg_b_n16, reg_b_n11, reg_b_n10, reg_b_n9, reg_b_n8,
         reg_b_n7, reg_b_n6, reg_b_n5, reg_b_n4, reg_b_n3, reg_b_n2, reg_b_n15,
         reg_b_n14, reg_b_n13, reg_b_n12, reg_c_n40, reg_c_n39, reg_c_n38,
         reg_c_n37, reg_c_n36, reg_c_n35, reg_c_n34, reg_c_n33, reg_c_n32,
         reg_c_n31, reg_c_n30, reg_c_n19, reg_c_n18, reg_c_n17, reg_c_n16,
         reg_d_n40, reg_d_n39, reg_d_n38, reg_d_n37, reg_d_n36, reg_d_n35,
         reg_d_n34, reg_d_n33, reg_d_n32, reg_d_n31, reg_d_n30, reg_d_n19,
         reg_d_n18, reg_d_n17, reg_d_n16, cntrl_inst_n222, cntrl_inst_n221,
         cntrl_inst_n220, cntrl_inst_n219, cntrl_inst_n218, cntrl_inst_n217,
         cntrl_inst_n216, cntrl_inst_n215, cntrl_inst_n214, cntrl_inst_n213,
         cntrl_inst_n212, cntrl_inst_n211, cntrl_inst_n210, cntrl_inst_n209,
         cntrl_inst_n208, cntrl_inst_n207, cntrl_inst_n206, cntrl_inst_n205,
         cntrl_inst_n204, cntrl_inst_n203, cntrl_inst_n202, cntrl_inst_n201,
         cntrl_inst_n200, cntrl_inst_n199, cntrl_inst_n198, cntrl_inst_n197,
         cntrl_inst_n196, cntrl_inst_n195, cntrl_inst_n194, cntrl_inst_n193,
         cntrl_inst_n192, cntrl_inst_n191, cntrl_inst_n190, cntrl_inst_n189,
         cntrl_inst_n188, cntrl_inst_n187, cntrl_inst_n186, cntrl_inst_n185,
         cntrl_inst_n184, cntrl_inst_n183, cntrl_inst_n182, cntrl_inst_n181,
         cntrl_inst_n180, cntrl_inst_n179, cntrl_inst_n178, cntrl_inst_n177,
         cntrl_inst_n176, cntrl_inst_n175, cntrl_inst_n174, cntrl_inst_n173,
         cntrl_inst_n172, cntrl_inst_n171, cntrl_inst_n170, cntrl_inst_n169,
         cntrl_inst_n168, cntrl_inst_n167, cntrl_inst_n166, cntrl_inst_n165,
         cntrl_inst_n164, cntrl_inst_n163, cntrl_inst_n162, cntrl_inst_n161,
         cntrl_inst_n160, cntrl_inst_n159, cntrl_inst_n158, cntrl_inst_n157,
         cntrl_inst_n156, cntrl_inst_n155, cntrl_inst_n154, cntrl_inst_n153,
         cntrl_inst_n152, cntrl_inst_n151, cntrl_inst_n150, cntrl_inst_n149,
         cntrl_inst_n148, cntrl_inst_n147, cntrl_inst_n146, cntrl_inst_n145,
         cntrl_inst_n144, cntrl_inst_n143, cntrl_inst_n142, cntrl_inst_n141,
         cntrl_inst_n140, cntrl_inst_n139, cntrl_inst_n138, cntrl_inst_n137,
         cntrl_inst_n136, cntrl_inst_n135, cntrl_inst_n134, cntrl_inst_n133,
         cntrl_inst_n132, cntrl_inst_n131, cntrl_inst_n130, cntrl_inst_n129,
         cntrl_inst_n128, cntrl_inst_n127, cntrl_inst_n126, cntrl_inst_n125,
         cntrl_inst_n124, cntrl_inst_n123, cntrl_inst_n122, cntrl_inst_n121,
         cntrl_inst_n120, cntrl_inst_n119, cntrl_inst_n118, cntrl_inst_n117,
         cntrl_inst_n116, cntrl_inst_n115, cntrl_inst_n114, cntrl_inst_n113,
         cntrl_inst_n112, cntrl_inst_n111, cntrl_inst_n110, cntrl_inst_n109,
         cntrl_inst_n108, cntrl_inst_n102, cntrl_inst_n100, cntrl_inst_n99,
         cntrl_inst_n98, round_inst_n70, round_inst_n69, round_inst_n68,
         round_inst_n67, round_inst_n66, round_inst_n65, round_inst_n64,
         round_inst_n63, round_inst_n62, round_inst_n61, round_inst_n60,
         round_inst_n59, round_inst_n58, round_inst_n57, round_inst_n56,
         round_inst_n55, round_inst_n54, round_inst_n53, round_inst_n52,
         round_inst_n51, round_inst_n50, round_inst_n49, round_inst_n48,
         round_inst_n47, round_inst_n46, round_inst_n45, round_inst_n44,
         round_inst_n43, round_inst_n42, round_inst_n41, round_inst_n40,
         round_inst_n39, round_inst_n38, round_inst_n37, round_inst_n36,
         round_inst_n35, round_inst_n34, round_inst_n33, round_inst_n32,
         round_inst_n31, round_inst_n30, round_inst_n29, round_inst_n28,
         round_inst_n27, round_inst_n26, round_inst_n25, round_inst_n24,
         round_inst_n23, round_inst_n22, round_inst_n21, round_inst_n20,
         round_inst_n19, round_inst_n18, round_inst_n17, round_inst_n16,
         round_inst_n15, round_inst_n14, round_inst_n13, round_inst_n12,
         round_inst_n11, round_inst_n10, round_inst_n9, round_inst_n8,
         round_inst_n7, round_inst_n6, round_inst_n72, round_inst_A_0__aw_n3,
         round_inst_A_0__ax_n1, round_inst_A_0__ay_n3, round_inst_A_0__az_n3,
         round_inst_A_1__aw_n5, round_inst_A_1__ax_n3, round_inst_A_1__ay_n3,
         round_inst_A_1__az_n3, round_inst_A_2__aw_n5, round_inst_A_2__ax_n3,
         round_inst_A_2__ay_n3, round_inst_A_2__az_n3, round_inst_A_3__aw_n5,
         round_inst_A_3__ax_n3, round_inst_A_3__ay_n3, round_inst_A_3__az_n3,
         round_inst_A_4__aw_n5, round_inst_A_4__ax_n3, round_inst_A_4__ay_n3,
         round_inst_A_4__az_n3, round_inst_A_5__aw_n5, round_inst_A_5__ax_n3,
         round_inst_A_5__ay_n3, round_inst_A_5__az_n3, round_inst_A_6__aw_n5,
         round_inst_A_6__ax_n3, round_inst_A_6__ay_n3, round_inst_A_6__az_n3,
         round_inst_A_7__aw_n5, round_inst_A_7__ax_n3, round_inst_A_7__ay_n3,
         round_inst_A_7__az_n3, round_inst_A_8__aw_n5, round_inst_A_8__ax_n3,
         round_inst_A_8__ay_n3, round_inst_A_8__az_n3, round_inst_A_9__aw_n5,
         round_inst_A_9__ax_n3, round_inst_A_9__ay_n3, round_inst_A_9__az_n3,
         round_inst_A_10__aw_n5, round_inst_A_10__ax_n3,
         round_inst_A_10__ay_n3, round_inst_A_10__az_n3,
         round_inst_A_11__aw_n5, round_inst_A_11__ax_n3,
         round_inst_A_11__ay_n3, round_inst_A_11__az_n3,
         round_inst_A_12__aw_n5, round_inst_A_12__ax_n3,
         round_inst_A_12__ay_n3, round_inst_A_12__az_n3,
         round_inst_A_13__aw_n5, round_inst_A_13__ax_n3,
         round_inst_A_13__ay_n3, round_inst_A_13__az_n3,
         round_inst_A_14__aw_n5, round_inst_A_14__ax_n3,
         round_inst_A_14__ay_n3, round_inst_A_14__az_n3,
         round_inst_A_15__aw_n5, round_inst_A_15__ax_n3,
         round_inst_A_15__ay_n3, round_inst_A_15__az_n3,
         round_inst_mux_inv_w_n266, round_inst_mux_inv_w_n265,
         round_inst_mux_inv_w_n264, round_inst_mux_inv_w_n263,
         round_inst_mux_inv_x_n266, round_inst_mux_inv_x_n265,
         round_inst_mux_inv_x_n264, round_inst_mux_inv_x_n263,
         round_inst_mux_inv_y_n268, round_inst_mux_inv_y_n267,
         round_inst_mux_inv_y_n266, round_inst_mux_inv_y_n265,
         round_inst_mux_inv_y_n263, round_inst_mux_inv_y_n269,
         round_inst_mux_inv_z_n267, round_inst_mux_inv_z_n266,
         round_inst_mux_inv_z_n265, round_inst_mux_inv_z_n264,
         round_inst_mux_inv_z_n263, round_inst_sbox_inst0_com_w_inst_n160,
         round_inst_sbox_inst0_com_w_inst_n159,
         round_inst_sbox_inst0_com_w_inst_n158,
         round_inst_sbox_inst0_com_w_inst_n157,
         round_inst_sbox_inst0_com_w_inst_n156,
         round_inst_sbox_inst0_com_w_inst_n155,
         round_inst_sbox_inst0_com_w_inst_n154,
         round_inst_sbox_inst0_com_w_inst_n153,
         round_inst_sbox_inst0_com_w_inst_n152,
         round_inst_sbox_inst0_com_w_inst_n151,
         round_inst_sbox_inst0_com_w_inst_n150,
         round_inst_sbox_inst0_com_w_inst_n149,
         round_inst_sbox_inst0_com_w_inst_n148,
         round_inst_sbox_inst0_com_w_inst_n147,
         round_inst_sbox_inst0_com_w_inst_n146,
         round_inst_sbox_inst0_com_w_inst_n145,
         round_inst_sbox_inst0_com_w_inst_n144,
         round_inst_sbox_inst0_com_w_inst_n143,
         round_inst_sbox_inst0_com_w_inst_n142,
         round_inst_sbox_inst0_com_w_inst_n141,
         round_inst_sbox_inst0_com_w_inst_n140,
         round_inst_sbox_inst0_com_w_inst_n139,
         round_inst_sbox_inst0_com_w_inst_n138,
         round_inst_sbox_inst0_com_w_inst_n137,
         round_inst_sbox_inst0_com_w_inst_n136,
         round_inst_sbox_inst0_com_w_inst_n135,
         round_inst_sbox_inst0_com_w_inst_n134,
         round_inst_sbox_inst0_com_w_inst_n133,
         round_inst_sbox_inst0_com_w_inst_n132,
         round_inst_sbox_inst0_com_w_inst_n131,
         round_inst_sbox_inst0_com_w_inst_n130,
         round_inst_sbox_inst0_com_w_inst_n129,
         round_inst_sbox_inst0_com_w_inst_n128,
         round_inst_sbox_inst0_com_w_inst_n127,
         round_inst_sbox_inst0_com_w_inst_n126,
         round_inst_sbox_inst0_com_w_inst_n125,
         round_inst_sbox_inst0_com_w_inst_n124,
         round_inst_sbox_inst0_com_w_inst_n123,
         round_inst_sbox_inst0_com_w_inst_n122,
         round_inst_sbox_inst0_com_w_inst_n121,
         round_inst_sbox_inst0_com_w_inst_n120,
         round_inst_sbox_inst0_com_w_inst_n119,
         round_inst_sbox_inst0_com_w_inst_n118,
         round_inst_sbox_inst0_com_w_inst_n117,
         round_inst_sbox_inst0_com_w_inst_n116,
         round_inst_sbox_inst0_com_w_inst_n115,
         round_inst_sbox_inst0_com_w_inst_n114,
         round_inst_sbox_inst0_com_w_inst_n113,
         round_inst_sbox_inst0_com_w_inst_n112,
         round_inst_sbox_inst0_com_w_inst_n111,
         round_inst_sbox_inst0_com_w_inst_n110,
         round_inst_sbox_inst0_com_w_inst_n109,
         round_inst_sbox_inst0_com_w_inst_n108,
         round_inst_sbox_inst0_com_w_inst_n107,
         round_inst_sbox_inst0_com_w_inst_n106,
         round_inst_sbox_inst0_com_w_inst_n105,
         round_inst_sbox_inst0_com_w_inst_n104,
         round_inst_sbox_inst0_com_w_inst_n103,
         round_inst_sbox_inst0_com_w_inst_n102,
         round_inst_sbox_inst0_com_w_inst_n101,
         round_inst_sbox_inst0_com_w_inst_n100,
         round_inst_sbox_inst0_com_w_inst_n99,
         round_inst_sbox_inst0_com_w_inst_n98,
         round_inst_sbox_inst0_com_w_inst_n97,
         round_inst_sbox_inst0_com_w_inst_n96,
         round_inst_sbox_inst0_com_w_inst_n95,
         round_inst_sbox_inst0_com_w_inst_n94,
         round_inst_sbox_inst0_com_w_inst_n93,
         round_inst_sbox_inst0_com_w_inst_n92,
         round_inst_sbox_inst0_com_w_inst_n91,
         round_inst_sbox_inst0_com_w_inst_n90,
         round_inst_sbox_inst0_com_w_inst_n89,
         round_inst_sbox_inst0_com_w_inst_n88,
         round_inst_sbox_inst0_com_w_inst_n87,
         round_inst_sbox_inst0_com_w_inst_n86,
         round_inst_sbox_inst0_com_w_inst_n85,
         round_inst_sbox_inst0_com_w_inst_n84,
         round_inst_sbox_inst0_com_w_inst_n83,
         round_inst_sbox_inst0_com_w_inst_n82,
         round_inst_sbox_inst0_com_w_inst_n81,
         round_inst_sbox_inst0_com_w_inst_n80,
         round_inst_sbox_inst0_com_w_inst_n79,
         round_inst_sbox_inst0_com_w_inst_n78,
         round_inst_sbox_inst0_com_w_inst_n77,
         round_inst_sbox_inst0_com_w_inst_n76,
         round_inst_sbox_inst0_com_w_inst_n75,
         round_inst_sbox_inst0_com_w_inst_n74,
         round_inst_sbox_inst0_com_w_inst_n73,
         round_inst_sbox_inst0_com_w_inst_n72,
         round_inst_sbox_inst0_com_w_inst_n71,
         round_inst_sbox_inst0_com_w_inst_n70,
         round_inst_sbox_inst0_com_w_inst_n69,
         round_inst_sbox_inst0_com_w_inst_n68,
         round_inst_sbox_inst0_com_w_inst_n67,
         round_inst_sbox_inst0_com_w_inst_n66,
         round_inst_sbox_inst0_com_w_inst_n65,
         round_inst_sbox_inst0_com_w_inst_n64,
         round_inst_sbox_inst0_com_w_inst_n63,
         round_inst_sbox_inst0_com_w_inst_n62,
         round_inst_sbox_inst0_com_w_inst_n61,
         round_inst_sbox_inst0_com_w_inst_n60,
         round_inst_sbox_inst0_com_w_inst_n59,
         round_inst_sbox_inst0_com_w_inst_n58,
         round_inst_sbox_inst0_com_w_inst_n57,
         round_inst_sbox_inst0_com_w_inst_n56,
         round_inst_sbox_inst0_com_w_inst_n55,
         round_inst_sbox_inst0_com_w_inst_n54,
         round_inst_sbox_inst0_com_w_inst_n53,
         round_inst_sbox_inst0_com_w_inst_n52,
         round_inst_sbox_inst0_com_w_inst_n51,
         round_inst_sbox_inst0_com_w_inst_n50,
         round_inst_sbox_inst0_com_w_inst_n49,
         round_inst_sbox_inst0_com_w_inst_n48,
         round_inst_sbox_inst0_com_w_inst_n47,
         round_inst_sbox_inst0_com_w_inst_n46,
         round_inst_sbox_inst0_com_w_inst_n45,
         round_inst_sbox_inst0_com_w_inst_n44,
         round_inst_sbox_inst0_com_w_inst_n43,
         round_inst_sbox_inst0_com_w_inst_n42,
         round_inst_sbox_inst0_com_w_inst_n41,
         round_inst_sbox_inst0_com_w_inst_n40,
         round_inst_sbox_inst0_com_w_inst_n39,
         round_inst_sbox_inst0_com_w_inst_n38,
         round_inst_sbox_inst0_com_w_inst_n37,
         round_inst_sbox_inst0_com_w_inst_n36,
         round_inst_sbox_inst0_com_w_inst_n35,
         round_inst_sbox_inst0_com_w_inst_n34,
         round_inst_sbox_inst0_com_w_inst_n33,
         round_inst_sbox_inst0_com_w_inst_n32,
         round_inst_sbox_inst0_com_w_inst_n31,
         round_inst_sbox_inst0_com_w_inst_n30,
         round_inst_sbox_inst0_com_w_inst_n29,
         round_inst_sbox_inst0_com_w_inst_n28,
         round_inst_sbox_inst0_com_w_inst_n27,
         round_inst_sbox_inst0_com_w_inst_n26,
         round_inst_sbox_inst0_com_w_inst_n25,
         round_inst_sbox_inst0_com_w_inst_n24,
         round_inst_sbox_inst0_com_w_inst_n23,
         round_inst_sbox_inst0_com_w_inst_n22,
         round_inst_sbox_inst0_com_w_inst_n21,
         round_inst_sbox_inst0_com_w_inst_n20,
         round_inst_sbox_inst0_com_w_inst_n19,
         round_inst_sbox_inst0_com_w_inst_n18,
         round_inst_sbox_inst0_com_w_inst_n17,
         round_inst_sbox_inst0_com_w_inst_n16,
         round_inst_sbox_inst0_com_x_inst_n299,
         round_inst_sbox_inst0_com_x_inst_n298,
         round_inst_sbox_inst0_com_x_inst_n297,
         round_inst_sbox_inst0_com_x_inst_n296,
         round_inst_sbox_inst0_com_x_inst_n295,
         round_inst_sbox_inst0_com_x_inst_n294,
         round_inst_sbox_inst0_com_x_inst_n293,
         round_inst_sbox_inst0_com_x_inst_n292,
         round_inst_sbox_inst0_com_x_inst_n291,
         round_inst_sbox_inst0_com_x_inst_n290,
         round_inst_sbox_inst0_com_x_inst_n289,
         round_inst_sbox_inst0_com_x_inst_n288,
         round_inst_sbox_inst0_com_x_inst_n287,
         round_inst_sbox_inst0_com_x_inst_n286,
         round_inst_sbox_inst0_com_x_inst_n285,
         round_inst_sbox_inst0_com_x_inst_n284,
         round_inst_sbox_inst0_com_x_inst_n283,
         round_inst_sbox_inst0_com_x_inst_n282,
         round_inst_sbox_inst0_com_x_inst_n281,
         round_inst_sbox_inst0_com_x_inst_n280,
         round_inst_sbox_inst0_com_x_inst_n279,
         round_inst_sbox_inst0_com_x_inst_n278,
         round_inst_sbox_inst0_com_x_inst_n277,
         round_inst_sbox_inst0_com_x_inst_n276,
         round_inst_sbox_inst0_com_x_inst_n275,
         round_inst_sbox_inst0_com_x_inst_n274,
         round_inst_sbox_inst0_com_x_inst_n273,
         round_inst_sbox_inst0_com_x_inst_n272,
         round_inst_sbox_inst0_com_x_inst_n271,
         round_inst_sbox_inst0_com_x_inst_n270,
         round_inst_sbox_inst0_com_x_inst_n269,
         round_inst_sbox_inst0_com_x_inst_n268,
         round_inst_sbox_inst0_com_x_inst_n267,
         round_inst_sbox_inst0_com_x_inst_n266,
         round_inst_sbox_inst0_com_x_inst_n265,
         round_inst_sbox_inst0_com_x_inst_n264,
         round_inst_sbox_inst0_com_x_inst_n263,
         round_inst_sbox_inst0_com_x_inst_n262,
         round_inst_sbox_inst0_com_x_inst_n261,
         round_inst_sbox_inst0_com_x_inst_n260,
         round_inst_sbox_inst0_com_x_inst_n259,
         round_inst_sbox_inst0_com_x_inst_n258,
         round_inst_sbox_inst0_com_x_inst_n257,
         round_inst_sbox_inst0_com_x_inst_n256,
         round_inst_sbox_inst0_com_x_inst_n255,
         round_inst_sbox_inst0_com_x_inst_n254,
         round_inst_sbox_inst0_com_x_inst_n253,
         round_inst_sbox_inst0_com_x_inst_n252,
         round_inst_sbox_inst0_com_x_inst_n251,
         round_inst_sbox_inst0_com_x_inst_n250,
         round_inst_sbox_inst0_com_x_inst_n249,
         round_inst_sbox_inst0_com_x_inst_n248,
         round_inst_sbox_inst0_com_x_inst_n247,
         round_inst_sbox_inst0_com_x_inst_n246,
         round_inst_sbox_inst0_com_x_inst_n245,
         round_inst_sbox_inst0_com_x_inst_n244,
         round_inst_sbox_inst0_com_x_inst_n243,
         round_inst_sbox_inst0_com_x_inst_n242,
         round_inst_sbox_inst0_com_x_inst_n241,
         round_inst_sbox_inst0_com_x_inst_n240,
         round_inst_sbox_inst0_com_x_inst_n239,
         round_inst_sbox_inst0_com_x_inst_n238,
         round_inst_sbox_inst0_com_x_inst_n237,
         round_inst_sbox_inst0_com_x_inst_n236,
         round_inst_sbox_inst0_com_x_inst_n235,
         round_inst_sbox_inst0_com_x_inst_n234,
         round_inst_sbox_inst0_com_x_inst_n233,
         round_inst_sbox_inst0_com_x_inst_n232,
         round_inst_sbox_inst0_com_x_inst_n231,
         round_inst_sbox_inst0_com_x_inst_n230,
         round_inst_sbox_inst0_com_x_inst_n229,
         round_inst_sbox_inst0_com_x_inst_n228,
         round_inst_sbox_inst0_com_x_inst_n227,
         round_inst_sbox_inst0_com_x_inst_n226,
         round_inst_sbox_inst0_com_x_inst_n225,
         round_inst_sbox_inst0_com_x_inst_n224,
         round_inst_sbox_inst0_com_x_inst_n223,
         round_inst_sbox_inst0_com_x_inst_n222,
         round_inst_sbox_inst0_com_x_inst_n221,
         round_inst_sbox_inst0_com_x_inst_n220,
         round_inst_sbox_inst0_com_x_inst_n219,
         round_inst_sbox_inst0_com_x_inst_n218,
         round_inst_sbox_inst0_com_x_inst_n217,
         round_inst_sbox_inst0_com_x_inst_n216,
         round_inst_sbox_inst0_com_x_inst_n215,
         round_inst_sbox_inst0_com_x_inst_n214,
         round_inst_sbox_inst0_com_x_inst_n213,
         round_inst_sbox_inst0_com_x_inst_n212,
         round_inst_sbox_inst0_com_x_inst_n211,
         round_inst_sbox_inst0_com_x_inst_n210,
         round_inst_sbox_inst0_com_x_inst_n209,
         round_inst_sbox_inst0_com_x_inst_n208,
         round_inst_sbox_inst0_com_x_inst_n207,
         round_inst_sbox_inst0_com_x_inst_n206,
         round_inst_sbox_inst0_com_x_inst_n205,
         round_inst_sbox_inst0_com_x_inst_n204,
         round_inst_sbox_inst0_com_x_inst_n203,
         round_inst_sbox_inst0_com_x_inst_n202,
         round_inst_sbox_inst0_com_x_inst_n201,
         round_inst_sbox_inst0_com_x_inst_n200,
         round_inst_sbox_inst0_com_x_inst_n199,
         round_inst_sbox_inst0_com_x_inst_n198,
         round_inst_sbox_inst0_com_x_inst_n197,
         round_inst_sbox_inst0_com_x_inst_n196,
         round_inst_sbox_inst0_com_x_inst_n195,
         round_inst_sbox_inst0_com_x_inst_n194,
         round_inst_sbox_inst0_com_x_inst_n193,
         round_inst_sbox_inst0_com_x_inst_n192,
         round_inst_sbox_inst0_com_x_inst_n191,
         round_inst_sbox_inst0_com_x_inst_n190,
         round_inst_sbox_inst0_com_x_inst_n189,
         round_inst_sbox_inst0_com_x_inst_n188,
         round_inst_sbox_inst0_com_x_inst_n187,
         round_inst_sbox_inst0_com_x_inst_n186,
         round_inst_sbox_inst0_com_x_inst_n185,
         round_inst_sbox_inst0_com_x_inst_n184,
         round_inst_sbox_inst0_com_x_inst_n183,
         round_inst_sbox_inst0_com_x_inst_n182,
         round_inst_sbox_inst0_com_x_inst_n181,
         round_inst_sbox_inst0_com_x_inst_n180,
         round_inst_sbox_inst0_com_x_inst_n179,
         round_inst_sbox_inst0_com_x_inst_n178,
         round_inst_sbox_inst0_com_x_inst_n177,
         round_inst_sbox_inst0_com_x_inst_n176,
         round_inst_sbox_inst0_com_x_inst_n175,
         round_inst_sbox_inst0_com_x_inst_n174,
         round_inst_sbox_inst0_com_x_inst_n173,
         round_inst_sbox_inst0_com_x_inst_n172,
         round_inst_sbox_inst0_com_x_inst_n171,
         round_inst_sbox_inst0_com_x_inst_n170,
         round_inst_sbox_inst0_com_x_inst_n169,
         round_inst_sbox_inst0_com_x_inst_n168,
         round_inst_sbox_inst0_com_x_inst_n167,
         round_inst_sbox_inst0_com_x_inst_n166,
         round_inst_sbox_inst0_com_x_inst_n165,
         round_inst_sbox_inst0_com_x_inst_n164,
         round_inst_sbox_inst0_com_x_inst_n163,
         round_inst_sbox_inst0_com_x_inst_n162,
         round_inst_sbox_inst0_com_x_inst_n161,
         round_inst_sbox_inst0_com_x_inst_n160,
         round_inst_sbox_inst0_com_x_inst_n159,
         round_inst_sbox_inst0_com_y_inst_n155,
         round_inst_sbox_inst0_com_y_inst_n154,
         round_inst_sbox_inst0_com_y_inst_n153,
         round_inst_sbox_inst0_com_y_inst_n152,
         round_inst_sbox_inst0_com_y_inst_n151,
         round_inst_sbox_inst0_com_y_inst_n150,
         round_inst_sbox_inst0_com_y_inst_n149,
         round_inst_sbox_inst0_com_y_inst_n148,
         round_inst_sbox_inst0_com_y_inst_n147,
         round_inst_sbox_inst0_com_y_inst_n146,
         round_inst_sbox_inst0_com_y_inst_n145,
         round_inst_sbox_inst0_com_y_inst_n144,
         round_inst_sbox_inst0_com_y_inst_n143,
         round_inst_sbox_inst0_com_y_inst_n142,
         round_inst_sbox_inst0_com_y_inst_n141,
         round_inst_sbox_inst0_com_y_inst_n140,
         round_inst_sbox_inst0_com_y_inst_n139,
         round_inst_sbox_inst0_com_y_inst_n138,
         round_inst_sbox_inst0_com_y_inst_n137,
         round_inst_sbox_inst0_com_y_inst_n136,
         round_inst_sbox_inst0_com_y_inst_n135,
         round_inst_sbox_inst0_com_y_inst_n134,
         round_inst_sbox_inst0_com_y_inst_n133,
         round_inst_sbox_inst0_com_y_inst_n132,
         round_inst_sbox_inst0_com_y_inst_n131,
         round_inst_sbox_inst0_com_y_inst_n130,
         round_inst_sbox_inst0_com_y_inst_n129,
         round_inst_sbox_inst0_com_y_inst_n128,
         round_inst_sbox_inst0_com_y_inst_n127,
         round_inst_sbox_inst0_com_y_inst_n126,
         round_inst_sbox_inst0_com_y_inst_n125,
         round_inst_sbox_inst0_com_y_inst_n124,
         round_inst_sbox_inst0_com_y_inst_n123,
         round_inst_sbox_inst0_com_y_inst_n122,
         round_inst_sbox_inst0_com_y_inst_n121,
         round_inst_sbox_inst0_com_y_inst_n120,
         round_inst_sbox_inst0_com_y_inst_n119,
         round_inst_sbox_inst0_com_y_inst_n118,
         round_inst_sbox_inst0_com_y_inst_n117,
         round_inst_sbox_inst0_com_y_inst_n116,
         round_inst_sbox_inst0_com_y_inst_n115,
         round_inst_sbox_inst0_com_y_inst_n114,
         round_inst_sbox_inst0_com_y_inst_n113,
         round_inst_sbox_inst0_com_y_inst_n112,
         round_inst_sbox_inst0_com_y_inst_n111,
         round_inst_sbox_inst0_com_y_inst_n110,
         round_inst_sbox_inst0_com_y_inst_n109,
         round_inst_sbox_inst0_com_y_inst_n108,
         round_inst_sbox_inst0_com_y_inst_n107,
         round_inst_sbox_inst0_com_y_inst_n106,
         round_inst_sbox_inst0_com_y_inst_n105,
         round_inst_sbox_inst0_com_y_inst_n104,
         round_inst_sbox_inst0_com_y_inst_n103,
         round_inst_sbox_inst0_com_y_inst_n102,
         round_inst_sbox_inst0_com_y_inst_n101,
         round_inst_sbox_inst0_com_y_inst_n100,
         round_inst_sbox_inst0_com_y_inst_n99,
         round_inst_sbox_inst0_com_y_inst_n98,
         round_inst_sbox_inst0_com_y_inst_n97,
         round_inst_sbox_inst0_com_y_inst_n96,
         round_inst_sbox_inst0_com_y_inst_n95,
         round_inst_sbox_inst0_com_y_inst_n94,
         round_inst_sbox_inst0_com_y_inst_n93,
         round_inst_sbox_inst0_com_y_inst_n92,
         round_inst_sbox_inst0_com_y_inst_n91,
         round_inst_sbox_inst0_com_y_inst_n90,
         round_inst_sbox_inst0_com_y_inst_n89,
         round_inst_sbox_inst0_com_y_inst_n88,
         round_inst_sbox_inst0_com_y_inst_n87,
         round_inst_sbox_inst0_com_y_inst_n86,
         round_inst_sbox_inst0_com_y_inst_n85,
         round_inst_sbox_inst0_com_y_inst_n84,
         round_inst_sbox_inst0_com_y_inst_n83,
         round_inst_sbox_inst0_com_y_inst_n82,
         round_inst_sbox_inst0_com_y_inst_n81,
         round_inst_sbox_inst0_com_y_inst_n80,
         round_inst_sbox_inst0_com_y_inst_n79,
         round_inst_sbox_inst0_com_y_inst_n78,
         round_inst_sbox_inst0_com_y_inst_n77,
         round_inst_sbox_inst0_com_y_inst_n76,
         round_inst_sbox_inst0_com_y_inst_n75,
         round_inst_sbox_inst0_com_y_inst_n74,
         round_inst_sbox_inst0_com_y_inst_n73,
         round_inst_sbox_inst0_com_y_inst_n72,
         round_inst_sbox_inst0_com_y_inst_n71,
         round_inst_sbox_inst0_com_y_inst_n70,
         round_inst_sbox_inst0_com_y_inst_n69,
         round_inst_sbox_inst0_com_y_inst_n68,
         round_inst_sbox_inst0_com_y_inst_n67,
         round_inst_sbox_inst0_com_y_inst_n66,
         round_inst_sbox_inst0_com_y_inst_n65,
         round_inst_sbox_inst0_com_y_inst_n64,
         round_inst_sbox_inst0_com_y_inst_n63,
         round_inst_sbox_inst0_com_y_inst_n62,
         round_inst_sbox_inst0_com_y_inst_n61,
         round_inst_sbox_inst0_com_y_inst_n60,
         round_inst_sbox_inst0_com_y_inst_n59,
         round_inst_sbox_inst0_com_y_inst_n58,
         round_inst_sbox_inst0_com_y_inst_n57,
         round_inst_sbox_inst0_com_y_inst_n56,
         round_inst_sbox_inst0_com_y_inst_n55,
         round_inst_sbox_inst0_com_y_inst_n54,
         round_inst_sbox_inst0_com_y_inst_n53,
         round_inst_sbox_inst0_com_y_inst_n52,
         round_inst_sbox_inst0_com_y_inst_n51,
         round_inst_sbox_inst0_com_y_inst_n50,
         round_inst_sbox_inst0_com_y_inst_n49,
         round_inst_sbox_inst0_com_y_inst_n48,
         round_inst_sbox_inst0_com_y_inst_n47,
         round_inst_sbox_inst0_com_y_inst_n46,
         round_inst_sbox_inst0_com_y_inst_n45,
         round_inst_sbox_inst0_com_y_inst_n44,
         round_inst_sbox_inst0_com_y_inst_n43,
         round_inst_sbox_inst0_com_y_inst_n42,
         round_inst_sbox_inst0_com_y_inst_n41,
         round_inst_sbox_inst0_com_y_inst_n40,
         round_inst_sbox_inst0_com_y_inst_n39,
         round_inst_sbox_inst0_com_y_inst_n38,
         round_inst_sbox_inst0_com_y_inst_n37,
         round_inst_sbox_inst0_com_y_inst_n36,
         round_inst_sbox_inst0_com_y_inst_n35,
         round_inst_sbox_inst0_com_y_inst_n34,
         round_inst_sbox_inst0_com_y_inst_n33,
         round_inst_sbox_inst0_com_y_inst_n32,
         round_inst_sbox_inst0_com_y_inst_n31,
         round_inst_sbox_inst0_com_y_inst_n30,
         round_inst_sbox_inst0_com_y_inst_n29,
         round_inst_sbox_inst0_com_y_inst_n28,
         round_inst_sbox_inst0_com_y_inst_n27,
         round_inst_sbox_inst0_com_y_inst_n26,
         round_inst_sbox_inst0_com_y_inst_n25,
         round_inst_sbox_inst0_com_y_inst_n24,
         round_inst_sbox_inst0_com_y_inst_n23,
         round_inst_sbox_inst0_com_y_inst_n22,
         round_inst_sbox_inst0_com_y_inst_n21,
         round_inst_sbox_inst0_com_y_inst_n20,
         round_inst_sbox_inst0_com_y_inst_n19,
         round_inst_sbox_inst0_com_y_inst_n18,
         round_inst_sbox_inst0_com_y_inst_n17,
         round_inst_sbox_inst0_com_y_inst_n16,
         round_inst_sbox_inst0_com_z_inst_n274,
         round_inst_sbox_inst0_com_z_inst_n273,
         round_inst_sbox_inst0_com_z_inst_n272,
         round_inst_sbox_inst0_com_z_inst_n271,
         round_inst_sbox_inst0_com_z_inst_n270,
         round_inst_sbox_inst0_com_z_inst_n269,
         round_inst_sbox_inst0_com_z_inst_n268,
         round_inst_sbox_inst0_com_z_inst_n267,
         round_inst_sbox_inst0_com_z_inst_n266,
         round_inst_sbox_inst0_com_z_inst_n265,
         round_inst_sbox_inst0_com_z_inst_n264,
         round_inst_sbox_inst0_com_z_inst_n263,
         round_inst_sbox_inst0_com_z_inst_n262,
         round_inst_sbox_inst0_com_z_inst_n261,
         round_inst_sbox_inst0_com_z_inst_n260,
         round_inst_sbox_inst0_com_z_inst_n259,
         round_inst_sbox_inst0_com_z_inst_n258,
         round_inst_sbox_inst0_com_z_inst_n257,
         round_inst_sbox_inst0_com_z_inst_n256,
         round_inst_sbox_inst0_com_z_inst_n255,
         round_inst_sbox_inst0_com_z_inst_n254,
         round_inst_sbox_inst0_com_z_inst_n253,
         round_inst_sbox_inst0_com_z_inst_n252,
         round_inst_sbox_inst0_com_z_inst_n251,
         round_inst_sbox_inst0_com_z_inst_n250,
         round_inst_sbox_inst0_com_z_inst_n249,
         round_inst_sbox_inst0_com_z_inst_n248,
         round_inst_sbox_inst0_com_z_inst_n247,
         round_inst_sbox_inst0_com_z_inst_n246,
         round_inst_sbox_inst0_com_z_inst_n245,
         round_inst_sbox_inst0_com_z_inst_n244,
         round_inst_sbox_inst0_com_z_inst_n243,
         round_inst_sbox_inst0_com_z_inst_n242,
         round_inst_sbox_inst0_com_z_inst_n241,
         round_inst_sbox_inst0_com_z_inst_n240,
         round_inst_sbox_inst0_com_z_inst_n239,
         round_inst_sbox_inst0_com_z_inst_n238,
         round_inst_sbox_inst0_com_z_inst_n237,
         round_inst_sbox_inst0_com_z_inst_n236,
         round_inst_sbox_inst0_com_z_inst_n235,
         round_inst_sbox_inst0_com_z_inst_n234,
         round_inst_sbox_inst0_com_z_inst_n233,
         round_inst_sbox_inst0_com_z_inst_n232,
         round_inst_sbox_inst0_com_z_inst_n231,
         round_inst_sbox_inst0_com_z_inst_n230,
         round_inst_sbox_inst0_com_z_inst_n229,
         round_inst_sbox_inst0_com_z_inst_n228,
         round_inst_sbox_inst0_com_z_inst_n227,
         round_inst_sbox_inst0_com_z_inst_n226,
         round_inst_sbox_inst0_com_z_inst_n225,
         round_inst_sbox_inst0_com_z_inst_n224,
         round_inst_sbox_inst0_com_z_inst_n223,
         round_inst_sbox_inst0_com_z_inst_n222,
         round_inst_sbox_inst0_com_z_inst_n221,
         round_inst_sbox_inst0_com_z_inst_n220,
         round_inst_sbox_inst0_com_z_inst_n219,
         round_inst_sbox_inst0_com_z_inst_n218,
         round_inst_sbox_inst0_com_z_inst_n217,
         round_inst_sbox_inst0_com_z_inst_n216,
         round_inst_sbox_inst0_com_z_inst_n215,
         round_inst_sbox_inst0_com_z_inst_n214,
         round_inst_sbox_inst0_com_z_inst_n213,
         round_inst_sbox_inst0_com_z_inst_n212,
         round_inst_sbox_inst0_com_z_inst_n211,
         round_inst_sbox_inst0_com_z_inst_n210,
         round_inst_sbox_inst0_com_z_inst_n209,
         round_inst_sbox_inst0_com_z_inst_n208,
         round_inst_sbox_inst0_com_z_inst_n207,
         round_inst_sbox_inst0_com_z_inst_n206,
         round_inst_sbox_inst0_com_z_inst_n205,
         round_inst_sbox_inst0_com_z_inst_n204,
         round_inst_sbox_inst0_com_z_inst_n203,
         round_inst_sbox_inst0_com_z_inst_n202,
         round_inst_sbox_inst0_com_z_inst_n201,
         round_inst_sbox_inst0_com_z_inst_n200,
         round_inst_sbox_inst0_com_z_inst_n199,
         round_inst_sbox_inst0_com_z_inst_n198,
         round_inst_sbox_inst0_com_z_inst_n197,
         round_inst_sbox_inst0_com_z_inst_n196,
         round_inst_sbox_inst0_com_z_inst_n195,
         round_inst_sbox_inst0_com_z_inst_n194,
         round_inst_sbox_inst0_com_z_inst_n193,
         round_inst_sbox_inst0_com_z_inst_n192,
         round_inst_sbox_inst0_com_z_inst_n191,
         round_inst_sbox_inst0_com_z_inst_n190,
         round_inst_sbox_inst0_com_z_inst_n189,
         round_inst_sbox_inst0_com_z_inst_n188,
         round_inst_sbox_inst0_com_z_inst_n187,
         round_inst_sbox_inst0_com_z_inst_n186,
         round_inst_sbox_inst0_com_z_inst_n185,
         round_inst_sbox_inst0_com_z_inst_n184,
         round_inst_sbox_inst0_com_z_inst_n183,
         round_inst_sbox_inst0_com_z_inst_n182,
         round_inst_sbox_inst0_com_z_inst_n181,
         round_inst_sbox_inst0_com_z_inst_n180,
         round_inst_sbox_inst0_com_z_inst_n179,
         round_inst_sbox_inst0_com_z_inst_n178,
         round_inst_sbox_inst0_com_z_inst_n177,
         round_inst_sbox_inst0_com_z_inst_n176,
         round_inst_sbox_inst0_com_z_inst_n175,
         round_inst_sbox_inst0_com_z_inst_n174,
         round_inst_sbox_inst0_com_z_inst_n173,
         round_inst_sbox_inst0_com_z_inst_n172,
         round_inst_sbox_inst0_com_z_inst_n171,
         round_inst_sbox_inst0_com_z_inst_n170,
         round_inst_sbox_inst0_com_z_inst_n169,
         round_inst_sbox_inst0_com_z_inst_n168,
         round_inst_sbox_inst0_com_z_inst_n167,
         round_inst_sbox_inst0_com_z_inst_n166,
         round_inst_sbox_inst0_com_z_inst_n165,
         round_inst_sbox_inst0_com_z_inst_n164,
         round_inst_sbox_inst0_com_z_inst_n163,
         round_inst_sbox_inst0_com_z_inst_n162,
         round_inst_sbox_inst0_com_z_inst_n161,
         round_inst_sbox_inst0_com_z_inst_n160,
         round_inst_sbox_inst0_com_z_inst_n159,
         round_inst_sbox_inst0_com_z_inst_n158,
         round_inst_sbox_inst0_com_z_inst_n157,
         round_inst_sbox_inst0_com_z_inst_n156,
         round_inst_sbox_inst0_com_z_inst_n155,
         round_inst_sbox_inst0_com_z_inst_n154,
         round_inst_sbox_inst0_com_z_inst_n153,
         round_inst_sbox_inst0_com_z_inst_n152,
         round_inst_sbox_inst0_com_z_inst_n151,
         round_inst_sbox_inst0_com_z_inst_n150,
         round_inst_sbox_inst0_com_z_inst_n149,
         round_inst_sbox_inst0_com_z_inst_n148,
         round_inst_sbox_inst0_com_z_inst_n147,
         round_inst_sbox_inst0_com_z_inst_n146,
         round_inst_sbox_inst0_com_z_inst_n145,
         round_inst_sbox_inst0_com_z_inst_n144, round_inst_S_1__sbox_inst_n2,
         round_inst_S_1__sbox_inst_n1,
         round_inst_S_1__sbox_inst_com_w_inst_n538,
         round_inst_S_1__sbox_inst_com_w_inst_n537,
         round_inst_S_1__sbox_inst_com_w_inst_n536,
         round_inst_S_1__sbox_inst_com_w_inst_n535,
         round_inst_S_1__sbox_inst_com_w_inst_n534,
         round_inst_S_1__sbox_inst_com_w_inst_n533,
         round_inst_S_1__sbox_inst_com_w_inst_n532,
         round_inst_S_1__sbox_inst_com_w_inst_n531,
         round_inst_S_1__sbox_inst_com_w_inst_n530,
         round_inst_S_1__sbox_inst_com_w_inst_n529,
         round_inst_S_1__sbox_inst_com_w_inst_n528,
         round_inst_S_1__sbox_inst_com_w_inst_n527,
         round_inst_S_1__sbox_inst_com_w_inst_n526,
         round_inst_S_1__sbox_inst_com_w_inst_n525,
         round_inst_S_1__sbox_inst_com_w_inst_n524,
         round_inst_S_1__sbox_inst_com_w_inst_n523,
         round_inst_S_1__sbox_inst_com_w_inst_n522,
         round_inst_S_1__sbox_inst_com_w_inst_n521,
         round_inst_S_1__sbox_inst_com_w_inst_n520,
         round_inst_S_1__sbox_inst_com_w_inst_n519,
         round_inst_S_1__sbox_inst_com_w_inst_n518,
         round_inst_S_1__sbox_inst_com_w_inst_n517,
         round_inst_S_1__sbox_inst_com_w_inst_n516,
         round_inst_S_1__sbox_inst_com_w_inst_n515,
         round_inst_S_1__sbox_inst_com_w_inst_n514,
         round_inst_S_1__sbox_inst_com_w_inst_n513,
         round_inst_S_1__sbox_inst_com_w_inst_n512,
         round_inst_S_1__sbox_inst_com_w_inst_n511,
         round_inst_S_1__sbox_inst_com_w_inst_n510,
         round_inst_S_1__sbox_inst_com_w_inst_n509,
         round_inst_S_1__sbox_inst_com_w_inst_n508,
         round_inst_S_1__sbox_inst_com_w_inst_n507,
         round_inst_S_1__sbox_inst_com_w_inst_n506,
         round_inst_S_1__sbox_inst_com_w_inst_n505,
         round_inst_S_1__sbox_inst_com_w_inst_n504,
         round_inst_S_1__sbox_inst_com_w_inst_n503,
         round_inst_S_1__sbox_inst_com_w_inst_n502,
         round_inst_S_1__sbox_inst_com_w_inst_n501,
         round_inst_S_1__sbox_inst_com_w_inst_n500,
         round_inst_S_1__sbox_inst_com_w_inst_n499,
         round_inst_S_1__sbox_inst_com_w_inst_n498,
         round_inst_S_1__sbox_inst_com_w_inst_n497,
         round_inst_S_1__sbox_inst_com_w_inst_n496,
         round_inst_S_1__sbox_inst_com_w_inst_n495,
         round_inst_S_1__sbox_inst_com_w_inst_n494,
         round_inst_S_1__sbox_inst_com_w_inst_n493,
         round_inst_S_1__sbox_inst_com_w_inst_n492,
         round_inst_S_1__sbox_inst_com_w_inst_n491,
         round_inst_S_1__sbox_inst_com_w_inst_n490,
         round_inst_S_1__sbox_inst_com_w_inst_n489,
         round_inst_S_1__sbox_inst_com_w_inst_n488,
         round_inst_S_1__sbox_inst_com_w_inst_n487,
         round_inst_S_1__sbox_inst_com_w_inst_n486,
         round_inst_S_1__sbox_inst_com_w_inst_n485,
         round_inst_S_1__sbox_inst_com_w_inst_n484,
         round_inst_S_1__sbox_inst_com_w_inst_n483,
         round_inst_S_1__sbox_inst_com_w_inst_n482,
         round_inst_S_1__sbox_inst_com_w_inst_n481,
         round_inst_S_1__sbox_inst_com_w_inst_n480,
         round_inst_S_1__sbox_inst_com_w_inst_n479,
         round_inst_S_1__sbox_inst_com_w_inst_n478,
         round_inst_S_1__sbox_inst_com_w_inst_n477,
         round_inst_S_1__sbox_inst_com_w_inst_n476,
         round_inst_S_1__sbox_inst_com_w_inst_n475,
         round_inst_S_1__sbox_inst_com_w_inst_n474,
         round_inst_S_1__sbox_inst_com_w_inst_n473,
         round_inst_S_1__sbox_inst_com_w_inst_n472,
         round_inst_S_1__sbox_inst_com_w_inst_n471,
         round_inst_S_1__sbox_inst_com_w_inst_n470,
         round_inst_S_1__sbox_inst_com_w_inst_n469,
         round_inst_S_1__sbox_inst_com_w_inst_n468,
         round_inst_S_1__sbox_inst_com_w_inst_n467,
         round_inst_S_1__sbox_inst_com_w_inst_n466,
         round_inst_S_1__sbox_inst_com_w_inst_n465,
         round_inst_S_1__sbox_inst_com_w_inst_n464,
         round_inst_S_1__sbox_inst_com_w_inst_n463,
         round_inst_S_1__sbox_inst_com_w_inst_n462,
         round_inst_S_1__sbox_inst_com_w_inst_n461,
         round_inst_S_1__sbox_inst_com_w_inst_n460,
         round_inst_S_1__sbox_inst_com_w_inst_n459,
         round_inst_S_1__sbox_inst_com_w_inst_n458,
         round_inst_S_1__sbox_inst_com_w_inst_n457,
         round_inst_S_1__sbox_inst_com_w_inst_n456,
         round_inst_S_1__sbox_inst_com_w_inst_n455,
         round_inst_S_1__sbox_inst_com_w_inst_n454,
         round_inst_S_1__sbox_inst_com_w_inst_n453,
         round_inst_S_1__sbox_inst_com_w_inst_n452,
         round_inst_S_1__sbox_inst_com_w_inst_n451,
         round_inst_S_1__sbox_inst_com_w_inst_n450,
         round_inst_S_1__sbox_inst_com_w_inst_n449,
         round_inst_S_1__sbox_inst_com_w_inst_n448,
         round_inst_S_1__sbox_inst_com_w_inst_n447,
         round_inst_S_1__sbox_inst_com_w_inst_n446,
         round_inst_S_1__sbox_inst_com_w_inst_n445,
         round_inst_S_1__sbox_inst_com_w_inst_n444,
         round_inst_S_1__sbox_inst_com_w_inst_n443,
         round_inst_S_1__sbox_inst_com_w_inst_n442,
         round_inst_S_1__sbox_inst_com_w_inst_n441,
         round_inst_S_1__sbox_inst_com_w_inst_n440,
         round_inst_S_1__sbox_inst_com_w_inst_n439,
         round_inst_S_1__sbox_inst_com_w_inst_n438,
         round_inst_S_1__sbox_inst_com_w_inst_n437,
         round_inst_S_1__sbox_inst_com_w_inst_n436,
         round_inst_S_1__sbox_inst_com_w_inst_n435,
         round_inst_S_1__sbox_inst_com_w_inst_n434,
         round_inst_S_1__sbox_inst_com_w_inst_n433,
         round_inst_S_1__sbox_inst_com_w_inst_n432,
         round_inst_S_1__sbox_inst_com_w_inst_n431,
         round_inst_S_1__sbox_inst_com_w_inst_n430,
         round_inst_S_1__sbox_inst_com_w_inst_n429,
         round_inst_S_1__sbox_inst_com_w_inst_n428,
         round_inst_S_1__sbox_inst_com_w_inst_n427,
         round_inst_S_1__sbox_inst_com_w_inst_n426,
         round_inst_S_1__sbox_inst_com_w_inst_n425,
         round_inst_S_1__sbox_inst_com_w_inst_n424,
         round_inst_S_1__sbox_inst_com_w_inst_n423,
         round_inst_S_1__sbox_inst_com_w_inst_n422,
         round_inst_S_1__sbox_inst_com_w_inst_n421,
         round_inst_S_1__sbox_inst_com_w_inst_n420,
         round_inst_S_1__sbox_inst_com_w_inst_n419,
         round_inst_S_1__sbox_inst_com_w_inst_n418,
         round_inst_S_1__sbox_inst_com_w_inst_n417,
         round_inst_S_1__sbox_inst_com_w_inst_n416,
         round_inst_S_1__sbox_inst_com_w_inst_n415,
         round_inst_S_1__sbox_inst_com_w_inst_n414,
         round_inst_S_1__sbox_inst_com_w_inst_n413,
         round_inst_S_1__sbox_inst_com_w_inst_n412,
         round_inst_S_1__sbox_inst_com_w_inst_n411,
         round_inst_S_1__sbox_inst_com_w_inst_n410,
         round_inst_S_1__sbox_inst_com_w_inst_n409,
         round_inst_S_1__sbox_inst_com_w_inst_n408,
         round_inst_S_1__sbox_inst_com_w_inst_n407,
         round_inst_S_1__sbox_inst_com_w_inst_n406,
         round_inst_S_1__sbox_inst_com_w_inst_n405,
         round_inst_S_1__sbox_inst_com_w_inst_n404,
         round_inst_S_1__sbox_inst_com_w_inst_n403,
         round_inst_S_1__sbox_inst_com_w_inst_n402,
         round_inst_S_1__sbox_inst_com_w_inst_n401,
         round_inst_S_1__sbox_inst_com_w_inst_n400,
         round_inst_S_1__sbox_inst_com_w_inst_n399,
         round_inst_S_1__sbox_inst_com_w_inst_n398,
         round_inst_S_1__sbox_inst_com_w_inst_n397,
         round_inst_S_1__sbox_inst_com_w_inst_n396,
         round_inst_S_1__sbox_inst_com_w_inst_n395,
         round_inst_S_1__sbox_inst_com_x_inst_n512,
         round_inst_S_1__sbox_inst_com_x_inst_n511,
         round_inst_S_1__sbox_inst_com_x_inst_n510,
         round_inst_S_1__sbox_inst_com_x_inst_n509,
         round_inst_S_1__sbox_inst_com_x_inst_n508,
         round_inst_S_1__sbox_inst_com_x_inst_n507,
         round_inst_S_1__sbox_inst_com_x_inst_n506,
         round_inst_S_1__sbox_inst_com_x_inst_n505,
         round_inst_S_1__sbox_inst_com_x_inst_n504,
         round_inst_S_1__sbox_inst_com_x_inst_n503,
         round_inst_S_1__sbox_inst_com_x_inst_n502,
         round_inst_S_1__sbox_inst_com_x_inst_n501,
         round_inst_S_1__sbox_inst_com_x_inst_n500,
         round_inst_S_1__sbox_inst_com_x_inst_n499,
         round_inst_S_1__sbox_inst_com_x_inst_n498,
         round_inst_S_1__sbox_inst_com_x_inst_n497,
         round_inst_S_1__sbox_inst_com_x_inst_n496,
         round_inst_S_1__sbox_inst_com_x_inst_n495,
         round_inst_S_1__sbox_inst_com_x_inst_n494,
         round_inst_S_1__sbox_inst_com_x_inst_n493,
         round_inst_S_1__sbox_inst_com_x_inst_n492,
         round_inst_S_1__sbox_inst_com_x_inst_n491,
         round_inst_S_1__sbox_inst_com_x_inst_n490,
         round_inst_S_1__sbox_inst_com_x_inst_n489,
         round_inst_S_1__sbox_inst_com_x_inst_n488,
         round_inst_S_1__sbox_inst_com_x_inst_n487,
         round_inst_S_1__sbox_inst_com_x_inst_n486,
         round_inst_S_1__sbox_inst_com_x_inst_n485,
         round_inst_S_1__sbox_inst_com_x_inst_n484,
         round_inst_S_1__sbox_inst_com_x_inst_n483,
         round_inst_S_1__sbox_inst_com_x_inst_n482,
         round_inst_S_1__sbox_inst_com_x_inst_n481,
         round_inst_S_1__sbox_inst_com_x_inst_n480,
         round_inst_S_1__sbox_inst_com_x_inst_n479,
         round_inst_S_1__sbox_inst_com_x_inst_n478,
         round_inst_S_1__sbox_inst_com_x_inst_n477,
         round_inst_S_1__sbox_inst_com_x_inst_n476,
         round_inst_S_1__sbox_inst_com_x_inst_n475,
         round_inst_S_1__sbox_inst_com_x_inst_n474,
         round_inst_S_1__sbox_inst_com_x_inst_n473,
         round_inst_S_1__sbox_inst_com_x_inst_n472,
         round_inst_S_1__sbox_inst_com_x_inst_n471,
         round_inst_S_1__sbox_inst_com_x_inst_n470,
         round_inst_S_1__sbox_inst_com_x_inst_n469,
         round_inst_S_1__sbox_inst_com_x_inst_n468,
         round_inst_S_1__sbox_inst_com_x_inst_n467,
         round_inst_S_1__sbox_inst_com_x_inst_n466,
         round_inst_S_1__sbox_inst_com_x_inst_n465,
         round_inst_S_1__sbox_inst_com_x_inst_n464,
         round_inst_S_1__sbox_inst_com_x_inst_n463,
         round_inst_S_1__sbox_inst_com_x_inst_n462,
         round_inst_S_1__sbox_inst_com_x_inst_n461,
         round_inst_S_1__sbox_inst_com_x_inst_n460,
         round_inst_S_1__sbox_inst_com_x_inst_n459,
         round_inst_S_1__sbox_inst_com_x_inst_n458,
         round_inst_S_1__sbox_inst_com_x_inst_n457,
         round_inst_S_1__sbox_inst_com_x_inst_n456,
         round_inst_S_1__sbox_inst_com_x_inst_n455,
         round_inst_S_1__sbox_inst_com_x_inst_n454,
         round_inst_S_1__sbox_inst_com_x_inst_n453,
         round_inst_S_1__sbox_inst_com_x_inst_n452,
         round_inst_S_1__sbox_inst_com_x_inst_n451,
         round_inst_S_1__sbox_inst_com_x_inst_n450,
         round_inst_S_1__sbox_inst_com_x_inst_n449,
         round_inst_S_1__sbox_inst_com_x_inst_n448,
         round_inst_S_1__sbox_inst_com_x_inst_n447,
         round_inst_S_1__sbox_inst_com_x_inst_n446,
         round_inst_S_1__sbox_inst_com_x_inst_n445,
         round_inst_S_1__sbox_inst_com_x_inst_n444,
         round_inst_S_1__sbox_inst_com_x_inst_n443,
         round_inst_S_1__sbox_inst_com_x_inst_n442,
         round_inst_S_1__sbox_inst_com_x_inst_n441,
         round_inst_S_1__sbox_inst_com_x_inst_n440,
         round_inst_S_1__sbox_inst_com_x_inst_n439,
         round_inst_S_1__sbox_inst_com_x_inst_n438,
         round_inst_S_1__sbox_inst_com_x_inst_n437,
         round_inst_S_1__sbox_inst_com_x_inst_n436,
         round_inst_S_1__sbox_inst_com_x_inst_n435,
         round_inst_S_1__sbox_inst_com_x_inst_n434,
         round_inst_S_1__sbox_inst_com_x_inst_n433,
         round_inst_S_1__sbox_inst_com_x_inst_n432,
         round_inst_S_1__sbox_inst_com_x_inst_n431,
         round_inst_S_1__sbox_inst_com_x_inst_n430,
         round_inst_S_1__sbox_inst_com_x_inst_n429,
         round_inst_S_1__sbox_inst_com_x_inst_n428,
         round_inst_S_1__sbox_inst_com_x_inst_n427,
         round_inst_S_1__sbox_inst_com_x_inst_n426,
         round_inst_S_1__sbox_inst_com_x_inst_n425,
         round_inst_S_1__sbox_inst_com_x_inst_n424,
         round_inst_S_1__sbox_inst_com_x_inst_n423,
         round_inst_S_1__sbox_inst_com_x_inst_n422,
         round_inst_S_1__sbox_inst_com_x_inst_n421,
         round_inst_S_1__sbox_inst_com_x_inst_n420,
         round_inst_S_1__sbox_inst_com_x_inst_n419,
         round_inst_S_1__sbox_inst_com_x_inst_n418,
         round_inst_S_1__sbox_inst_com_x_inst_n417,
         round_inst_S_1__sbox_inst_com_x_inst_n416,
         round_inst_S_1__sbox_inst_com_x_inst_n415,
         round_inst_S_1__sbox_inst_com_x_inst_n414,
         round_inst_S_1__sbox_inst_com_x_inst_n413,
         round_inst_S_1__sbox_inst_com_x_inst_n412,
         round_inst_S_1__sbox_inst_com_x_inst_n411,
         round_inst_S_1__sbox_inst_com_x_inst_n410,
         round_inst_S_1__sbox_inst_com_x_inst_n409,
         round_inst_S_1__sbox_inst_com_x_inst_n408,
         round_inst_S_1__sbox_inst_com_x_inst_n407,
         round_inst_S_1__sbox_inst_com_x_inst_n406,
         round_inst_S_1__sbox_inst_com_x_inst_n405,
         round_inst_S_1__sbox_inst_com_x_inst_n404,
         round_inst_S_1__sbox_inst_com_x_inst_n403,
         round_inst_S_1__sbox_inst_com_x_inst_n402,
         round_inst_S_1__sbox_inst_com_x_inst_n401,
         round_inst_S_1__sbox_inst_com_x_inst_n400,
         round_inst_S_1__sbox_inst_com_x_inst_n399,
         round_inst_S_1__sbox_inst_com_x_inst_n398,
         round_inst_S_1__sbox_inst_com_x_inst_n397,
         round_inst_S_1__sbox_inst_com_x_inst_n396,
         round_inst_S_1__sbox_inst_com_x_inst_n395,
         round_inst_S_1__sbox_inst_com_x_inst_n394,
         round_inst_S_1__sbox_inst_com_x_inst_n393,
         round_inst_S_1__sbox_inst_com_x_inst_n392,
         round_inst_S_1__sbox_inst_com_x_inst_n391,
         round_inst_S_1__sbox_inst_com_x_inst_n390,
         round_inst_S_1__sbox_inst_com_x_inst_n389,
         round_inst_S_1__sbox_inst_com_x_inst_n388,
         round_inst_S_1__sbox_inst_com_x_inst_n387,
         round_inst_S_1__sbox_inst_com_x_inst_n386,
         round_inst_S_1__sbox_inst_com_x_inst_n385,
         round_inst_S_1__sbox_inst_com_x_inst_n384,
         round_inst_S_1__sbox_inst_com_x_inst_n383,
         round_inst_S_1__sbox_inst_com_x_inst_n382,
         round_inst_S_1__sbox_inst_com_x_inst_n381,
         round_inst_S_1__sbox_inst_com_y_inst_n518,
         round_inst_S_1__sbox_inst_com_y_inst_n517,
         round_inst_S_1__sbox_inst_com_y_inst_n516,
         round_inst_S_1__sbox_inst_com_y_inst_n515,
         round_inst_S_1__sbox_inst_com_y_inst_n514,
         round_inst_S_1__sbox_inst_com_y_inst_n513,
         round_inst_S_1__sbox_inst_com_y_inst_n512,
         round_inst_S_1__sbox_inst_com_y_inst_n511,
         round_inst_S_1__sbox_inst_com_y_inst_n510,
         round_inst_S_1__sbox_inst_com_y_inst_n509,
         round_inst_S_1__sbox_inst_com_y_inst_n508,
         round_inst_S_1__sbox_inst_com_y_inst_n507,
         round_inst_S_1__sbox_inst_com_y_inst_n506,
         round_inst_S_1__sbox_inst_com_y_inst_n505,
         round_inst_S_1__sbox_inst_com_y_inst_n504,
         round_inst_S_1__sbox_inst_com_y_inst_n503,
         round_inst_S_1__sbox_inst_com_y_inst_n502,
         round_inst_S_1__sbox_inst_com_y_inst_n501,
         round_inst_S_1__sbox_inst_com_y_inst_n500,
         round_inst_S_1__sbox_inst_com_y_inst_n499,
         round_inst_S_1__sbox_inst_com_y_inst_n498,
         round_inst_S_1__sbox_inst_com_y_inst_n497,
         round_inst_S_1__sbox_inst_com_y_inst_n496,
         round_inst_S_1__sbox_inst_com_y_inst_n495,
         round_inst_S_1__sbox_inst_com_y_inst_n494,
         round_inst_S_1__sbox_inst_com_y_inst_n493,
         round_inst_S_1__sbox_inst_com_y_inst_n492,
         round_inst_S_1__sbox_inst_com_y_inst_n491,
         round_inst_S_1__sbox_inst_com_y_inst_n490,
         round_inst_S_1__sbox_inst_com_y_inst_n489,
         round_inst_S_1__sbox_inst_com_y_inst_n488,
         round_inst_S_1__sbox_inst_com_y_inst_n487,
         round_inst_S_1__sbox_inst_com_y_inst_n486,
         round_inst_S_1__sbox_inst_com_y_inst_n485,
         round_inst_S_1__sbox_inst_com_y_inst_n484,
         round_inst_S_1__sbox_inst_com_y_inst_n483,
         round_inst_S_1__sbox_inst_com_y_inst_n482,
         round_inst_S_1__sbox_inst_com_y_inst_n481,
         round_inst_S_1__sbox_inst_com_y_inst_n480,
         round_inst_S_1__sbox_inst_com_y_inst_n479,
         round_inst_S_1__sbox_inst_com_y_inst_n478,
         round_inst_S_1__sbox_inst_com_y_inst_n477,
         round_inst_S_1__sbox_inst_com_y_inst_n476,
         round_inst_S_1__sbox_inst_com_y_inst_n475,
         round_inst_S_1__sbox_inst_com_y_inst_n474,
         round_inst_S_1__sbox_inst_com_y_inst_n473,
         round_inst_S_1__sbox_inst_com_y_inst_n472,
         round_inst_S_1__sbox_inst_com_y_inst_n471,
         round_inst_S_1__sbox_inst_com_y_inst_n470,
         round_inst_S_1__sbox_inst_com_y_inst_n469,
         round_inst_S_1__sbox_inst_com_y_inst_n468,
         round_inst_S_1__sbox_inst_com_y_inst_n467,
         round_inst_S_1__sbox_inst_com_y_inst_n466,
         round_inst_S_1__sbox_inst_com_y_inst_n465,
         round_inst_S_1__sbox_inst_com_y_inst_n464,
         round_inst_S_1__sbox_inst_com_y_inst_n463,
         round_inst_S_1__sbox_inst_com_y_inst_n462,
         round_inst_S_1__sbox_inst_com_y_inst_n461,
         round_inst_S_1__sbox_inst_com_y_inst_n460,
         round_inst_S_1__sbox_inst_com_y_inst_n459,
         round_inst_S_1__sbox_inst_com_y_inst_n458,
         round_inst_S_1__sbox_inst_com_y_inst_n457,
         round_inst_S_1__sbox_inst_com_y_inst_n456,
         round_inst_S_1__sbox_inst_com_y_inst_n455,
         round_inst_S_1__sbox_inst_com_y_inst_n454,
         round_inst_S_1__sbox_inst_com_y_inst_n453,
         round_inst_S_1__sbox_inst_com_y_inst_n452,
         round_inst_S_1__sbox_inst_com_y_inst_n451,
         round_inst_S_1__sbox_inst_com_y_inst_n450,
         round_inst_S_1__sbox_inst_com_y_inst_n449,
         round_inst_S_1__sbox_inst_com_y_inst_n448,
         round_inst_S_1__sbox_inst_com_y_inst_n447,
         round_inst_S_1__sbox_inst_com_y_inst_n446,
         round_inst_S_1__sbox_inst_com_y_inst_n445,
         round_inst_S_1__sbox_inst_com_y_inst_n444,
         round_inst_S_1__sbox_inst_com_y_inst_n443,
         round_inst_S_1__sbox_inst_com_y_inst_n442,
         round_inst_S_1__sbox_inst_com_y_inst_n441,
         round_inst_S_1__sbox_inst_com_y_inst_n440,
         round_inst_S_1__sbox_inst_com_y_inst_n439,
         round_inst_S_1__sbox_inst_com_y_inst_n438,
         round_inst_S_1__sbox_inst_com_y_inst_n437,
         round_inst_S_1__sbox_inst_com_y_inst_n436,
         round_inst_S_1__sbox_inst_com_y_inst_n435,
         round_inst_S_1__sbox_inst_com_y_inst_n434,
         round_inst_S_1__sbox_inst_com_y_inst_n433,
         round_inst_S_1__sbox_inst_com_y_inst_n432,
         round_inst_S_1__sbox_inst_com_y_inst_n431,
         round_inst_S_1__sbox_inst_com_y_inst_n430,
         round_inst_S_1__sbox_inst_com_y_inst_n429,
         round_inst_S_1__sbox_inst_com_y_inst_n428,
         round_inst_S_1__sbox_inst_com_y_inst_n427,
         round_inst_S_1__sbox_inst_com_y_inst_n426,
         round_inst_S_1__sbox_inst_com_y_inst_n425,
         round_inst_S_1__sbox_inst_com_y_inst_n424,
         round_inst_S_1__sbox_inst_com_y_inst_n423,
         round_inst_S_1__sbox_inst_com_y_inst_n422,
         round_inst_S_1__sbox_inst_com_y_inst_n421,
         round_inst_S_1__sbox_inst_com_y_inst_n420,
         round_inst_S_1__sbox_inst_com_y_inst_n419,
         round_inst_S_1__sbox_inst_com_y_inst_n418,
         round_inst_S_1__sbox_inst_com_y_inst_n417,
         round_inst_S_1__sbox_inst_com_y_inst_n416,
         round_inst_S_1__sbox_inst_com_y_inst_n415,
         round_inst_S_1__sbox_inst_com_y_inst_n414,
         round_inst_S_1__sbox_inst_com_y_inst_n413,
         round_inst_S_1__sbox_inst_com_y_inst_n412,
         round_inst_S_1__sbox_inst_com_y_inst_n411,
         round_inst_S_1__sbox_inst_com_y_inst_n410,
         round_inst_S_1__sbox_inst_com_y_inst_n409,
         round_inst_S_1__sbox_inst_com_y_inst_n408,
         round_inst_S_1__sbox_inst_com_y_inst_n407,
         round_inst_S_1__sbox_inst_com_y_inst_n406,
         round_inst_S_1__sbox_inst_com_y_inst_n405,
         round_inst_S_1__sbox_inst_com_y_inst_n404,
         round_inst_S_1__sbox_inst_com_y_inst_n403,
         round_inst_S_1__sbox_inst_com_y_inst_n402,
         round_inst_S_1__sbox_inst_com_y_inst_n401,
         round_inst_S_1__sbox_inst_com_y_inst_n400,
         round_inst_S_1__sbox_inst_com_y_inst_n399,
         round_inst_S_1__sbox_inst_com_y_inst_n398,
         round_inst_S_1__sbox_inst_com_y_inst_n397,
         round_inst_S_1__sbox_inst_com_y_inst_n396,
         round_inst_S_1__sbox_inst_com_y_inst_n395,
         round_inst_S_1__sbox_inst_com_y_inst_n394,
         round_inst_S_1__sbox_inst_com_y_inst_n393,
         round_inst_S_1__sbox_inst_com_y_inst_n392,
         round_inst_S_1__sbox_inst_com_y_inst_n391,
         round_inst_S_1__sbox_inst_com_y_inst_n390,
         round_inst_S_1__sbox_inst_com_y_inst_n389,
         round_inst_S_1__sbox_inst_com_y_inst_n388,
         round_inst_S_1__sbox_inst_com_y_inst_n387,
         round_inst_S_1__sbox_inst_com_y_inst_n386,
         round_inst_S_1__sbox_inst_com_z_inst_n517,
         round_inst_S_1__sbox_inst_com_z_inst_n516,
         round_inst_S_1__sbox_inst_com_z_inst_n515,
         round_inst_S_1__sbox_inst_com_z_inst_n514,
         round_inst_S_1__sbox_inst_com_z_inst_n513,
         round_inst_S_1__sbox_inst_com_z_inst_n512,
         round_inst_S_1__sbox_inst_com_z_inst_n511,
         round_inst_S_1__sbox_inst_com_z_inst_n510,
         round_inst_S_1__sbox_inst_com_z_inst_n509,
         round_inst_S_1__sbox_inst_com_z_inst_n508,
         round_inst_S_1__sbox_inst_com_z_inst_n507,
         round_inst_S_1__sbox_inst_com_z_inst_n506,
         round_inst_S_1__sbox_inst_com_z_inst_n505,
         round_inst_S_1__sbox_inst_com_z_inst_n504,
         round_inst_S_1__sbox_inst_com_z_inst_n503,
         round_inst_S_1__sbox_inst_com_z_inst_n502,
         round_inst_S_1__sbox_inst_com_z_inst_n501,
         round_inst_S_1__sbox_inst_com_z_inst_n500,
         round_inst_S_1__sbox_inst_com_z_inst_n499,
         round_inst_S_1__sbox_inst_com_z_inst_n498,
         round_inst_S_1__sbox_inst_com_z_inst_n497,
         round_inst_S_1__sbox_inst_com_z_inst_n496,
         round_inst_S_1__sbox_inst_com_z_inst_n495,
         round_inst_S_1__sbox_inst_com_z_inst_n494,
         round_inst_S_1__sbox_inst_com_z_inst_n493,
         round_inst_S_1__sbox_inst_com_z_inst_n492,
         round_inst_S_1__sbox_inst_com_z_inst_n491,
         round_inst_S_1__sbox_inst_com_z_inst_n490,
         round_inst_S_1__sbox_inst_com_z_inst_n489,
         round_inst_S_1__sbox_inst_com_z_inst_n488,
         round_inst_S_1__sbox_inst_com_z_inst_n487,
         round_inst_S_1__sbox_inst_com_z_inst_n486,
         round_inst_S_1__sbox_inst_com_z_inst_n485,
         round_inst_S_1__sbox_inst_com_z_inst_n484,
         round_inst_S_1__sbox_inst_com_z_inst_n483,
         round_inst_S_1__sbox_inst_com_z_inst_n482,
         round_inst_S_1__sbox_inst_com_z_inst_n481,
         round_inst_S_1__sbox_inst_com_z_inst_n480,
         round_inst_S_1__sbox_inst_com_z_inst_n479,
         round_inst_S_1__sbox_inst_com_z_inst_n478,
         round_inst_S_1__sbox_inst_com_z_inst_n477,
         round_inst_S_1__sbox_inst_com_z_inst_n476,
         round_inst_S_1__sbox_inst_com_z_inst_n475,
         round_inst_S_1__sbox_inst_com_z_inst_n474,
         round_inst_S_1__sbox_inst_com_z_inst_n473,
         round_inst_S_1__sbox_inst_com_z_inst_n472,
         round_inst_S_1__sbox_inst_com_z_inst_n471,
         round_inst_S_1__sbox_inst_com_z_inst_n470,
         round_inst_S_1__sbox_inst_com_z_inst_n469,
         round_inst_S_1__sbox_inst_com_z_inst_n468,
         round_inst_S_1__sbox_inst_com_z_inst_n467,
         round_inst_S_1__sbox_inst_com_z_inst_n466,
         round_inst_S_1__sbox_inst_com_z_inst_n465,
         round_inst_S_1__sbox_inst_com_z_inst_n464,
         round_inst_S_1__sbox_inst_com_z_inst_n463,
         round_inst_S_1__sbox_inst_com_z_inst_n462,
         round_inst_S_1__sbox_inst_com_z_inst_n461,
         round_inst_S_1__sbox_inst_com_z_inst_n460,
         round_inst_S_1__sbox_inst_com_z_inst_n459,
         round_inst_S_1__sbox_inst_com_z_inst_n458,
         round_inst_S_1__sbox_inst_com_z_inst_n457,
         round_inst_S_1__sbox_inst_com_z_inst_n456,
         round_inst_S_1__sbox_inst_com_z_inst_n455,
         round_inst_S_1__sbox_inst_com_z_inst_n454,
         round_inst_S_1__sbox_inst_com_z_inst_n453,
         round_inst_S_1__sbox_inst_com_z_inst_n452,
         round_inst_S_1__sbox_inst_com_z_inst_n451,
         round_inst_S_1__sbox_inst_com_z_inst_n450,
         round_inst_S_1__sbox_inst_com_z_inst_n449,
         round_inst_S_1__sbox_inst_com_z_inst_n448,
         round_inst_S_1__sbox_inst_com_z_inst_n447,
         round_inst_S_1__sbox_inst_com_z_inst_n446,
         round_inst_S_1__sbox_inst_com_z_inst_n445,
         round_inst_S_1__sbox_inst_com_z_inst_n444,
         round_inst_S_1__sbox_inst_com_z_inst_n443,
         round_inst_S_1__sbox_inst_com_z_inst_n442,
         round_inst_S_1__sbox_inst_com_z_inst_n441,
         round_inst_S_1__sbox_inst_com_z_inst_n440,
         round_inst_S_1__sbox_inst_com_z_inst_n439,
         round_inst_S_1__sbox_inst_com_z_inst_n438,
         round_inst_S_1__sbox_inst_com_z_inst_n437,
         round_inst_S_1__sbox_inst_com_z_inst_n436,
         round_inst_S_1__sbox_inst_com_z_inst_n435,
         round_inst_S_1__sbox_inst_com_z_inst_n434,
         round_inst_S_1__sbox_inst_com_z_inst_n433,
         round_inst_S_1__sbox_inst_com_z_inst_n432,
         round_inst_S_1__sbox_inst_com_z_inst_n431,
         round_inst_S_1__sbox_inst_com_z_inst_n430,
         round_inst_S_1__sbox_inst_com_z_inst_n429,
         round_inst_S_1__sbox_inst_com_z_inst_n428,
         round_inst_S_1__sbox_inst_com_z_inst_n427,
         round_inst_S_1__sbox_inst_com_z_inst_n426,
         round_inst_S_1__sbox_inst_com_z_inst_n425,
         round_inst_S_1__sbox_inst_com_z_inst_n424,
         round_inst_S_1__sbox_inst_com_z_inst_n423,
         round_inst_S_1__sbox_inst_com_z_inst_n422,
         round_inst_S_1__sbox_inst_com_z_inst_n421,
         round_inst_S_1__sbox_inst_com_z_inst_n420,
         round_inst_S_1__sbox_inst_com_z_inst_n419,
         round_inst_S_1__sbox_inst_com_z_inst_n418,
         round_inst_S_1__sbox_inst_com_z_inst_n417,
         round_inst_S_1__sbox_inst_com_z_inst_n416,
         round_inst_S_1__sbox_inst_com_z_inst_n415,
         round_inst_S_1__sbox_inst_com_z_inst_n414,
         round_inst_S_1__sbox_inst_com_z_inst_n413,
         round_inst_S_1__sbox_inst_com_z_inst_n412,
         round_inst_S_1__sbox_inst_com_z_inst_n411,
         round_inst_S_1__sbox_inst_com_z_inst_n410,
         round_inst_S_1__sbox_inst_com_z_inst_n409,
         round_inst_S_1__sbox_inst_com_z_inst_n408,
         round_inst_S_1__sbox_inst_com_z_inst_n407,
         round_inst_S_1__sbox_inst_com_z_inst_n406,
         round_inst_S_1__sbox_inst_com_z_inst_n405,
         round_inst_S_1__sbox_inst_com_z_inst_n404,
         round_inst_S_1__sbox_inst_com_z_inst_n403,
         round_inst_S_1__sbox_inst_com_z_inst_n402,
         round_inst_S_1__sbox_inst_com_z_inst_n401,
         round_inst_S_1__sbox_inst_com_z_inst_n400,
         round_inst_S_1__sbox_inst_com_z_inst_n399,
         round_inst_S_1__sbox_inst_com_z_inst_n398,
         round_inst_S_1__sbox_inst_com_z_inst_n397,
         round_inst_S_1__sbox_inst_com_z_inst_n396,
         round_inst_S_1__sbox_inst_com_z_inst_n395,
         round_inst_S_1__sbox_inst_com_z_inst_n394,
         round_inst_S_1__sbox_inst_com_z_inst_n393,
         round_inst_S_1__sbox_inst_com_z_inst_n392,
         round_inst_S_1__sbox_inst_com_z_inst_n391,
         round_inst_S_1__sbox_inst_com_z_inst_n390,
         round_inst_S_2__sbox_inst_n6, round_inst_S_2__sbox_inst_n5,
         round_inst_S_2__sbox_inst_n4, round_inst_S_2__sbox_inst_n3,
         round_inst_S_2__sbox_inst_n2, round_inst_S_2__sbox_inst_n1,
         round_inst_S_2__sbox_inst_com_w_inst_n532,
         round_inst_S_2__sbox_inst_com_w_inst_n531,
         round_inst_S_2__sbox_inst_com_w_inst_n530,
         round_inst_S_2__sbox_inst_com_w_inst_n529,
         round_inst_S_2__sbox_inst_com_w_inst_n528,
         round_inst_S_2__sbox_inst_com_w_inst_n527,
         round_inst_S_2__sbox_inst_com_w_inst_n526,
         round_inst_S_2__sbox_inst_com_w_inst_n525,
         round_inst_S_2__sbox_inst_com_w_inst_n524,
         round_inst_S_2__sbox_inst_com_w_inst_n523,
         round_inst_S_2__sbox_inst_com_w_inst_n522,
         round_inst_S_2__sbox_inst_com_w_inst_n521,
         round_inst_S_2__sbox_inst_com_w_inst_n520,
         round_inst_S_2__sbox_inst_com_w_inst_n519,
         round_inst_S_2__sbox_inst_com_w_inst_n518,
         round_inst_S_2__sbox_inst_com_w_inst_n517,
         round_inst_S_2__sbox_inst_com_w_inst_n516,
         round_inst_S_2__sbox_inst_com_w_inst_n515,
         round_inst_S_2__sbox_inst_com_w_inst_n514,
         round_inst_S_2__sbox_inst_com_w_inst_n513,
         round_inst_S_2__sbox_inst_com_w_inst_n512,
         round_inst_S_2__sbox_inst_com_w_inst_n511,
         round_inst_S_2__sbox_inst_com_w_inst_n510,
         round_inst_S_2__sbox_inst_com_w_inst_n509,
         round_inst_S_2__sbox_inst_com_w_inst_n508,
         round_inst_S_2__sbox_inst_com_w_inst_n507,
         round_inst_S_2__sbox_inst_com_w_inst_n506,
         round_inst_S_2__sbox_inst_com_w_inst_n505,
         round_inst_S_2__sbox_inst_com_w_inst_n504,
         round_inst_S_2__sbox_inst_com_w_inst_n503,
         round_inst_S_2__sbox_inst_com_w_inst_n502,
         round_inst_S_2__sbox_inst_com_w_inst_n501,
         round_inst_S_2__sbox_inst_com_w_inst_n500,
         round_inst_S_2__sbox_inst_com_w_inst_n499,
         round_inst_S_2__sbox_inst_com_w_inst_n498,
         round_inst_S_2__sbox_inst_com_w_inst_n497,
         round_inst_S_2__sbox_inst_com_w_inst_n496,
         round_inst_S_2__sbox_inst_com_w_inst_n495,
         round_inst_S_2__sbox_inst_com_w_inst_n494,
         round_inst_S_2__sbox_inst_com_w_inst_n493,
         round_inst_S_2__sbox_inst_com_w_inst_n492,
         round_inst_S_2__sbox_inst_com_w_inst_n491,
         round_inst_S_2__sbox_inst_com_w_inst_n490,
         round_inst_S_2__sbox_inst_com_w_inst_n489,
         round_inst_S_2__sbox_inst_com_w_inst_n488,
         round_inst_S_2__sbox_inst_com_w_inst_n487,
         round_inst_S_2__sbox_inst_com_w_inst_n486,
         round_inst_S_2__sbox_inst_com_w_inst_n485,
         round_inst_S_2__sbox_inst_com_w_inst_n484,
         round_inst_S_2__sbox_inst_com_w_inst_n483,
         round_inst_S_2__sbox_inst_com_w_inst_n482,
         round_inst_S_2__sbox_inst_com_w_inst_n481,
         round_inst_S_2__sbox_inst_com_w_inst_n480,
         round_inst_S_2__sbox_inst_com_w_inst_n479,
         round_inst_S_2__sbox_inst_com_w_inst_n478,
         round_inst_S_2__sbox_inst_com_w_inst_n477,
         round_inst_S_2__sbox_inst_com_w_inst_n476,
         round_inst_S_2__sbox_inst_com_w_inst_n475,
         round_inst_S_2__sbox_inst_com_w_inst_n474,
         round_inst_S_2__sbox_inst_com_w_inst_n473,
         round_inst_S_2__sbox_inst_com_w_inst_n472,
         round_inst_S_2__sbox_inst_com_w_inst_n471,
         round_inst_S_2__sbox_inst_com_w_inst_n470,
         round_inst_S_2__sbox_inst_com_w_inst_n469,
         round_inst_S_2__sbox_inst_com_w_inst_n468,
         round_inst_S_2__sbox_inst_com_w_inst_n467,
         round_inst_S_2__sbox_inst_com_w_inst_n466,
         round_inst_S_2__sbox_inst_com_w_inst_n465,
         round_inst_S_2__sbox_inst_com_w_inst_n464,
         round_inst_S_2__sbox_inst_com_w_inst_n463,
         round_inst_S_2__sbox_inst_com_w_inst_n462,
         round_inst_S_2__sbox_inst_com_w_inst_n461,
         round_inst_S_2__sbox_inst_com_w_inst_n460,
         round_inst_S_2__sbox_inst_com_w_inst_n459,
         round_inst_S_2__sbox_inst_com_w_inst_n458,
         round_inst_S_2__sbox_inst_com_w_inst_n457,
         round_inst_S_2__sbox_inst_com_w_inst_n456,
         round_inst_S_2__sbox_inst_com_w_inst_n455,
         round_inst_S_2__sbox_inst_com_w_inst_n454,
         round_inst_S_2__sbox_inst_com_w_inst_n453,
         round_inst_S_2__sbox_inst_com_w_inst_n452,
         round_inst_S_2__sbox_inst_com_w_inst_n451,
         round_inst_S_2__sbox_inst_com_w_inst_n450,
         round_inst_S_2__sbox_inst_com_w_inst_n449,
         round_inst_S_2__sbox_inst_com_w_inst_n448,
         round_inst_S_2__sbox_inst_com_w_inst_n447,
         round_inst_S_2__sbox_inst_com_w_inst_n446,
         round_inst_S_2__sbox_inst_com_w_inst_n445,
         round_inst_S_2__sbox_inst_com_w_inst_n444,
         round_inst_S_2__sbox_inst_com_w_inst_n443,
         round_inst_S_2__sbox_inst_com_w_inst_n442,
         round_inst_S_2__sbox_inst_com_w_inst_n441,
         round_inst_S_2__sbox_inst_com_w_inst_n440,
         round_inst_S_2__sbox_inst_com_w_inst_n439,
         round_inst_S_2__sbox_inst_com_w_inst_n438,
         round_inst_S_2__sbox_inst_com_w_inst_n437,
         round_inst_S_2__sbox_inst_com_w_inst_n436,
         round_inst_S_2__sbox_inst_com_w_inst_n435,
         round_inst_S_2__sbox_inst_com_w_inst_n434,
         round_inst_S_2__sbox_inst_com_w_inst_n433,
         round_inst_S_2__sbox_inst_com_w_inst_n432,
         round_inst_S_2__sbox_inst_com_w_inst_n431,
         round_inst_S_2__sbox_inst_com_w_inst_n430,
         round_inst_S_2__sbox_inst_com_w_inst_n429,
         round_inst_S_2__sbox_inst_com_w_inst_n428,
         round_inst_S_2__sbox_inst_com_w_inst_n427,
         round_inst_S_2__sbox_inst_com_w_inst_n426,
         round_inst_S_2__sbox_inst_com_w_inst_n425,
         round_inst_S_2__sbox_inst_com_w_inst_n424,
         round_inst_S_2__sbox_inst_com_w_inst_n423,
         round_inst_S_2__sbox_inst_com_w_inst_n422,
         round_inst_S_2__sbox_inst_com_w_inst_n421,
         round_inst_S_2__sbox_inst_com_w_inst_n420,
         round_inst_S_2__sbox_inst_com_w_inst_n419,
         round_inst_S_2__sbox_inst_com_w_inst_n418,
         round_inst_S_2__sbox_inst_com_w_inst_n417,
         round_inst_S_2__sbox_inst_com_w_inst_n416,
         round_inst_S_2__sbox_inst_com_w_inst_n415,
         round_inst_S_2__sbox_inst_com_w_inst_n414,
         round_inst_S_2__sbox_inst_com_w_inst_n413,
         round_inst_S_2__sbox_inst_com_w_inst_n412,
         round_inst_S_2__sbox_inst_com_w_inst_n411,
         round_inst_S_2__sbox_inst_com_w_inst_n410,
         round_inst_S_2__sbox_inst_com_w_inst_n409,
         round_inst_S_2__sbox_inst_com_w_inst_n408,
         round_inst_S_2__sbox_inst_com_w_inst_n407,
         round_inst_S_2__sbox_inst_com_w_inst_n406,
         round_inst_S_2__sbox_inst_com_w_inst_n405,
         round_inst_S_2__sbox_inst_com_w_inst_n404,
         round_inst_S_2__sbox_inst_com_w_inst_n403,
         round_inst_S_2__sbox_inst_com_w_inst_n402,
         round_inst_S_2__sbox_inst_com_w_inst_n401,
         round_inst_S_2__sbox_inst_com_w_inst_n400,
         round_inst_S_2__sbox_inst_com_w_inst_n399,
         round_inst_S_2__sbox_inst_com_w_inst_n398,
         round_inst_S_2__sbox_inst_com_w_inst_n397,
         round_inst_S_2__sbox_inst_com_w_inst_n396,
         round_inst_S_2__sbox_inst_com_x_inst_n511,
         round_inst_S_2__sbox_inst_com_x_inst_n510,
         round_inst_S_2__sbox_inst_com_x_inst_n509,
         round_inst_S_2__sbox_inst_com_x_inst_n508,
         round_inst_S_2__sbox_inst_com_x_inst_n507,
         round_inst_S_2__sbox_inst_com_x_inst_n506,
         round_inst_S_2__sbox_inst_com_x_inst_n505,
         round_inst_S_2__sbox_inst_com_x_inst_n504,
         round_inst_S_2__sbox_inst_com_x_inst_n503,
         round_inst_S_2__sbox_inst_com_x_inst_n502,
         round_inst_S_2__sbox_inst_com_x_inst_n501,
         round_inst_S_2__sbox_inst_com_x_inst_n500,
         round_inst_S_2__sbox_inst_com_x_inst_n499,
         round_inst_S_2__sbox_inst_com_x_inst_n498,
         round_inst_S_2__sbox_inst_com_x_inst_n497,
         round_inst_S_2__sbox_inst_com_x_inst_n496,
         round_inst_S_2__sbox_inst_com_x_inst_n495,
         round_inst_S_2__sbox_inst_com_x_inst_n494,
         round_inst_S_2__sbox_inst_com_x_inst_n493,
         round_inst_S_2__sbox_inst_com_x_inst_n492,
         round_inst_S_2__sbox_inst_com_x_inst_n491,
         round_inst_S_2__sbox_inst_com_x_inst_n490,
         round_inst_S_2__sbox_inst_com_x_inst_n489,
         round_inst_S_2__sbox_inst_com_x_inst_n488,
         round_inst_S_2__sbox_inst_com_x_inst_n487,
         round_inst_S_2__sbox_inst_com_x_inst_n486,
         round_inst_S_2__sbox_inst_com_x_inst_n485,
         round_inst_S_2__sbox_inst_com_x_inst_n484,
         round_inst_S_2__sbox_inst_com_x_inst_n483,
         round_inst_S_2__sbox_inst_com_x_inst_n482,
         round_inst_S_2__sbox_inst_com_x_inst_n481,
         round_inst_S_2__sbox_inst_com_x_inst_n480,
         round_inst_S_2__sbox_inst_com_x_inst_n479,
         round_inst_S_2__sbox_inst_com_x_inst_n478,
         round_inst_S_2__sbox_inst_com_x_inst_n477,
         round_inst_S_2__sbox_inst_com_x_inst_n476,
         round_inst_S_2__sbox_inst_com_x_inst_n475,
         round_inst_S_2__sbox_inst_com_x_inst_n474,
         round_inst_S_2__sbox_inst_com_x_inst_n473,
         round_inst_S_2__sbox_inst_com_x_inst_n472,
         round_inst_S_2__sbox_inst_com_x_inst_n471,
         round_inst_S_2__sbox_inst_com_x_inst_n470,
         round_inst_S_2__sbox_inst_com_x_inst_n469,
         round_inst_S_2__sbox_inst_com_x_inst_n468,
         round_inst_S_2__sbox_inst_com_x_inst_n467,
         round_inst_S_2__sbox_inst_com_x_inst_n466,
         round_inst_S_2__sbox_inst_com_x_inst_n465,
         round_inst_S_2__sbox_inst_com_x_inst_n464,
         round_inst_S_2__sbox_inst_com_x_inst_n463,
         round_inst_S_2__sbox_inst_com_x_inst_n462,
         round_inst_S_2__sbox_inst_com_x_inst_n461,
         round_inst_S_2__sbox_inst_com_x_inst_n460,
         round_inst_S_2__sbox_inst_com_x_inst_n459,
         round_inst_S_2__sbox_inst_com_x_inst_n458,
         round_inst_S_2__sbox_inst_com_x_inst_n457,
         round_inst_S_2__sbox_inst_com_x_inst_n456,
         round_inst_S_2__sbox_inst_com_x_inst_n455,
         round_inst_S_2__sbox_inst_com_x_inst_n454,
         round_inst_S_2__sbox_inst_com_x_inst_n453,
         round_inst_S_2__sbox_inst_com_x_inst_n452,
         round_inst_S_2__sbox_inst_com_x_inst_n451,
         round_inst_S_2__sbox_inst_com_x_inst_n450,
         round_inst_S_2__sbox_inst_com_x_inst_n449,
         round_inst_S_2__sbox_inst_com_x_inst_n448,
         round_inst_S_2__sbox_inst_com_x_inst_n447,
         round_inst_S_2__sbox_inst_com_x_inst_n446,
         round_inst_S_2__sbox_inst_com_x_inst_n445,
         round_inst_S_2__sbox_inst_com_x_inst_n444,
         round_inst_S_2__sbox_inst_com_x_inst_n443,
         round_inst_S_2__sbox_inst_com_x_inst_n442,
         round_inst_S_2__sbox_inst_com_x_inst_n441,
         round_inst_S_2__sbox_inst_com_x_inst_n440,
         round_inst_S_2__sbox_inst_com_x_inst_n439,
         round_inst_S_2__sbox_inst_com_x_inst_n438,
         round_inst_S_2__sbox_inst_com_x_inst_n437,
         round_inst_S_2__sbox_inst_com_x_inst_n436,
         round_inst_S_2__sbox_inst_com_x_inst_n435,
         round_inst_S_2__sbox_inst_com_x_inst_n434,
         round_inst_S_2__sbox_inst_com_x_inst_n433,
         round_inst_S_2__sbox_inst_com_x_inst_n432,
         round_inst_S_2__sbox_inst_com_x_inst_n431,
         round_inst_S_2__sbox_inst_com_x_inst_n430,
         round_inst_S_2__sbox_inst_com_x_inst_n429,
         round_inst_S_2__sbox_inst_com_x_inst_n428,
         round_inst_S_2__sbox_inst_com_x_inst_n427,
         round_inst_S_2__sbox_inst_com_x_inst_n426,
         round_inst_S_2__sbox_inst_com_x_inst_n425,
         round_inst_S_2__sbox_inst_com_x_inst_n424,
         round_inst_S_2__sbox_inst_com_x_inst_n423,
         round_inst_S_2__sbox_inst_com_x_inst_n422,
         round_inst_S_2__sbox_inst_com_x_inst_n421,
         round_inst_S_2__sbox_inst_com_x_inst_n420,
         round_inst_S_2__sbox_inst_com_x_inst_n419,
         round_inst_S_2__sbox_inst_com_x_inst_n418,
         round_inst_S_2__sbox_inst_com_x_inst_n417,
         round_inst_S_2__sbox_inst_com_x_inst_n416,
         round_inst_S_2__sbox_inst_com_x_inst_n415,
         round_inst_S_2__sbox_inst_com_x_inst_n414,
         round_inst_S_2__sbox_inst_com_x_inst_n413,
         round_inst_S_2__sbox_inst_com_x_inst_n412,
         round_inst_S_2__sbox_inst_com_x_inst_n411,
         round_inst_S_2__sbox_inst_com_x_inst_n410,
         round_inst_S_2__sbox_inst_com_x_inst_n409,
         round_inst_S_2__sbox_inst_com_x_inst_n408,
         round_inst_S_2__sbox_inst_com_x_inst_n407,
         round_inst_S_2__sbox_inst_com_x_inst_n406,
         round_inst_S_2__sbox_inst_com_x_inst_n405,
         round_inst_S_2__sbox_inst_com_x_inst_n404,
         round_inst_S_2__sbox_inst_com_x_inst_n403,
         round_inst_S_2__sbox_inst_com_x_inst_n402,
         round_inst_S_2__sbox_inst_com_x_inst_n401,
         round_inst_S_2__sbox_inst_com_x_inst_n400,
         round_inst_S_2__sbox_inst_com_x_inst_n399,
         round_inst_S_2__sbox_inst_com_x_inst_n398,
         round_inst_S_2__sbox_inst_com_x_inst_n397,
         round_inst_S_2__sbox_inst_com_x_inst_n396,
         round_inst_S_2__sbox_inst_com_x_inst_n395,
         round_inst_S_2__sbox_inst_com_x_inst_n394,
         round_inst_S_2__sbox_inst_com_x_inst_n393,
         round_inst_S_2__sbox_inst_com_x_inst_n392,
         round_inst_S_2__sbox_inst_com_x_inst_n391,
         round_inst_S_2__sbox_inst_com_x_inst_n390,
         round_inst_S_2__sbox_inst_com_x_inst_n389,
         round_inst_S_2__sbox_inst_com_x_inst_n388,
         round_inst_S_2__sbox_inst_com_x_inst_n387,
         round_inst_S_2__sbox_inst_com_x_inst_n386,
         round_inst_S_2__sbox_inst_com_x_inst_n385,
         round_inst_S_2__sbox_inst_com_x_inst_n384,
         round_inst_S_2__sbox_inst_com_x_inst_n383,
         round_inst_S_2__sbox_inst_com_x_inst_n382,
         round_inst_S_2__sbox_inst_com_x_inst_n381,
         round_inst_S_2__sbox_inst_com_y_inst_n518,
         round_inst_S_2__sbox_inst_com_y_inst_n517,
         round_inst_S_2__sbox_inst_com_y_inst_n516,
         round_inst_S_2__sbox_inst_com_y_inst_n515,
         round_inst_S_2__sbox_inst_com_y_inst_n514,
         round_inst_S_2__sbox_inst_com_y_inst_n513,
         round_inst_S_2__sbox_inst_com_y_inst_n512,
         round_inst_S_2__sbox_inst_com_y_inst_n511,
         round_inst_S_2__sbox_inst_com_y_inst_n510,
         round_inst_S_2__sbox_inst_com_y_inst_n509,
         round_inst_S_2__sbox_inst_com_y_inst_n508,
         round_inst_S_2__sbox_inst_com_y_inst_n507,
         round_inst_S_2__sbox_inst_com_y_inst_n506,
         round_inst_S_2__sbox_inst_com_y_inst_n505,
         round_inst_S_2__sbox_inst_com_y_inst_n504,
         round_inst_S_2__sbox_inst_com_y_inst_n503,
         round_inst_S_2__sbox_inst_com_y_inst_n502,
         round_inst_S_2__sbox_inst_com_y_inst_n501,
         round_inst_S_2__sbox_inst_com_y_inst_n500,
         round_inst_S_2__sbox_inst_com_y_inst_n499,
         round_inst_S_2__sbox_inst_com_y_inst_n498,
         round_inst_S_2__sbox_inst_com_y_inst_n497,
         round_inst_S_2__sbox_inst_com_y_inst_n496,
         round_inst_S_2__sbox_inst_com_y_inst_n495,
         round_inst_S_2__sbox_inst_com_y_inst_n494,
         round_inst_S_2__sbox_inst_com_y_inst_n493,
         round_inst_S_2__sbox_inst_com_y_inst_n492,
         round_inst_S_2__sbox_inst_com_y_inst_n491,
         round_inst_S_2__sbox_inst_com_y_inst_n490,
         round_inst_S_2__sbox_inst_com_y_inst_n489,
         round_inst_S_2__sbox_inst_com_y_inst_n488,
         round_inst_S_2__sbox_inst_com_y_inst_n487,
         round_inst_S_2__sbox_inst_com_y_inst_n486,
         round_inst_S_2__sbox_inst_com_y_inst_n485,
         round_inst_S_2__sbox_inst_com_y_inst_n484,
         round_inst_S_2__sbox_inst_com_y_inst_n483,
         round_inst_S_2__sbox_inst_com_y_inst_n482,
         round_inst_S_2__sbox_inst_com_y_inst_n481,
         round_inst_S_2__sbox_inst_com_y_inst_n480,
         round_inst_S_2__sbox_inst_com_y_inst_n479,
         round_inst_S_2__sbox_inst_com_y_inst_n478,
         round_inst_S_2__sbox_inst_com_y_inst_n477,
         round_inst_S_2__sbox_inst_com_y_inst_n476,
         round_inst_S_2__sbox_inst_com_y_inst_n475,
         round_inst_S_2__sbox_inst_com_y_inst_n474,
         round_inst_S_2__sbox_inst_com_y_inst_n473,
         round_inst_S_2__sbox_inst_com_y_inst_n472,
         round_inst_S_2__sbox_inst_com_y_inst_n471,
         round_inst_S_2__sbox_inst_com_y_inst_n470,
         round_inst_S_2__sbox_inst_com_y_inst_n469,
         round_inst_S_2__sbox_inst_com_y_inst_n468,
         round_inst_S_2__sbox_inst_com_y_inst_n467,
         round_inst_S_2__sbox_inst_com_y_inst_n466,
         round_inst_S_2__sbox_inst_com_y_inst_n465,
         round_inst_S_2__sbox_inst_com_y_inst_n464,
         round_inst_S_2__sbox_inst_com_y_inst_n463,
         round_inst_S_2__sbox_inst_com_y_inst_n462,
         round_inst_S_2__sbox_inst_com_y_inst_n461,
         round_inst_S_2__sbox_inst_com_y_inst_n460,
         round_inst_S_2__sbox_inst_com_y_inst_n459,
         round_inst_S_2__sbox_inst_com_y_inst_n458,
         round_inst_S_2__sbox_inst_com_y_inst_n457,
         round_inst_S_2__sbox_inst_com_y_inst_n456,
         round_inst_S_2__sbox_inst_com_y_inst_n455,
         round_inst_S_2__sbox_inst_com_y_inst_n454,
         round_inst_S_2__sbox_inst_com_y_inst_n453,
         round_inst_S_2__sbox_inst_com_y_inst_n452,
         round_inst_S_2__sbox_inst_com_y_inst_n451,
         round_inst_S_2__sbox_inst_com_y_inst_n450,
         round_inst_S_2__sbox_inst_com_y_inst_n449,
         round_inst_S_2__sbox_inst_com_y_inst_n448,
         round_inst_S_2__sbox_inst_com_y_inst_n447,
         round_inst_S_2__sbox_inst_com_y_inst_n446,
         round_inst_S_2__sbox_inst_com_y_inst_n445,
         round_inst_S_2__sbox_inst_com_y_inst_n444,
         round_inst_S_2__sbox_inst_com_y_inst_n443,
         round_inst_S_2__sbox_inst_com_y_inst_n442,
         round_inst_S_2__sbox_inst_com_y_inst_n441,
         round_inst_S_2__sbox_inst_com_y_inst_n440,
         round_inst_S_2__sbox_inst_com_y_inst_n439,
         round_inst_S_2__sbox_inst_com_y_inst_n438,
         round_inst_S_2__sbox_inst_com_y_inst_n437,
         round_inst_S_2__sbox_inst_com_y_inst_n436,
         round_inst_S_2__sbox_inst_com_y_inst_n435,
         round_inst_S_2__sbox_inst_com_y_inst_n434,
         round_inst_S_2__sbox_inst_com_y_inst_n433,
         round_inst_S_2__sbox_inst_com_y_inst_n432,
         round_inst_S_2__sbox_inst_com_y_inst_n431,
         round_inst_S_2__sbox_inst_com_y_inst_n430,
         round_inst_S_2__sbox_inst_com_y_inst_n429,
         round_inst_S_2__sbox_inst_com_y_inst_n428,
         round_inst_S_2__sbox_inst_com_y_inst_n427,
         round_inst_S_2__sbox_inst_com_y_inst_n426,
         round_inst_S_2__sbox_inst_com_y_inst_n425,
         round_inst_S_2__sbox_inst_com_y_inst_n424,
         round_inst_S_2__sbox_inst_com_y_inst_n423,
         round_inst_S_2__sbox_inst_com_y_inst_n422,
         round_inst_S_2__sbox_inst_com_y_inst_n421,
         round_inst_S_2__sbox_inst_com_y_inst_n420,
         round_inst_S_2__sbox_inst_com_y_inst_n419,
         round_inst_S_2__sbox_inst_com_y_inst_n418,
         round_inst_S_2__sbox_inst_com_y_inst_n417,
         round_inst_S_2__sbox_inst_com_y_inst_n416,
         round_inst_S_2__sbox_inst_com_y_inst_n415,
         round_inst_S_2__sbox_inst_com_y_inst_n414,
         round_inst_S_2__sbox_inst_com_y_inst_n413,
         round_inst_S_2__sbox_inst_com_y_inst_n412,
         round_inst_S_2__sbox_inst_com_y_inst_n411,
         round_inst_S_2__sbox_inst_com_y_inst_n410,
         round_inst_S_2__sbox_inst_com_y_inst_n409,
         round_inst_S_2__sbox_inst_com_y_inst_n408,
         round_inst_S_2__sbox_inst_com_y_inst_n407,
         round_inst_S_2__sbox_inst_com_y_inst_n406,
         round_inst_S_2__sbox_inst_com_y_inst_n405,
         round_inst_S_2__sbox_inst_com_y_inst_n404,
         round_inst_S_2__sbox_inst_com_y_inst_n403,
         round_inst_S_2__sbox_inst_com_y_inst_n402,
         round_inst_S_2__sbox_inst_com_y_inst_n401,
         round_inst_S_2__sbox_inst_com_y_inst_n400,
         round_inst_S_2__sbox_inst_com_y_inst_n399,
         round_inst_S_2__sbox_inst_com_y_inst_n398,
         round_inst_S_2__sbox_inst_com_y_inst_n397,
         round_inst_S_2__sbox_inst_com_y_inst_n396,
         round_inst_S_2__sbox_inst_com_y_inst_n395,
         round_inst_S_2__sbox_inst_com_y_inst_n394,
         round_inst_S_2__sbox_inst_com_y_inst_n393,
         round_inst_S_2__sbox_inst_com_y_inst_n392,
         round_inst_S_2__sbox_inst_com_y_inst_n391,
         round_inst_S_2__sbox_inst_com_y_inst_n390,
         round_inst_S_2__sbox_inst_com_y_inst_n389,
         round_inst_S_2__sbox_inst_com_y_inst_n388,
         round_inst_S_2__sbox_inst_com_y_inst_n387,
         round_inst_S_2__sbox_inst_com_y_inst_n386,
         round_inst_S_2__sbox_inst_com_z_inst_n516,
         round_inst_S_2__sbox_inst_com_z_inst_n515,
         round_inst_S_2__sbox_inst_com_z_inst_n514,
         round_inst_S_2__sbox_inst_com_z_inst_n513,
         round_inst_S_2__sbox_inst_com_z_inst_n512,
         round_inst_S_2__sbox_inst_com_z_inst_n511,
         round_inst_S_2__sbox_inst_com_z_inst_n510,
         round_inst_S_2__sbox_inst_com_z_inst_n509,
         round_inst_S_2__sbox_inst_com_z_inst_n508,
         round_inst_S_2__sbox_inst_com_z_inst_n507,
         round_inst_S_2__sbox_inst_com_z_inst_n506,
         round_inst_S_2__sbox_inst_com_z_inst_n505,
         round_inst_S_2__sbox_inst_com_z_inst_n504,
         round_inst_S_2__sbox_inst_com_z_inst_n503,
         round_inst_S_2__sbox_inst_com_z_inst_n502,
         round_inst_S_2__sbox_inst_com_z_inst_n501,
         round_inst_S_2__sbox_inst_com_z_inst_n500,
         round_inst_S_2__sbox_inst_com_z_inst_n499,
         round_inst_S_2__sbox_inst_com_z_inst_n498,
         round_inst_S_2__sbox_inst_com_z_inst_n497,
         round_inst_S_2__sbox_inst_com_z_inst_n496,
         round_inst_S_2__sbox_inst_com_z_inst_n495,
         round_inst_S_2__sbox_inst_com_z_inst_n494,
         round_inst_S_2__sbox_inst_com_z_inst_n493,
         round_inst_S_2__sbox_inst_com_z_inst_n492,
         round_inst_S_2__sbox_inst_com_z_inst_n491,
         round_inst_S_2__sbox_inst_com_z_inst_n490,
         round_inst_S_2__sbox_inst_com_z_inst_n489,
         round_inst_S_2__sbox_inst_com_z_inst_n488,
         round_inst_S_2__sbox_inst_com_z_inst_n487,
         round_inst_S_2__sbox_inst_com_z_inst_n486,
         round_inst_S_2__sbox_inst_com_z_inst_n485,
         round_inst_S_2__sbox_inst_com_z_inst_n484,
         round_inst_S_2__sbox_inst_com_z_inst_n483,
         round_inst_S_2__sbox_inst_com_z_inst_n482,
         round_inst_S_2__sbox_inst_com_z_inst_n481,
         round_inst_S_2__sbox_inst_com_z_inst_n480,
         round_inst_S_2__sbox_inst_com_z_inst_n479,
         round_inst_S_2__sbox_inst_com_z_inst_n478,
         round_inst_S_2__sbox_inst_com_z_inst_n477,
         round_inst_S_2__sbox_inst_com_z_inst_n476,
         round_inst_S_2__sbox_inst_com_z_inst_n475,
         round_inst_S_2__sbox_inst_com_z_inst_n474,
         round_inst_S_2__sbox_inst_com_z_inst_n473,
         round_inst_S_2__sbox_inst_com_z_inst_n472,
         round_inst_S_2__sbox_inst_com_z_inst_n471,
         round_inst_S_2__sbox_inst_com_z_inst_n470,
         round_inst_S_2__sbox_inst_com_z_inst_n469,
         round_inst_S_2__sbox_inst_com_z_inst_n468,
         round_inst_S_2__sbox_inst_com_z_inst_n467,
         round_inst_S_2__sbox_inst_com_z_inst_n466,
         round_inst_S_2__sbox_inst_com_z_inst_n465,
         round_inst_S_2__sbox_inst_com_z_inst_n464,
         round_inst_S_2__sbox_inst_com_z_inst_n463,
         round_inst_S_2__sbox_inst_com_z_inst_n462,
         round_inst_S_2__sbox_inst_com_z_inst_n461,
         round_inst_S_2__sbox_inst_com_z_inst_n460,
         round_inst_S_2__sbox_inst_com_z_inst_n459,
         round_inst_S_2__sbox_inst_com_z_inst_n458,
         round_inst_S_2__sbox_inst_com_z_inst_n457,
         round_inst_S_2__sbox_inst_com_z_inst_n456,
         round_inst_S_2__sbox_inst_com_z_inst_n455,
         round_inst_S_2__sbox_inst_com_z_inst_n454,
         round_inst_S_2__sbox_inst_com_z_inst_n453,
         round_inst_S_2__sbox_inst_com_z_inst_n452,
         round_inst_S_2__sbox_inst_com_z_inst_n451,
         round_inst_S_2__sbox_inst_com_z_inst_n450,
         round_inst_S_2__sbox_inst_com_z_inst_n449,
         round_inst_S_2__sbox_inst_com_z_inst_n448,
         round_inst_S_2__sbox_inst_com_z_inst_n447,
         round_inst_S_2__sbox_inst_com_z_inst_n446,
         round_inst_S_2__sbox_inst_com_z_inst_n445,
         round_inst_S_2__sbox_inst_com_z_inst_n444,
         round_inst_S_2__sbox_inst_com_z_inst_n443,
         round_inst_S_2__sbox_inst_com_z_inst_n442,
         round_inst_S_2__sbox_inst_com_z_inst_n441,
         round_inst_S_2__sbox_inst_com_z_inst_n440,
         round_inst_S_2__sbox_inst_com_z_inst_n439,
         round_inst_S_2__sbox_inst_com_z_inst_n438,
         round_inst_S_2__sbox_inst_com_z_inst_n437,
         round_inst_S_2__sbox_inst_com_z_inst_n436,
         round_inst_S_2__sbox_inst_com_z_inst_n435,
         round_inst_S_2__sbox_inst_com_z_inst_n434,
         round_inst_S_2__sbox_inst_com_z_inst_n433,
         round_inst_S_2__sbox_inst_com_z_inst_n432,
         round_inst_S_2__sbox_inst_com_z_inst_n431,
         round_inst_S_2__sbox_inst_com_z_inst_n430,
         round_inst_S_2__sbox_inst_com_z_inst_n429,
         round_inst_S_2__sbox_inst_com_z_inst_n428,
         round_inst_S_2__sbox_inst_com_z_inst_n427,
         round_inst_S_2__sbox_inst_com_z_inst_n426,
         round_inst_S_2__sbox_inst_com_z_inst_n425,
         round_inst_S_2__sbox_inst_com_z_inst_n424,
         round_inst_S_2__sbox_inst_com_z_inst_n423,
         round_inst_S_2__sbox_inst_com_z_inst_n422,
         round_inst_S_2__sbox_inst_com_z_inst_n421,
         round_inst_S_2__sbox_inst_com_z_inst_n420,
         round_inst_S_2__sbox_inst_com_z_inst_n419,
         round_inst_S_2__sbox_inst_com_z_inst_n418,
         round_inst_S_2__sbox_inst_com_z_inst_n417,
         round_inst_S_2__sbox_inst_com_z_inst_n416,
         round_inst_S_2__sbox_inst_com_z_inst_n415,
         round_inst_S_2__sbox_inst_com_z_inst_n414,
         round_inst_S_2__sbox_inst_com_z_inst_n413,
         round_inst_S_2__sbox_inst_com_z_inst_n412,
         round_inst_S_2__sbox_inst_com_z_inst_n411,
         round_inst_S_2__sbox_inst_com_z_inst_n410,
         round_inst_S_2__sbox_inst_com_z_inst_n409,
         round_inst_S_2__sbox_inst_com_z_inst_n408,
         round_inst_S_2__sbox_inst_com_z_inst_n407,
         round_inst_S_2__sbox_inst_com_z_inst_n406,
         round_inst_S_2__sbox_inst_com_z_inst_n405,
         round_inst_S_2__sbox_inst_com_z_inst_n404,
         round_inst_S_2__sbox_inst_com_z_inst_n403,
         round_inst_S_2__sbox_inst_com_z_inst_n402,
         round_inst_S_2__sbox_inst_com_z_inst_n401,
         round_inst_S_2__sbox_inst_com_z_inst_n400,
         round_inst_S_2__sbox_inst_com_z_inst_n399,
         round_inst_S_2__sbox_inst_com_z_inst_n398,
         round_inst_S_2__sbox_inst_com_z_inst_n397,
         round_inst_S_2__sbox_inst_com_z_inst_n396,
         round_inst_S_2__sbox_inst_com_z_inst_n395,
         round_inst_S_2__sbox_inst_com_z_inst_n394,
         round_inst_S_2__sbox_inst_com_z_inst_n393,
         round_inst_S_2__sbox_inst_com_z_inst_n392,
         round_inst_S_2__sbox_inst_com_z_inst_n391,
         round_inst_S_2__sbox_inst_com_z_inst_n390,
         round_inst_S_3__sbox_inst_n6, round_inst_S_3__sbox_inst_n5,
         round_inst_S_3__sbox_inst_n4, round_inst_S_3__sbox_inst_n3,
         round_inst_S_3__sbox_inst_n2, round_inst_S_3__sbox_inst_n1,
         round_inst_S_3__sbox_inst_com_w_inst_n532,
         round_inst_S_3__sbox_inst_com_w_inst_n531,
         round_inst_S_3__sbox_inst_com_w_inst_n530,
         round_inst_S_3__sbox_inst_com_w_inst_n529,
         round_inst_S_3__sbox_inst_com_w_inst_n528,
         round_inst_S_3__sbox_inst_com_w_inst_n527,
         round_inst_S_3__sbox_inst_com_w_inst_n526,
         round_inst_S_3__sbox_inst_com_w_inst_n525,
         round_inst_S_3__sbox_inst_com_w_inst_n524,
         round_inst_S_3__sbox_inst_com_w_inst_n523,
         round_inst_S_3__sbox_inst_com_w_inst_n522,
         round_inst_S_3__sbox_inst_com_w_inst_n521,
         round_inst_S_3__sbox_inst_com_w_inst_n520,
         round_inst_S_3__sbox_inst_com_w_inst_n519,
         round_inst_S_3__sbox_inst_com_w_inst_n518,
         round_inst_S_3__sbox_inst_com_w_inst_n517,
         round_inst_S_3__sbox_inst_com_w_inst_n516,
         round_inst_S_3__sbox_inst_com_w_inst_n515,
         round_inst_S_3__sbox_inst_com_w_inst_n514,
         round_inst_S_3__sbox_inst_com_w_inst_n513,
         round_inst_S_3__sbox_inst_com_w_inst_n512,
         round_inst_S_3__sbox_inst_com_w_inst_n511,
         round_inst_S_3__sbox_inst_com_w_inst_n510,
         round_inst_S_3__sbox_inst_com_w_inst_n509,
         round_inst_S_3__sbox_inst_com_w_inst_n508,
         round_inst_S_3__sbox_inst_com_w_inst_n507,
         round_inst_S_3__sbox_inst_com_w_inst_n506,
         round_inst_S_3__sbox_inst_com_w_inst_n505,
         round_inst_S_3__sbox_inst_com_w_inst_n504,
         round_inst_S_3__sbox_inst_com_w_inst_n503,
         round_inst_S_3__sbox_inst_com_w_inst_n502,
         round_inst_S_3__sbox_inst_com_w_inst_n501,
         round_inst_S_3__sbox_inst_com_w_inst_n500,
         round_inst_S_3__sbox_inst_com_w_inst_n499,
         round_inst_S_3__sbox_inst_com_w_inst_n498,
         round_inst_S_3__sbox_inst_com_w_inst_n497,
         round_inst_S_3__sbox_inst_com_w_inst_n496,
         round_inst_S_3__sbox_inst_com_w_inst_n495,
         round_inst_S_3__sbox_inst_com_w_inst_n494,
         round_inst_S_3__sbox_inst_com_w_inst_n493,
         round_inst_S_3__sbox_inst_com_w_inst_n492,
         round_inst_S_3__sbox_inst_com_w_inst_n491,
         round_inst_S_3__sbox_inst_com_w_inst_n490,
         round_inst_S_3__sbox_inst_com_w_inst_n489,
         round_inst_S_3__sbox_inst_com_w_inst_n488,
         round_inst_S_3__sbox_inst_com_w_inst_n487,
         round_inst_S_3__sbox_inst_com_w_inst_n486,
         round_inst_S_3__sbox_inst_com_w_inst_n485,
         round_inst_S_3__sbox_inst_com_w_inst_n484,
         round_inst_S_3__sbox_inst_com_w_inst_n483,
         round_inst_S_3__sbox_inst_com_w_inst_n482,
         round_inst_S_3__sbox_inst_com_w_inst_n481,
         round_inst_S_3__sbox_inst_com_w_inst_n480,
         round_inst_S_3__sbox_inst_com_w_inst_n479,
         round_inst_S_3__sbox_inst_com_w_inst_n478,
         round_inst_S_3__sbox_inst_com_w_inst_n477,
         round_inst_S_3__sbox_inst_com_w_inst_n476,
         round_inst_S_3__sbox_inst_com_w_inst_n475,
         round_inst_S_3__sbox_inst_com_w_inst_n474,
         round_inst_S_3__sbox_inst_com_w_inst_n473,
         round_inst_S_3__sbox_inst_com_w_inst_n472,
         round_inst_S_3__sbox_inst_com_w_inst_n471,
         round_inst_S_3__sbox_inst_com_w_inst_n470,
         round_inst_S_3__sbox_inst_com_w_inst_n469,
         round_inst_S_3__sbox_inst_com_w_inst_n468,
         round_inst_S_3__sbox_inst_com_w_inst_n467,
         round_inst_S_3__sbox_inst_com_w_inst_n466,
         round_inst_S_3__sbox_inst_com_w_inst_n465,
         round_inst_S_3__sbox_inst_com_w_inst_n464,
         round_inst_S_3__sbox_inst_com_w_inst_n463,
         round_inst_S_3__sbox_inst_com_w_inst_n462,
         round_inst_S_3__sbox_inst_com_w_inst_n461,
         round_inst_S_3__sbox_inst_com_w_inst_n460,
         round_inst_S_3__sbox_inst_com_w_inst_n459,
         round_inst_S_3__sbox_inst_com_w_inst_n458,
         round_inst_S_3__sbox_inst_com_w_inst_n457,
         round_inst_S_3__sbox_inst_com_w_inst_n456,
         round_inst_S_3__sbox_inst_com_w_inst_n455,
         round_inst_S_3__sbox_inst_com_w_inst_n454,
         round_inst_S_3__sbox_inst_com_w_inst_n453,
         round_inst_S_3__sbox_inst_com_w_inst_n452,
         round_inst_S_3__sbox_inst_com_w_inst_n451,
         round_inst_S_3__sbox_inst_com_w_inst_n450,
         round_inst_S_3__sbox_inst_com_w_inst_n449,
         round_inst_S_3__sbox_inst_com_w_inst_n448,
         round_inst_S_3__sbox_inst_com_w_inst_n447,
         round_inst_S_3__sbox_inst_com_w_inst_n446,
         round_inst_S_3__sbox_inst_com_w_inst_n445,
         round_inst_S_3__sbox_inst_com_w_inst_n444,
         round_inst_S_3__sbox_inst_com_w_inst_n443,
         round_inst_S_3__sbox_inst_com_w_inst_n442,
         round_inst_S_3__sbox_inst_com_w_inst_n441,
         round_inst_S_3__sbox_inst_com_w_inst_n440,
         round_inst_S_3__sbox_inst_com_w_inst_n439,
         round_inst_S_3__sbox_inst_com_w_inst_n438,
         round_inst_S_3__sbox_inst_com_w_inst_n437,
         round_inst_S_3__sbox_inst_com_w_inst_n436,
         round_inst_S_3__sbox_inst_com_w_inst_n435,
         round_inst_S_3__sbox_inst_com_w_inst_n434,
         round_inst_S_3__sbox_inst_com_w_inst_n433,
         round_inst_S_3__sbox_inst_com_w_inst_n432,
         round_inst_S_3__sbox_inst_com_w_inst_n431,
         round_inst_S_3__sbox_inst_com_w_inst_n430,
         round_inst_S_3__sbox_inst_com_w_inst_n429,
         round_inst_S_3__sbox_inst_com_w_inst_n428,
         round_inst_S_3__sbox_inst_com_w_inst_n427,
         round_inst_S_3__sbox_inst_com_w_inst_n426,
         round_inst_S_3__sbox_inst_com_w_inst_n425,
         round_inst_S_3__sbox_inst_com_w_inst_n424,
         round_inst_S_3__sbox_inst_com_w_inst_n423,
         round_inst_S_3__sbox_inst_com_w_inst_n422,
         round_inst_S_3__sbox_inst_com_w_inst_n421,
         round_inst_S_3__sbox_inst_com_w_inst_n420,
         round_inst_S_3__sbox_inst_com_w_inst_n419,
         round_inst_S_3__sbox_inst_com_w_inst_n418,
         round_inst_S_3__sbox_inst_com_w_inst_n417,
         round_inst_S_3__sbox_inst_com_w_inst_n416,
         round_inst_S_3__sbox_inst_com_w_inst_n415,
         round_inst_S_3__sbox_inst_com_w_inst_n414,
         round_inst_S_3__sbox_inst_com_w_inst_n413,
         round_inst_S_3__sbox_inst_com_w_inst_n412,
         round_inst_S_3__sbox_inst_com_w_inst_n411,
         round_inst_S_3__sbox_inst_com_w_inst_n410,
         round_inst_S_3__sbox_inst_com_w_inst_n409,
         round_inst_S_3__sbox_inst_com_w_inst_n408,
         round_inst_S_3__sbox_inst_com_w_inst_n407,
         round_inst_S_3__sbox_inst_com_w_inst_n406,
         round_inst_S_3__sbox_inst_com_w_inst_n405,
         round_inst_S_3__sbox_inst_com_w_inst_n404,
         round_inst_S_3__sbox_inst_com_w_inst_n403,
         round_inst_S_3__sbox_inst_com_w_inst_n402,
         round_inst_S_3__sbox_inst_com_w_inst_n401,
         round_inst_S_3__sbox_inst_com_w_inst_n400,
         round_inst_S_3__sbox_inst_com_w_inst_n399,
         round_inst_S_3__sbox_inst_com_w_inst_n398,
         round_inst_S_3__sbox_inst_com_w_inst_n397,
         round_inst_S_3__sbox_inst_com_w_inst_n396,
         round_inst_S_3__sbox_inst_com_x_inst_n520,
         round_inst_S_3__sbox_inst_com_x_inst_n519,
         round_inst_S_3__sbox_inst_com_x_inst_n518,
         round_inst_S_3__sbox_inst_com_x_inst_n517,
         round_inst_S_3__sbox_inst_com_x_inst_n516,
         round_inst_S_3__sbox_inst_com_x_inst_n515,
         round_inst_S_3__sbox_inst_com_x_inst_n514,
         round_inst_S_3__sbox_inst_com_x_inst_n513,
         round_inst_S_3__sbox_inst_com_x_inst_n512,
         round_inst_S_3__sbox_inst_com_x_inst_n511,
         round_inst_S_3__sbox_inst_com_x_inst_n510,
         round_inst_S_3__sbox_inst_com_x_inst_n509,
         round_inst_S_3__sbox_inst_com_x_inst_n508,
         round_inst_S_3__sbox_inst_com_x_inst_n507,
         round_inst_S_3__sbox_inst_com_x_inst_n506,
         round_inst_S_3__sbox_inst_com_x_inst_n505,
         round_inst_S_3__sbox_inst_com_x_inst_n504,
         round_inst_S_3__sbox_inst_com_x_inst_n503,
         round_inst_S_3__sbox_inst_com_x_inst_n502,
         round_inst_S_3__sbox_inst_com_x_inst_n501,
         round_inst_S_3__sbox_inst_com_x_inst_n500,
         round_inst_S_3__sbox_inst_com_x_inst_n499,
         round_inst_S_3__sbox_inst_com_x_inst_n498,
         round_inst_S_3__sbox_inst_com_x_inst_n497,
         round_inst_S_3__sbox_inst_com_x_inst_n496,
         round_inst_S_3__sbox_inst_com_x_inst_n495,
         round_inst_S_3__sbox_inst_com_x_inst_n494,
         round_inst_S_3__sbox_inst_com_x_inst_n493,
         round_inst_S_3__sbox_inst_com_x_inst_n492,
         round_inst_S_3__sbox_inst_com_x_inst_n491,
         round_inst_S_3__sbox_inst_com_x_inst_n490,
         round_inst_S_3__sbox_inst_com_x_inst_n489,
         round_inst_S_3__sbox_inst_com_x_inst_n488,
         round_inst_S_3__sbox_inst_com_x_inst_n487,
         round_inst_S_3__sbox_inst_com_x_inst_n486,
         round_inst_S_3__sbox_inst_com_x_inst_n485,
         round_inst_S_3__sbox_inst_com_x_inst_n484,
         round_inst_S_3__sbox_inst_com_x_inst_n483,
         round_inst_S_3__sbox_inst_com_x_inst_n482,
         round_inst_S_3__sbox_inst_com_x_inst_n481,
         round_inst_S_3__sbox_inst_com_x_inst_n480,
         round_inst_S_3__sbox_inst_com_x_inst_n479,
         round_inst_S_3__sbox_inst_com_x_inst_n478,
         round_inst_S_3__sbox_inst_com_x_inst_n477,
         round_inst_S_3__sbox_inst_com_x_inst_n476,
         round_inst_S_3__sbox_inst_com_x_inst_n475,
         round_inst_S_3__sbox_inst_com_x_inst_n474,
         round_inst_S_3__sbox_inst_com_x_inst_n473,
         round_inst_S_3__sbox_inst_com_x_inst_n472,
         round_inst_S_3__sbox_inst_com_x_inst_n471,
         round_inst_S_3__sbox_inst_com_x_inst_n470,
         round_inst_S_3__sbox_inst_com_x_inst_n469,
         round_inst_S_3__sbox_inst_com_x_inst_n468,
         round_inst_S_3__sbox_inst_com_x_inst_n467,
         round_inst_S_3__sbox_inst_com_x_inst_n466,
         round_inst_S_3__sbox_inst_com_x_inst_n465,
         round_inst_S_3__sbox_inst_com_x_inst_n464,
         round_inst_S_3__sbox_inst_com_x_inst_n463,
         round_inst_S_3__sbox_inst_com_x_inst_n462,
         round_inst_S_3__sbox_inst_com_x_inst_n461,
         round_inst_S_3__sbox_inst_com_x_inst_n460,
         round_inst_S_3__sbox_inst_com_x_inst_n459,
         round_inst_S_3__sbox_inst_com_x_inst_n458,
         round_inst_S_3__sbox_inst_com_x_inst_n457,
         round_inst_S_3__sbox_inst_com_x_inst_n456,
         round_inst_S_3__sbox_inst_com_x_inst_n455,
         round_inst_S_3__sbox_inst_com_x_inst_n454,
         round_inst_S_3__sbox_inst_com_x_inst_n453,
         round_inst_S_3__sbox_inst_com_x_inst_n452,
         round_inst_S_3__sbox_inst_com_x_inst_n451,
         round_inst_S_3__sbox_inst_com_x_inst_n450,
         round_inst_S_3__sbox_inst_com_x_inst_n449,
         round_inst_S_3__sbox_inst_com_x_inst_n448,
         round_inst_S_3__sbox_inst_com_x_inst_n447,
         round_inst_S_3__sbox_inst_com_x_inst_n446,
         round_inst_S_3__sbox_inst_com_x_inst_n445,
         round_inst_S_3__sbox_inst_com_x_inst_n444,
         round_inst_S_3__sbox_inst_com_x_inst_n443,
         round_inst_S_3__sbox_inst_com_x_inst_n442,
         round_inst_S_3__sbox_inst_com_x_inst_n441,
         round_inst_S_3__sbox_inst_com_x_inst_n440,
         round_inst_S_3__sbox_inst_com_x_inst_n439,
         round_inst_S_3__sbox_inst_com_x_inst_n438,
         round_inst_S_3__sbox_inst_com_x_inst_n437,
         round_inst_S_3__sbox_inst_com_x_inst_n436,
         round_inst_S_3__sbox_inst_com_x_inst_n435,
         round_inst_S_3__sbox_inst_com_x_inst_n434,
         round_inst_S_3__sbox_inst_com_x_inst_n433,
         round_inst_S_3__sbox_inst_com_x_inst_n432,
         round_inst_S_3__sbox_inst_com_x_inst_n431,
         round_inst_S_3__sbox_inst_com_x_inst_n430,
         round_inst_S_3__sbox_inst_com_x_inst_n429,
         round_inst_S_3__sbox_inst_com_x_inst_n428,
         round_inst_S_3__sbox_inst_com_x_inst_n427,
         round_inst_S_3__sbox_inst_com_x_inst_n426,
         round_inst_S_3__sbox_inst_com_x_inst_n425,
         round_inst_S_3__sbox_inst_com_x_inst_n424,
         round_inst_S_3__sbox_inst_com_x_inst_n423,
         round_inst_S_3__sbox_inst_com_x_inst_n422,
         round_inst_S_3__sbox_inst_com_x_inst_n421,
         round_inst_S_3__sbox_inst_com_x_inst_n420,
         round_inst_S_3__sbox_inst_com_x_inst_n419,
         round_inst_S_3__sbox_inst_com_x_inst_n418,
         round_inst_S_3__sbox_inst_com_x_inst_n417,
         round_inst_S_3__sbox_inst_com_x_inst_n416,
         round_inst_S_3__sbox_inst_com_x_inst_n415,
         round_inst_S_3__sbox_inst_com_x_inst_n414,
         round_inst_S_3__sbox_inst_com_x_inst_n413,
         round_inst_S_3__sbox_inst_com_x_inst_n412,
         round_inst_S_3__sbox_inst_com_x_inst_n411,
         round_inst_S_3__sbox_inst_com_x_inst_n410,
         round_inst_S_3__sbox_inst_com_x_inst_n409,
         round_inst_S_3__sbox_inst_com_x_inst_n408,
         round_inst_S_3__sbox_inst_com_x_inst_n407,
         round_inst_S_3__sbox_inst_com_x_inst_n406,
         round_inst_S_3__sbox_inst_com_x_inst_n405,
         round_inst_S_3__sbox_inst_com_x_inst_n404,
         round_inst_S_3__sbox_inst_com_x_inst_n403,
         round_inst_S_3__sbox_inst_com_x_inst_n402,
         round_inst_S_3__sbox_inst_com_x_inst_n401,
         round_inst_S_3__sbox_inst_com_x_inst_n400,
         round_inst_S_3__sbox_inst_com_x_inst_n399,
         round_inst_S_3__sbox_inst_com_x_inst_n398,
         round_inst_S_3__sbox_inst_com_x_inst_n397,
         round_inst_S_3__sbox_inst_com_x_inst_n396,
         round_inst_S_3__sbox_inst_com_x_inst_n395,
         round_inst_S_3__sbox_inst_com_x_inst_n394,
         round_inst_S_3__sbox_inst_com_x_inst_n393,
         round_inst_S_3__sbox_inst_com_x_inst_n392,
         round_inst_S_3__sbox_inst_com_x_inst_n391,
         round_inst_S_3__sbox_inst_com_x_inst_n390,
         round_inst_S_3__sbox_inst_com_x_inst_n389,
         round_inst_S_3__sbox_inst_com_x_inst_n388,
         round_inst_S_3__sbox_inst_com_x_inst_n387,
         round_inst_S_3__sbox_inst_com_x_inst_n386,
         round_inst_S_3__sbox_inst_com_x_inst_n385,
         round_inst_S_3__sbox_inst_com_x_inst_n384,
         round_inst_S_3__sbox_inst_com_x_inst_n383,
         round_inst_S_3__sbox_inst_com_x_inst_n382,
         round_inst_S_3__sbox_inst_com_x_inst_n381,
         round_inst_S_3__sbox_inst_com_y_inst_n517,
         round_inst_S_3__sbox_inst_com_y_inst_n516,
         round_inst_S_3__sbox_inst_com_y_inst_n515,
         round_inst_S_3__sbox_inst_com_y_inst_n514,
         round_inst_S_3__sbox_inst_com_y_inst_n513,
         round_inst_S_3__sbox_inst_com_y_inst_n512,
         round_inst_S_3__sbox_inst_com_y_inst_n511,
         round_inst_S_3__sbox_inst_com_y_inst_n510,
         round_inst_S_3__sbox_inst_com_y_inst_n509,
         round_inst_S_3__sbox_inst_com_y_inst_n508,
         round_inst_S_3__sbox_inst_com_y_inst_n507,
         round_inst_S_3__sbox_inst_com_y_inst_n506,
         round_inst_S_3__sbox_inst_com_y_inst_n505,
         round_inst_S_3__sbox_inst_com_y_inst_n504,
         round_inst_S_3__sbox_inst_com_y_inst_n503,
         round_inst_S_3__sbox_inst_com_y_inst_n502,
         round_inst_S_3__sbox_inst_com_y_inst_n501,
         round_inst_S_3__sbox_inst_com_y_inst_n500,
         round_inst_S_3__sbox_inst_com_y_inst_n499,
         round_inst_S_3__sbox_inst_com_y_inst_n498,
         round_inst_S_3__sbox_inst_com_y_inst_n497,
         round_inst_S_3__sbox_inst_com_y_inst_n496,
         round_inst_S_3__sbox_inst_com_y_inst_n495,
         round_inst_S_3__sbox_inst_com_y_inst_n494,
         round_inst_S_3__sbox_inst_com_y_inst_n493,
         round_inst_S_3__sbox_inst_com_y_inst_n492,
         round_inst_S_3__sbox_inst_com_y_inst_n491,
         round_inst_S_3__sbox_inst_com_y_inst_n490,
         round_inst_S_3__sbox_inst_com_y_inst_n489,
         round_inst_S_3__sbox_inst_com_y_inst_n488,
         round_inst_S_3__sbox_inst_com_y_inst_n487,
         round_inst_S_3__sbox_inst_com_y_inst_n486,
         round_inst_S_3__sbox_inst_com_y_inst_n485,
         round_inst_S_3__sbox_inst_com_y_inst_n484,
         round_inst_S_3__sbox_inst_com_y_inst_n483,
         round_inst_S_3__sbox_inst_com_y_inst_n482,
         round_inst_S_3__sbox_inst_com_y_inst_n481,
         round_inst_S_3__sbox_inst_com_y_inst_n480,
         round_inst_S_3__sbox_inst_com_y_inst_n479,
         round_inst_S_3__sbox_inst_com_y_inst_n478,
         round_inst_S_3__sbox_inst_com_y_inst_n477,
         round_inst_S_3__sbox_inst_com_y_inst_n476,
         round_inst_S_3__sbox_inst_com_y_inst_n475,
         round_inst_S_3__sbox_inst_com_y_inst_n474,
         round_inst_S_3__sbox_inst_com_y_inst_n473,
         round_inst_S_3__sbox_inst_com_y_inst_n472,
         round_inst_S_3__sbox_inst_com_y_inst_n471,
         round_inst_S_3__sbox_inst_com_y_inst_n470,
         round_inst_S_3__sbox_inst_com_y_inst_n469,
         round_inst_S_3__sbox_inst_com_y_inst_n468,
         round_inst_S_3__sbox_inst_com_y_inst_n467,
         round_inst_S_3__sbox_inst_com_y_inst_n466,
         round_inst_S_3__sbox_inst_com_y_inst_n465,
         round_inst_S_3__sbox_inst_com_y_inst_n464,
         round_inst_S_3__sbox_inst_com_y_inst_n463,
         round_inst_S_3__sbox_inst_com_y_inst_n462,
         round_inst_S_3__sbox_inst_com_y_inst_n461,
         round_inst_S_3__sbox_inst_com_y_inst_n460,
         round_inst_S_3__sbox_inst_com_y_inst_n459,
         round_inst_S_3__sbox_inst_com_y_inst_n458,
         round_inst_S_3__sbox_inst_com_y_inst_n457,
         round_inst_S_3__sbox_inst_com_y_inst_n456,
         round_inst_S_3__sbox_inst_com_y_inst_n455,
         round_inst_S_3__sbox_inst_com_y_inst_n454,
         round_inst_S_3__sbox_inst_com_y_inst_n453,
         round_inst_S_3__sbox_inst_com_y_inst_n452,
         round_inst_S_3__sbox_inst_com_y_inst_n451,
         round_inst_S_3__sbox_inst_com_y_inst_n450,
         round_inst_S_3__sbox_inst_com_y_inst_n449,
         round_inst_S_3__sbox_inst_com_y_inst_n448,
         round_inst_S_3__sbox_inst_com_y_inst_n447,
         round_inst_S_3__sbox_inst_com_y_inst_n446,
         round_inst_S_3__sbox_inst_com_y_inst_n445,
         round_inst_S_3__sbox_inst_com_y_inst_n444,
         round_inst_S_3__sbox_inst_com_y_inst_n443,
         round_inst_S_3__sbox_inst_com_y_inst_n442,
         round_inst_S_3__sbox_inst_com_y_inst_n441,
         round_inst_S_3__sbox_inst_com_y_inst_n440,
         round_inst_S_3__sbox_inst_com_y_inst_n439,
         round_inst_S_3__sbox_inst_com_y_inst_n438,
         round_inst_S_3__sbox_inst_com_y_inst_n437,
         round_inst_S_3__sbox_inst_com_y_inst_n436,
         round_inst_S_3__sbox_inst_com_y_inst_n435,
         round_inst_S_3__sbox_inst_com_y_inst_n434,
         round_inst_S_3__sbox_inst_com_y_inst_n433,
         round_inst_S_3__sbox_inst_com_y_inst_n432,
         round_inst_S_3__sbox_inst_com_y_inst_n431,
         round_inst_S_3__sbox_inst_com_y_inst_n430,
         round_inst_S_3__sbox_inst_com_y_inst_n429,
         round_inst_S_3__sbox_inst_com_y_inst_n428,
         round_inst_S_3__sbox_inst_com_y_inst_n427,
         round_inst_S_3__sbox_inst_com_y_inst_n426,
         round_inst_S_3__sbox_inst_com_y_inst_n425,
         round_inst_S_3__sbox_inst_com_y_inst_n424,
         round_inst_S_3__sbox_inst_com_y_inst_n423,
         round_inst_S_3__sbox_inst_com_y_inst_n422,
         round_inst_S_3__sbox_inst_com_y_inst_n421,
         round_inst_S_3__sbox_inst_com_y_inst_n420,
         round_inst_S_3__sbox_inst_com_y_inst_n419,
         round_inst_S_3__sbox_inst_com_y_inst_n418,
         round_inst_S_3__sbox_inst_com_y_inst_n417,
         round_inst_S_3__sbox_inst_com_y_inst_n416,
         round_inst_S_3__sbox_inst_com_y_inst_n415,
         round_inst_S_3__sbox_inst_com_y_inst_n414,
         round_inst_S_3__sbox_inst_com_y_inst_n413,
         round_inst_S_3__sbox_inst_com_y_inst_n412,
         round_inst_S_3__sbox_inst_com_y_inst_n411,
         round_inst_S_3__sbox_inst_com_y_inst_n410,
         round_inst_S_3__sbox_inst_com_y_inst_n409,
         round_inst_S_3__sbox_inst_com_y_inst_n408,
         round_inst_S_3__sbox_inst_com_y_inst_n407,
         round_inst_S_3__sbox_inst_com_y_inst_n406,
         round_inst_S_3__sbox_inst_com_y_inst_n405,
         round_inst_S_3__sbox_inst_com_y_inst_n404,
         round_inst_S_3__sbox_inst_com_y_inst_n403,
         round_inst_S_3__sbox_inst_com_y_inst_n402,
         round_inst_S_3__sbox_inst_com_y_inst_n401,
         round_inst_S_3__sbox_inst_com_y_inst_n400,
         round_inst_S_3__sbox_inst_com_y_inst_n399,
         round_inst_S_3__sbox_inst_com_y_inst_n398,
         round_inst_S_3__sbox_inst_com_y_inst_n397,
         round_inst_S_3__sbox_inst_com_y_inst_n396,
         round_inst_S_3__sbox_inst_com_y_inst_n395,
         round_inst_S_3__sbox_inst_com_y_inst_n394,
         round_inst_S_3__sbox_inst_com_y_inst_n393,
         round_inst_S_3__sbox_inst_com_y_inst_n392,
         round_inst_S_3__sbox_inst_com_y_inst_n391,
         round_inst_S_3__sbox_inst_com_y_inst_n390,
         round_inst_S_3__sbox_inst_com_y_inst_n389,
         round_inst_S_3__sbox_inst_com_y_inst_n388,
         round_inst_S_3__sbox_inst_com_y_inst_n387,
         round_inst_S_3__sbox_inst_com_y_inst_n386,
         round_inst_S_3__sbox_inst_com_z_inst_n523,
         round_inst_S_3__sbox_inst_com_z_inst_n522,
         round_inst_S_3__sbox_inst_com_z_inst_n521,
         round_inst_S_3__sbox_inst_com_z_inst_n520,
         round_inst_S_3__sbox_inst_com_z_inst_n519,
         round_inst_S_3__sbox_inst_com_z_inst_n518,
         round_inst_S_3__sbox_inst_com_z_inst_n517,
         round_inst_S_3__sbox_inst_com_z_inst_n516,
         round_inst_S_3__sbox_inst_com_z_inst_n515,
         round_inst_S_3__sbox_inst_com_z_inst_n514,
         round_inst_S_3__sbox_inst_com_z_inst_n513,
         round_inst_S_3__sbox_inst_com_z_inst_n512,
         round_inst_S_3__sbox_inst_com_z_inst_n511,
         round_inst_S_3__sbox_inst_com_z_inst_n510,
         round_inst_S_3__sbox_inst_com_z_inst_n509,
         round_inst_S_3__sbox_inst_com_z_inst_n508,
         round_inst_S_3__sbox_inst_com_z_inst_n507,
         round_inst_S_3__sbox_inst_com_z_inst_n506,
         round_inst_S_3__sbox_inst_com_z_inst_n505,
         round_inst_S_3__sbox_inst_com_z_inst_n504,
         round_inst_S_3__sbox_inst_com_z_inst_n503,
         round_inst_S_3__sbox_inst_com_z_inst_n502,
         round_inst_S_3__sbox_inst_com_z_inst_n501,
         round_inst_S_3__sbox_inst_com_z_inst_n500,
         round_inst_S_3__sbox_inst_com_z_inst_n499,
         round_inst_S_3__sbox_inst_com_z_inst_n498,
         round_inst_S_3__sbox_inst_com_z_inst_n497,
         round_inst_S_3__sbox_inst_com_z_inst_n496,
         round_inst_S_3__sbox_inst_com_z_inst_n495,
         round_inst_S_3__sbox_inst_com_z_inst_n494,
         round_inst_S_3__sbox_inst_com_z_inst_n493,
         round_inst_S_3__sbox_inst_com_z_inst_n492,
         round_inst_S_3__sbox_inst_com_z_inst_n491,
         round_inst_S_3__sbox_inst_com_z_inst_n490,
         round_inst_S_3__sbox_inst_com_z_inst_n489,
         round_inst_S_3__sbox_inst_com_z_inst_n488,
         round_inst_S_3__sbox_inst_com_z_inst_n487,
         round_inst_S_3__sbox_inst_com_z_inst_n486,
         round_inst_S_3__sbox_inst_com_z_inst_n485,
         round_inst_S_3__sbox_inst_com_z_inst_n484,
         round_inst_S_3__sbox_inst_com_z_inst_n483,
         round_inst_S_3__sbox_inst_com_z_inst_n482,
         round_inst_S_3__sbox_inst_com_z_inst_n481,
         round_inst_S_3__sbox_inst_com_z_inst_n480,
         round_inst_S_3__sbox_inst_com_z_inst_n479,
         round_inst_S_3__sbox_inst_com_z_inst_n478,
         round_inst_S_3__sbox_inst_com_z_inst_n477,
         round_inst_S_3__sbox_inst_com_z_inst_n476,
         round_inst_S_3__sbox_inst_com_z_inst_n475,
         round_inst_S_3__sbox_inst_com_z_inst_n474,
         round_inst_S_3__sbox_inst_com_z_inst_n473,
         round_inst_S_3__sbox_inst_com_z_inst_n472,
         round_inst_S_3__sbox_inst_com_z_inst_n471,
         round_inst_S_3__sbox_inst_com_z_inst_n470,
         round_inst_S_3__sbox_inst_com_z_inst_n469,
         round_inst_S_3__sbox_inst_com_z_inst_n468,
         round_inst_S_3__sbox_inst_com_z_inst_n467,
         round_inst_S_3__sbox_inst_com_z_inst_n466,
         round_inst_S_3__sbox_inst_com_z_inst_n465,
         round_inst_S_3__sbox_inst_com_z_inst_n464,
         round_inst_S_3__sbox_inst_com_z_inst_n463,
         round_inst_S_3__sbox_inst_com_z_inst_n462,
         round_inst_S_3__sbox_inst_com_z_inst_n461,
         round_inst_S_3__sbox_inst_com_z_inst_n460,
         round_inst_S_3__sbox_inst_com_z_inst_n459,
         round_inst_S_3__sbox_inst_com_z_inst_n458,
         round_inst_S_3__sbox_inst_com_z_inst_n457,
         round_inst_S_3__sbox_inst_com_z_inst_n456,
         round_inst_S_3__sbox_inst_com_z_inst_n455,
         round_inst_S_3__sbox_inst_com_z_inst_n454,
         round_inst_S_3__sbox_inst_com_z_inst_n453,
         round_inst_S_3__sbox_inst_com_z_inst_n452,
         round_inst_S_3__sbox_inst_com_z_inst_n451,
         round_inst_S_3__sbox_inst_com_z_inst_n450,
         round_inst_S_3__sbox_inst_com_z_inst_n449,
         round_inst_S_3__sbox_inst_com_z_inst_n448,
         round_inst_S_3__sbox_inst_com_z_inst_n447,
         round_inst_S_3__sbox_inst_com_z_inst_n446,
         round_inst_S_3__sbox_inst_com_z_inst_n445,
         round_inst_S_3__sbox_inst_com_z_inst_n444,
         round_inst_S_3__sbox_inst_com_z_inst_n443,
         round_inst_S_3__sbox_inst_com_z_inst_n442,
         round_inst_S_3__sbox_inst_com_z_inst_n441,
         round_inst_S_3__sbox_inst_com_z_inst_n440,
         round_inst_S_3__sbox_inst_com_z_inst_n439,
         round_inst_S_3__sbox_inst_com_z_inst_n438,
         round_inst_S_3__sbox_inst_com_z_inst_n437,
         round_inst_S_3__sbox_inst_com_z_inst_n436,
         round_inst_S_3__sbox_inst_com_z_inst_n435,
         round_inst_S_3__sbox_inst_com_z_inst_n434,
         round_inst_S_3__sbox_inst_com_z_inst_n433,
         round_inst_S_3__sbox_inst_com_z_inst_n432,
         round_inst_S_3__sbox_inst_com_z_inst_n431,
         round_inst_S_3__sbox_inst_com_z_inst_n430,
         round_inst_S_3__sbox_inst_com_z_inst_n429,
         round_inst_S_3__sbox_inst_com_z_inst_n428,
         round_inst_S_3__sbox_inst_com_z_inst_n427,
         round_inst_S_3__sbox_inst_com_z_inst_n426,
         round_inst_S_3__sbox_inst_com_z_inst_n425,
         round_inst_S_3__sbox_inst_com_z_inst_n424,
         round_inst_S_3__sbox_inst_com_z_inst_n423,
         round_inst_S_3__sbox_inst_com_z_inst_n422,
         round_inst_S_3__sbox_inst_com_z_inst_n421,
         round_inst_S_3__sbox_inst_com_z_inst_n420,
         round_inst_S_3__sbox_inst_com_z_inst_n419,
         round_inst_S_3__sbox_inst_com_z_inst_n418,
         round_inst_S_3__sbox_inst_com_z_inst_n417,
         round_inst_S_3__sbox_inst_com_z_inst_n416,
         round_inst_S_3__sbox_inst_com_z_inst_n415,
         round_inst_S_3__sbox_inst_com_z_inst_n414,
         round_inst_S_3__sbox_inst_com_z_inst_n413,
         round_inst_S_3__sbox_inst_com_z_inst_n412,
         round_inst_S_3__sbox_inst_com_z_inst_n411,
         round_inst_S_3__sbox_inst_com_z_inst_n410,
         round_inst_S_3__sbox_inst_com_z_inst_n409,
         round_inst_S_3__sbox_inst_com_z_inst_n408,
         round_inst_S_3__sbox_inst_com_z_inst_n407,
         round_inst_S_3__sbox_inst_com_z_inst_n406,
         round_inst_S_3__sbox_inst_com_z_inst_n405,
         round_inst_S_3__sbox_inst_com_z_inst_n404,
         round_inst_S_3__sbox_inst_com_z_inst_n403,
         round_inst_S_3__sbox_inst_com_z_inst_n402,
         round_inst_S_3__sbox_inst_com_z_inst_n401,
         round_inst_S_3__sbox_inst_com_z_inst_n400,
         round_inst_S_3__sbox_inst_com_z_inst_n399,
         round_inst_S_3__sbox_inst_com_z_inst_n398,
         round_inst_S_3__sbox_inst_com_z_inst_n397,
         round_inst_S_3__sbox_inst_com_z_inst_n396,
         round_inst_S_3__sbox_inst_com_z_inst_n395,
         round_inst_S_3__sbox_inst_com_z_inst_n394,
         round_inst_S_3__sbox_inst_com_z_inst_n393,
         round_inst_S_3__sbox_inst_com_z_inst_n392,
         round_inst_S_3__sbox_inst_com_z_inst_n391,
         round_inst_S_4__sbox_inst_n6, round_inst_S_4__sbox_inst_n5,
         round_inst_S_4__sbox_inst_n4, round_inst_S_4__sbox_inst_n3,
         round_inst_S_4__sbox_inst_n2, round_inst_S_4__sbox_inst_n1,
         round_inst_S_4__sbox_inst_com_w_inst_n532,
         round_inst_S_4__sbox_inst_com_w_inst_n531,
         round_inst_S_4__sbox_inst_com_w_inst_n530,
         round_inst_S_4__sbox_inst_com_w_inst_n529,
         round_inst_S_4__sbox_inst_com_w_inst_n528,
         round_inst_S_4__sbox_inst_com_w_inst_n527,
         round_inst_S_4__sbox_inst_com_w_inst_n526,
         round_inst_S_4__sbox_inst_com_w_inst_n525,
         round_inst_S_4__sbox_inst_com_w_inst_n524,
         round_inst_S_4__sbox_inst_com_w_inst_n523,
         round_inst_S_4__sbox_inst_com_w_inst_n522,
         round_inst_S_4__sbox_inst_com_w_inst_n521,
         round_inst_S_4__sbox_inst_com_w_inst_n520,
         round_inst_S_4__sbox_inst_com_w_inst_n519,
         round_inst_S_4__sbox_inst_com_w_inst_n518,
         round_inst_S_4__sbox_inst_com_w_inst_n517,
         round_inst_S_4__sbox_inst_com_w_inst_n516,
         round_inst_S_4__sbox_inst_com_w_inst_n515,
         round_inst_S_4__sbox_inst_com_w_inst_n514,
         round_inst_S_4__sbox_inst_com_w_inst_n513,
         round_inst_S_4__sbox_inst_com_w_inst_n512,
         round_inst_S_4__sbox_inst_com_w_inst_n511,
         round_inst_S_4__sbox_inst_com_w_inst_n510,
         round_inst_S_4__sbox_inst_com_w_inst_n509,
         round_inst_S_4__sbox_inst_com_w_inst_n508,
         round_inst_S_4__sbox_inst_com_w_inst_n507,
         round_inst_S_4__sbox_inst_com_w_inst_n506,
         round_inst_S_4__sbox_inst_com_w_inst_n505,
         round_inst_S_4__sbox_inst_com_w_inst_n504,
         round_inst_S_4__sbox_inst_com_w_inst_n503,
         round_inst_S_4__sbox_inst_com_w_inst_n502,
         round_inst_S_4__sbox_inst_com_w_inst_n501,
         round_inst_S_4__sbox_inst_com_w_inst_n500,
         round_inst_S_4__sbox_inst_com_w_inst_n499,
         round_inst_S_4__sbox_inst_com_w_inst_n498,
         round_inst_S_4__sbox_inst_com_w_inst_n497,
         round_inst_S_4__sbox_inst_com_w_inst_n496,
         round_inst_S_4__sbox_inst_com_w_inst_n495,
         round_inst_S_4__sbox_inst_com_w_inst_n494,
         round_inst_S_4__sbox_inst_com_w_inst_n493,
         round_inst_S_4__sbox_inst_com_w_inst_n492,
         round_inst_S_4__sbox_inst_com_w_inst_n491,
         round_inst_S_4__sbox_inst_com_w_inst_n490,
         round_inst_S_4__sbox_inst_com_w_inst_n489,
         round_inst_S_4__sbox_inst_com_w_inst_n488,
         round_inst_S_4__sbox_inst_com_w_inst_n487,
         round_inst_S_4__sbox_inst_com_w_inst_n486,
         round_inst_S_4__sbox_inst_com_w_inst_n485,
         round_inst_S_4__sbox_inst_com_w_inst_n484,
         round_inst_S_4__sbox_inst_com_w_inst_n483,
         round_inst_S_4__sbox_inst_com_w_inst_n482,
         round_inst_S_4__sbox_inst_com_w_inst_n481,
         round_inst_S_4__sbox_inst_com_w_inst_n480,
         round_inst_S_4__sbox_inst_com_w_inst_n479,
         round_inst_S_4__sbox_inst_com_w_inst_n478,
         round_inst_S_4__sbox_inst_com_w_inst_n477,
         round_inst_S_4__sbox_inst_com_w_inst_n476,
         round_inst_S_4__sbox_inst_com_w_inst_n475,
         round_inst_S_4__sbox_inst_com_w_inst_n474,
         round_inst_S_4__sbox_inst_com_w_inst_n473,
         round_inst_S_4__sbox_inst_com_w_inst_n472,
         round_inst_S_4__sbox_inst_com_w_inst_n471,
         round_inst_S_4__sbox_inst_com_w_inst_n470,
         round_inst_S_4__sbox_inst_com_w_inst_n469,
         round_inst_S_4__sbox_inst_com_w_inst_n468,
         round_inst_S_4__sbox_inst_com_w_inst_n467,
         round_inst_S_4__sbox_inst_com_w_inst_n466,
         round_inst_S_4__sbox_inst_com_w_inst_n465,
         round_inst_S_4__sbox_inst_com_w_inst_n464,
         round_inst_S_4__sbox_inst_com_w_inst_n463,
         round_inst_S_4__sbox_inst_com_w_inst_n462,
         round_inst_S_4__sbox_inst_com_w_inst_n461,
         round_inst_S_4__sbox_inst_com_w_inst_n460,
         round_inst_S_4__sbox_inst_com_w_inst_n459,
         round_inst_S_4__sbox_inst_com_w_inst_n458,
         round_inst_S_4__sbox_inst_com_w_inst_n457,
         round_inst_S_4__sbox_inst_com_w_inst_n456,
         round_inst_S_4__sbox_inst_com_w_inst_n455,
         round_inst_S_4__sbox_inst_com_w_inst_n454,
         round_inst_S_4__sbox_inst_com_w_inst_n453,
         round_inst_S_4__sbox_inst_com_w_inst_n452,
         round_inst_S_4__sbox_inst_com_w_inst_n451,
         round_inst_S_4__sbox_inst_com_w_inst_n450,
         round_inst_S_4__sbox_inst_com_w_inst_n449,
         round_inst_S_4__sbox_inst_com_w_inst_n448,
         round_inst_S_4__sbox_inst_com_w_inst_n447,
         round_inst_S_4__sbox_inst_com_w_inst_n446,
         round_inst_S_4__sbox_inst_com_w_inst_n445,
         round_inst_S_4__sbox_inst_com_w_inst_n444,
         round_inst_S_4__sbox_inst_com_w_inst_n443,
         round_inst_S_4__sbox_inst_com_w_inst_n442,
         round_inst_S_4__sbox_inst_com_w_inst_n441,
         round_inst_S_4__sbox_inst_com_w_inst_n440,
         round_inst_S_4__sbox_inst_com_w_inst_n439,
         round_inst_S_4__sbox_inst_com_w_inst_n438,
         round_inst_S_4__sbox_inst_com_w_inst_n437,
         round_inst_S_4__sbox_inst_com_w_inst_n436,
         round_inst_S_4__sbox_inst_com_w_inst_n435,
         round_inst_S_4__sbox_inst_com_w_inst_n434,
         round_inst_S_4__sbox_inst_com_w_inst_n433,
         round_inst_S_4__sbox_inst_com_w_inst_n432,
         round_inst_S_4__sbox_inst_com_w_inst_n431,
         round_inst_S_4__sbox_inst_com_w_inst_n430,
         round_inst_S_4__sbox_inst_com_w_inst_n429,
         round_inst_S_4__sbox_inst_com_w_inst_n428,
         round_inst_S_4__sbox_inst_com_w_inst_n427,
         round_inst_S_4__sbox_inst_com_w_inst_n426,
         round_inst_S_4__sbox_inst_com_w_inst_n425,
         round_inst_S_4__sbox_inst_com_w_inst_n424,
         round_inst_S_4__sbox_inst_com_w_inst_n423,
         round_inst_S_4__sbox_inst_com_w_inst_n422,
         round_inst_S_4__sbox_inst_com_w_inst_n421,
         round_inst_S_4__sbox_inst_com_w_inst_n420,
         round_inst_S_4__sbox_inst_com_w_inst_n419,
         round_inst_S_4__sbox_inst_com_w_inst_n418,
         round_inst_S_4__sbox_inst_com_w_inst_n417,
         round_inst_S_4__sbox_inst_com_w_inst_n416,
         round_inst_S_4__sbox_inst_com_w_inst_n415,
         round_inst_S_4__sbox_inst_com_w_inst_n414,
         round_inst_S_4__sbox_inst_com_w_inst_n413,
         round_inst_S_4__sbox_inst_com_w_inst_n412,
         round_inst_S_4__sbox_inst_com_w_inst_n411,
         round_inst_S_4__sbox_inst_com_w_inst_n410,
         round_inst_S_4__sbox_inst_com_w_inst_n409,
         round_inst_S_4__sbox_inst_com_w_inst_n408,
         round_inst_S_4__sbox_inst_com_w_inst_n407,
         round_inst_S_4__sbox_inst_com_w_inst_n406,
         round_inst_S_4__sbox_inst_com_w_inst_n405,
         round_inst_S_4__sbox_inst_com_w_inst_n404,
         round_inst_S_4__sbox_inst_com_w_inst_n403,
         round_inst_S_4__sbox_inst_com_w_inst_n402,
         round_inst_S_4__sbox_inst_com_w_inst_n401,
         round_inst_S_4__sbox_inst_com_w_inst_n400,
         round_inst_S_4__sbox_inst_com_w_inst_n399,
         round_inst_S_4__sbox_inst_com_w_inst_n398,
         round_inst_S_4__sbox_inst_com_w_inst_n397,
         round_inst_S_4__sbox_inst_com_w_inst_n396,
         round_inst_S_4__sbox_inst_com_x_inst_n511,
         round_inst_S_4__sbox_inst_com_x_inst_n510,
         round_inst_S_4__sbox_inst_com_x_inst_n509,
         round_inst_S_4__sbox_inst_com_x_inst_n508,
         round_inst_S_4__sbox_inst_com_x_inst_n507,
         round_inst_S_4__sbox_inst_com_x_inst_n506,
         round_inst_S_4__sbox_inst_com_x_inst_n505,
         round_inst_S_4__sbox_inst_com_x_inst_n504,
         round_inst_S_4__sbox_inst_com_x_inst_n503,
         round_inst_S_4__sbox_inst_com_x_inst_n502,
         round_inst_S_4__sbox_inst_com_x_inst_n501,
         round_inst_S_4__sbox_inst_com_x_inst_n500,
         round_inst_S_4__sbox_inst_com_x_inst_n499,
         round_inst_S_4__sbox_inst_com_x_inst_n498,
         round_inst_S_4__sbox_inst_com_x_inst_n497,
         round_inst_S_4__sbox_inst_com_x_inst_n496,
         round_inst_S_4__sbox_inst_com_x_inst_n495,
         round_inst_S_4__sbox_inst_com_x_inst_n494,
         round_inst_S_4__sbox_inst_com_x_inst_n493,
         round_inst_S_4__sbox_inst_com_x_inst_n492,
         round_inst_S_4__sbox_inst_com_x_inst_n491,
         round_inst_S_4__sbox_inst_com_x_inst_n490,
         round_inst_S_4__sbox_inst_com_x_inst_n489,
         round_inst_S_4__sbox_inst_com_x_inst_n488,
         round_inst_S_4__sbox_inst_com_x_inst_n487,
         round_inst_S_4__sbox_inst_com_x_inst_n486,
         round_inst_S_4__sbox_inst_com_x_inst_n485,
         round_inst_S_4__sbox_inst_com_x_inst_n484,
         round_inst_S_4__sbox_inst_com_x_inst_n483,
         round_inst_S_4__sbox_inst_com_x_inst_n482,
         round_inst_S_4__sbox_inst_com_x_inst_n481,
         round_inst_S_4__sbox_inst_com_x_inst_n480,
         round_inst_S_4__sbox_inst_com_x_inst_n479,
         round_inst_S_4__sbox_inst_com_x_inst_n478,
         round_inst_S_4__sbox_inst_com_x_inst_n477,
         round_inst_S_4__sbox_inst_com_x_inst_n476,
         round_inst_S_4__sbox_inst_com_x_inst_n475,
         round_inst_S_4__sbox_inst_com_x_inst_n474,
         round_inst_S_4__sbox_inst_com_x_inst_n473,
         round_inst_S_4__sbox_inst_com_x_inst_n472,
         round_inst_S_4__sbox_inst_com_x_inst_n471,
         round_inst_S_4__sbox_inst_com_x_inst_n470,
         round_inst_S_4__sbox_inst_com_x_inst_n469,
         round_inst_S_4__sbox_inst_com_x_inst_n468,
         round_inst_S_4__sbox_inst_com_x_inst_n467,
         round_inst_S_4__sbox_inst_com_x_inst_n466,
         round_inst_S_4__sbox_inst_com_x_inst_n465,
         round_inst_S_4__sbox_inst_com_x_inst_n464,
         round_inst_S_4__sbox_inst_com_x_inst_n463,
         round_inst_S_4__sbox_inst_com_x_inst_n462,
         round_inst_S_4__sbox_inst_com_x_inst_n461,
         round_inst_S_4__sbox_inst_com_x_inst_n460,
         round_inst_S_4__sbox_inst_com_x_inst_n459,
         round_inst_S_4__sbox_inst_com_x_inst_n458,
         round_inst_S_4__sbox_inst_com_x_inst_n457,
         round_inst_S_4__sbox_inst_com_x_inst_n456,
         round_inst_S_4__sbox_inst_com_x_inst_n455,
         round_inst_S_4__sbox_inst_com_x_inst_n454,
         round_inst_S_4__sbox_inst_com_x_inst_n453,
         round_inst_S_4__sbox_inst_com_x_inst_n452,
         round_inst_S_4__sbox_inst_com_x_inst_n451,
         round_inst_S_4__sbox_inst_com_x_inst_n450,
         round_inst_S_4__sbox_inst_com_x_inst_n449,
         round_inst_S_4__sbox_inst_com_x_inst_n448,
         round_inst_S_4__sbox_inst_com_x_inst_n447,
         round_inst_S_4__sbox_inst_com_x_inst_n446,
         round_inst_S_4__sbox_inst_com_x_inst_n445,
         round_inst_S_4__sbox_inst_com_x_inst_n444,
         round_inst_S_4__sbox_inst_com_x_inst_n443,
         round_inst_S_4__sbox_inst_com_x_inst_n442,
         round_inst_S_4__sbox_inst_com_x_inst_n441,
         round_inst_S_4__sbox_inst_com_x_inst_n440,
         round_inst_S_4__sbox_inst_com_x_inst_n439,
         round_inst_S_4__sbox_inst_com_x_inst_n438,
         round_inst_S_4__sbox_inst_com_x_inst_n437,
         round_inst_S_4__sbox_inst_com_x_inst_n436,
         round_inst_S_4__sbox_inst_com_x_inst_n435,
         round_inst_S_4__sbox_inst_com_x_inst_n434,
         round_inst_S_4__sbox_inst_com_x_inst_n433,
         round_inst_S_4__sbox_inst_com_x_inst_n432,
         round_inst_S_4__sbox_inst_com_x_inst_n431,
         round_inst_S_4__sbox_inst_com_x_inst_n430,
         round_inst_S_4__sbox_inst_com_x_inst_n429,
         round_inst_S_4__sbox_inst_com_x_inst_n428,
         round_inst_S_4__sbox_inst_com_x_inst_n427,
         round_inst_S_4__sbox_inst_com_x_inst_n426,
         round_inst_S_4__sbox_inst_com_x_inst_n425,
         round_inst_S_4__sbox_inst_com_x_inst_n424,
         round_inst_S_4__sbox_inst_com_x_inst_n423,
         round_inst_S_4__sbox_inst_com_x_inst_n422,
         round_inst_S_4__sbox_inst_com_x_inst_n421,
         round_inst_S_4__sbox_inst_com_x_inst_n420,
         round_inst_S_4__sbox_inst_com_x_inst_n419,
         round_inst_S_4__sbox_inst_com_x_inst_n418,
         round_inst_S_4__sbox_inst_com_x_inst_n417,
         round_inst_S_4__sbox_inst_com_x_inst_n416,
         round_inst_S_4__sbox_inst_com_x_inst_n415,
         round_inst_S_4__sbox_inst_com_x_inst_n414,
         round_inst_S_4__sbox_inst_com_x_inst_n413,
         round_inst_S_4__sbox_inst_com_x_inst_n412,
         round_inst_S_4__sbox_inst_com_x_inst_n411,
         round_inst_S_4__sbox_inst_com_x_inst_n410,
         round_inst_S_4__sbox_inst_com_x_inst_n409,
         round_inst_S_4__sbox_inst_com_x_inst_n408,
         round_inst_S_4__sbox_inst_com_x_inst_n407,
         round_inst_S_4__sbox_inst_com_x_inst_n406,
         round_inst_S_4__sbox_inst_com_x_inst_n405,
         round_inst_S_4__sbox_inst_com_x_inst_n404,
         round_inst_S_4__sbox_inst_com_x_inst_n403,
         round_inst_S_4__sbox_inst_com_x_inst_n402,
         round_inst_S_4__sbox_inst_com_x_inst_n401,
         round_inst_S_4__sbox_inst_com_x_inst_n400,
         round_inst_S_4__sbox_inst_com_x_inst_n399,
         round_inst_S_4__sbox_inst_com_x_inst_n398,
         round_inst_S_4__sbox_inst_com_x_inst_n397,
         round_inst_S_4__sbox_inst_com_x_inst_n396,
         round_inst_S_4__sbox_inst_com_x_inst_n395,
         round_inst_S_4__sbox_inst_com_x_inst_n394,
         round_inst_S_4__sbox_inst_com_x_inst_n393,
         round_inst_S_4__sbox_inst_com_x_inst_n392,
         round_inst_S_4__sbox_inst_com_x_inst_n391,
         round_inst_S_4__sbox_inst_com_x_inst_n390,
         round_inst_S_4__sbox_inst_com_x_inst_n389,
         round_inst_S_4__sbox_inst_com_x_inst_n388,
         round_inst_S_4__sbox_inst_com_x_inst_n387,
         round_inst_S_4__sbox_inst_com_x_inst_n386,
         round_inst_S_4__sbox_inst_com_x_inst_n385,
         round_inst_S_4__sbox_inst_com_x_inst_n384,
         round_inst_S_4__sbox_inst_com_x_inst_n383,
         round_inst_S_4__sbox_inst_com_x_inst_n382,
         round_inst_S_4__sbox_inst_com_x_inst_n381,
         round_inst_S_4__sbox_inst_com_y_inst_n518,
         round_inst_S_4__sbox_inst_com_y_inst_n517,
         round_inst_S_4__sbox_inst_com_y_inst_n516,
         round_inst_S_4__sbox_inst_com_y_inst_n515,
         round_inst_S_4__sbox_inst_com_y_inst_n514,
         round_inst_S_4__sbox_inst_com_y_inst_n513,
         round_inst_S_4__sbox_inst_com_y_inst_n512,
         round_inst_S_4__sbox_inst_com_y_inst_n511,
         round_inst_S_4__sbox_inst_com_y_inst_n510,
         round_inst_S_4__sbox_inst_com_y_inst_n509,
         round_inst_S_4__sbox_inst_com_y_inst_n508,
         round_inst_S_4__sbox_inst_com_y_inst_n507,
         round_inst_S_4__sbox_inst_com_y_inst_n506,
         round_inst_S_4__sbox_inst_com_y_inst_n505,
         round_inst_S_4__sbox_inst_com_y_inst_n504,
         round_inst_S_4__sbox_inst_com_y_inst_n503,
         round_inst_S_4__sbox_inst_com_y_inst_n502,
         round_inst_S_4__sbox_inst_com_y_inst_n501,
         round_inst_S_4__sbox_inst_com_y_inst_n500,
         round_inst_S_4__sbox_inst_com_y_inst_n499,
         round_inst_S_4__sbox_inst_com_y_inst_n498,
         round_inst_S_4__sbox_inst_com_y_inst_n497,
         round_inst_S_4__sbox_inst_com_y_inst_n496,
         round_inst_S_4__sbox_inst_com_y_inst_n495,
         round_inst_S_4__sbox_inst_com_y_inst_n494,
         round_inst_S_4__sbox_inst_com_y_inst_n493,
         round_inst_S_4__sbox_inst_com_y_inst_n492,
         round_inst_S_4__sbox_inst_com_y_inst_n491,
         round_inst_S_4__sbox_inst_com_y_inst_n490,
         round_inst_S_4__sbox_inst_com_y_inst_n489,
         round_inst_S_4__sbox_inst_com_y_inst_n488,
         round_inst_S_4__sbox_inst_com_y_inst_n487,
         round_inst_S_4__sbox_inst_com_y_inst_n486,
         round_inst_S_4__sbox_inst_com_y_inst_n485,
         round_inst_S_4__sbox_inst_com_y_inst_n484,
         round_inst_S_4__sbox_inst_com_y_inst_n483,
         round_inst_S_4__sbox_inst_com_y_inst_n482,
         round_inst_S_4__sbox_inst_com_y_inst_n481,
         round_inst_S_4__sbox_inst_com_y_inst_n480,
         round_inst_S_4__sbox_inst_com_y_inst_n479,
         round_inst_S_4__sbox_inst_com_y_inst_n478,
         round_inst_S_4__sbox_inst_com_y_inst_n477,
         round_inst_S_4__sbox_inst_com_y_inst_n476,
         round_inst_S_4__sbox_inst_com_y_inst_n475,
         round_inst_S_4__sbox_inst_com_y_inst_n474,
         round_inst_S_4__sbox_inst_com_y_inst_n473,
         round_inst_S_4__sbox_inst_com_y_inst_n472,
         round_inst_S_4__sbox_inst_com_y_inst_n471,
         round_inst_S_4__sbox_inst_com_y_inst_n470,
         round_inst_S_4__sbox_inst_com_y_inst_n469,
         round_inst_S_4__sbox_inst_com_y_inst_n468,
         round_inst_S_4__sbox_inst_com_y_inst_n467,
         round_inst_S_4__sbox_inst_com_y_inst_n466,
         round_inst_S_4__sbox_inst_com_y_inst_n465,
         round_inst_S_4__sbox_inst_com_y_inst_n464,
         round_inst_S_4__sbox_inst_com_y_inst_n463,
         round_inst_S_4__sbox_inst_com_y_inst_n462,
         round_inst_S_4__sbox_inst_com_y_inst_n461,
         round_inst_S_4__sbox_inst_com_y_inst_n460,
         round_inst_S_4__sbox_inst_com_y_inst_n459,
         round_inst_S_4__sbox_inst_com_y_inst_n458,
         round_inst_S_4__sbox_inst_com_y_inst_n457,
         round_inst_S_4__sbox_inst_com_y_inst_n456,
         round_inst_S_4__sbox_inst_com_y_inst_n455,
         round_inst_S_4__sbox_inst_com_y_inst_n454,
         round_inst_S_4__sbox_inst_com_y_inst_n453,
         round_inst_S_4__sbox_inst_com_y_inst_n452,
         round_inst_S_4__sbox_inst_com_y_inst_n451,
         round_inst_S_4__sbox_inst_com_y_inst_n450,
         round_inst_S_4__sbox_inst_com_y_inst_n449,
         round_inst_S_4__sbox_inst_com_y_inst_n448,
         round_inst_S_4__sbox_inst_com_y_inst_n447,
         round_inst_S_4__sbox_inst_com_y_inst_n446,
         round_inst_S_4__sbox_inst_com_y_inst_n445,
         round_inst_S_4__sbox_inst_com_y_inst_n444,
         round_inst_S_4__sbox_inst_com_y_inst_n443,
         round_inst_S_4__sbox_inst_com_y_inst_n442,
         round_inst_S_4__sbox_inst_com_y_inst_n441,
         round_inst_S_4__sbox_inst_com_y_inst_n440,
         round_inst_S_4__sbox_inst_com_y_inst_n439,
         round_inst_S_4__sbox_inst_com_y_inst_n438,
         round_inst_S_4__sbox_inst_com_y_inst_n437,
         round_inst_S_4__sbox_inst_com_y_inst_n436,
         round_inst_S_4__sbox_inst_com_y_inst_n435,
         round_inst_S_4__sbox_inst_com_y_inst_n434,
         round_inst_S_4__sbox_inst_com_y_inst_n433,
         round_inst_S_4__sbox_inst_com_y_inst_n432,
         round_inst_S_4__sbox_inst_com_y_inst_n431,
         round_inst_S_4__sbox_inst_com_y_inst_n430,
         round_inst_S_4__sbox_inst_com_y_inst_n429,
         round_inst_S_4__sbox_inst_com_y_inst_n428,
         round_inst_S_4__sbox_inst_com_y_inst_n427,
         round_inst_S_4__sbox_inst_com_y_inst_n426,
         round_inst_S_4__sbox_inst_com_y_inst_n425,
         round_inst_S_4__sbox_inst_com_y_inst_n424,
         round_inst_S_4__sbox_inst_com_y_inst_n423,
         round_inst_S_4__sbox_inst_com_y_inst_n422,
         round_inst_S_4__sbox_inst_com_y_inst_n421,
         round_inst_S_4__sbox_inst_com_y_inst_n420,
         round_inst_S_4__sbox_inst_com_y_inst_n419,
         round_inst_S_4__sbox_inst_com_y_inst_n418,
         round_inst_S_4__sbox_inst_com_y_inst_n417,
         round_inst_S_4__sbox_inst_com_y_inst_n416,
         round_inst_S_4__sbox_inst_com_y_inst_n415,
         round_inst_S_4__sbox_inst_com_y_inst_n414,
         round_inst_S_4__sbox_inst_com_y_inst_n413,
         round_inst_S_4__sbox_inst_com_y_inst_n412,
         round_inst_S_4__sbox_inst_com_y_inst_n411,
         round_inst_S_4__sbox_inst_com_y_inst_n410,
         round_inst_S_4__sbox_inst_com_y_inst_n409,
         round_inst_S_4__sbox_inst_com_y_inst_n408,
         round_inst_S_4__sbox_inst_com_y_inst_n407,
         round_inst_S_4__sbox_inst_com_y_inst_n406,
         round_inst_S_4__sbox_inst_com_y_inst_n405,
         round_inst_S_4__sbox_inst_com_y_inst_n404,
         round_inst_S_4__sbox_inst_com_y_inst_n403,
         round_inst_S_4__sbox_inst_com_y_inst_n402,
         round_inst_S_4__sbox_inst_com_y_inst_n401,
         round_inst_S_4__sbox_inst_com_y_inst_n400,
         round_inst_S_4__sbox_inst_com_y_inst_n399,
         round_inst_S_4__sbox_inst_com_y_inst_n398,
         round_inst_S_4__sbox_inst_com_y_inst_n397,
         round_inst_S_4__sbox_inst_com_y_inst_n396,
         round_inst_S_4__sbox_inst_com_y_inst_n395,
         round_inst_S_4__sbox_inst_com_y_inst_n394,
         round_inst_S_4__sbox_inst_com_y_inst_n393,
         round_inst_S_4__sbox_inst_com_y_inst_n392,
         round_inst_S_4__sbox_inst_com_y_inst_n391,
         round_inst_S_4__sbox_inst_com_y_inst_n390,
         round_inst_S_4__sbox_inst_com_y_inst_n389,
         round_inst_S_4__sbox_inst_com_y_inst_n388,
         round_inst_S_4__sbox_inst_com_y_inst_n387,
         round_inst_S_4__sbox_inst_com_y_inst_n386,
         round_inst_S_4__sbox_inst_com_z_inst_n516,
         round_inst_S_4__sbox_inst_com_z_inst_n515,
         round_inst_S_4__sbox_inst_com_z_inst_n514,
         round_inst_S_4__sbox_inst_com_z_inst_n513,
         round_inst_S_4__sbox_inst_com_z_inst_n512,
         round_inst_S_4__sbox_inst_com_z_inst_n511,
         round_inst_S_4__sbox_inst_com_z_inst_n510,
         round_inst_S_4__sbox_inst_com_z_inst_n509,
         round_inst_S_4__sbox_inst_com_z_inst_n508,
         round_inst_S_4__sbox_inst_com_z_inst_n507,
         round_inst_S_4__sbox_inst_com_z_inst_n506,
         round_inst_S_4__sbox_inst_com_z_inst_n505,
         round_inst_S_4__sbox_inst_com_z_inst_n504,
         round_inst_S_4__sbox_inst_com_z_inst_n503,
         round_inst_S_4__sbox_inst_com_z_inst_n502,
         round_inst_S_4__sbox_inst_com_z_inst_n501,
         round_inst_S_4__sbox_inst_com_z_inst_n500,
         round_inst_S_4__sbox_inst_com_z_inst_n499,
         round_inst_S_4__sbox_inst_com_z_inst_n498,
         round_inst_S_4__sbox_inst_com_z_inst_n497,
         round_inst_S_4__sbox_inst_com_z_inst_n496,
         round_inst_S_4__sbox_inst_com_z_inst_n495,
         round_inst_S_4__sbox_inst_com_z_inst_n494,
         round_inst_S_4__sbox_inst_com_z_inst_n493,
         round_inst_S_4__sbox_inst_com_z_inst_n492,
         round_inst_S_4__sbox_inst_com_z_inst_n491,
         round_inst_S_4__sbox_inst_com_z_inst_n490,
         round_inst_S_4__sbox_inst_com_z_inst_n489,
         round_inst_S_4__sbox_inst_com_z_inst_n488,
         round_inst_S_4__sbox_inst_com_z_inst_n487,
         round_inst_S_4__sbox_inst_com_z_inst_n486,
         round_inst_S_4__sbox_inst_com_z_inst_n485,
         round_inst_S_4__sbox_inst_com_z_inst_n484,
         round_inst_S_4__sbox_inst_com_z_inst_n483,
         round_inst_S_4__sbox_inst_com_z_inst_n482,
         round_inst_S_4__sbox_inst_com_z_inst_n481,
         round_inst_S_4__sbox_inst_com_z_inst_n480,
         round_inst_S_4__sbox_inst_com_z_inst_n479,
         round_inst_S_4__sbox_inst_com_z_inst_n478,
         round_inst_S_4__sbox_inst_com_z_inst_n477,
         round_inst_S_4__sbox_inst_com_z_inst_n476,
         round_inst_S_4__sbox_inst_com_z_inst_n475,
         round_inst_S_4__sbox_inst_com_z_inst_n474,
         round_inst_S_4__sbox_inst_com_z_inst_n473,
         round_inst_S_4__sbox_inst_com_z_inst_n472,
         round_inst_S_4__sbox_inst_com_z_inst_n471,
         round_inst_S_4__sbox_inst_com_z_inst_n470,
         round_inst_S_4__sbox_inst_com_z_inst_n469,
         round_inst_S_4__sbox_inst_com_z_inst_n468,
         round_inst_S_4__sbox_inst_com_z_inst_n467,
         round_inst_S_4__sbox_inst_com_z_inst_n466,
         round_inst_S_4__sbox_inst_com_z_inst_n465,
         round_inst_S_4__sbox_inst_com_z_inst_n464,
         round_inst_S_4__sbox_inst_com_z_inst_n463,
         round_inst_S_4__sbox_inst_com_z_inst_n462,
         round_inst_S_4__sbox_inst_com_z_inst_n461,
         round_inst_S_4__sbox_inst_com_z_inst_n460,
         round_inst_S_4__sbox_inst_com_z_inst_n459,
         round_inst_S_4__sbox_inst_com_z_inst_n458,
         round_inst_S_4__sbox_inst_com_z_inst_n457,
         round_inst_S_4__sbox_inst_com_z_inst_n456,
         round_inst_S_4__sbox_inst_com_z_inst_n455,
         round_inst_S_4__sbox_inst_com_z_inst_n454,
         round_inst_S_4__sbox_inst_com_z_inst_n453,
         round_inst_S_4__sbox_inst_com_z_inst_n452,
         round_inst_S_4__sbox_inst_com_z_inst_n451,
         round_inst_S_4__sbox_inst_com_z_inst_n450,
         round_inst_S_4__sbox_inst_com_z_inst_n449,
         round_inst_S_4__sbox_inst_com_z_inst_n448,
         round_inst_S_4__sbox_inst_com_z_inst_n447,
         round_inst_S_4__sbox_inst_com_z_inst_n446,
         round_inst_S_4__sbox_inst_com_z_inst_n445,
         round_inst_S_4__sbox_inst_com_z_inst_n444,
         round_inst_S_4__sbox_inst_com_z_inst_n443,
         round_inst_S_4__sbox_inst_com_z_inst_n442,
         round_inst_S_4__sbox_inst_com_z_inst_n441,
         round_inst_S_4__sbox_inst_com_z_inst_n440,
         round_inst_S_4__sbox_inst_com_z_inst_n439,
         round_inst_S_4__sbox_inst_com_z_inst_n438,
         round_inst_S_4__sbox_inst_com_z_inst_n437,
         round_inst_S_4__sbox_inst_com_z_inst_n436,
         round_inst_S_4__sbox_inst_com_z_inst_n435,
         round_inst_S_4__sbox_inst_com_z_inst_n434,
         round_inst_S_4__sbox_inst_com_z_inst_n433,
         round_inst_S_4__sbox_inst_com_z_inst_n432,
         round_inst_S_4__sbox_inst_com_z_inst_n431,
         round_inst_S_4__sbox_inst_com_z_inst_n430,
         round_inst_S_4__sbox_inst_com_z_inst_n429,
         round_inst_S_4__sbox_inst_com_z_inst_n428,
         round_inst_S_4__sbox_inst_com_z_inst_n427,
         round_inst_S_4__sbox_inst_com_z_inst_n426,
         round_inst_S_4__sbox_inst_com_z_inst_n425,
         round_inst_S_4__sbox_inst_com_z_inst_n424,
         round_inst_S_4__sbox_inst_com_z_inst_n423,
         round_inst_S_4__sbox_inst_com_z_inst_n422,
         round_inst_S_4__sbox_inst_com_z_inst_n421,
         round_inst_S_4__sbox_inst_com_z_inst_n420,
         round_inst_S_4__sbox_inst_com_z_inst_n419,
         round_inst_S_4__sbox_inst_com_z_inst_n418,
         round_inst_S_4__sbox_inst_com_z_inst_n417,
         round_inst_S_4__sbox_inst_com_z_inst_n416,
         round_inst_S_4__sbox_inst_com_z_inst_n415,
         round_inst_S_4__sbox_inst_com_z_inst_n414,
         round_inst_S_4__sbox_inst_com_z_inst_n413,
         round_inst_S_4__sbox_inst_com_z_inst_n412,
         round_inst_S_4__sbox_inst_com_z_inst_n411,
         round_inst_S_4__sbox_inst_com_z_inst_n410,
         round_inst_S_4__sbox_inst_com_z_inst_n409,
         round_inst_S_4__sbox_inst_com_z_inst_n408,
         round_inst_S_4__sbox_inst_com_z_inst_n407,
         round_inst_S_4__sbox_inst_com_z_inst_n406,
         round_inst_S_4__sbox_inst_com_z_inst_n405,
         round_inst_S_4__sbox_inst_com_z_inst_n404,
         round_inst_S_4__sbox_inst_com_z_inst_n403,
         round_inst_S_4__sbox_inst_com_z_inst_n402,
         round_inst_S_4__sbox_inst_com_z_inst_n401,
         round_inst_S_4__sbox_inst_com_z_inst_n400,
         round_inst_S_4__sbox_inst_com_z_inst_n399,
         round_inst_S_4__sbox_inst_com_z_inst_n398,
         round_inst_S_4__sbox_inst_com_z_inst_n397,
         round_inst_S_4__sbox_inst_com_z_inst_n396,
         round_inst_S_4__sbox_inst_com_z_inst_n395,
         round_inst_S_4__sbox_inst_com_z_inst_n394,
         round_inst_S_4__sbox_inst_com_z_inst_n393,
         round_inst_S_4__sbox_inst_com_z_inst_n392,
         round_inst_S_4__sbox_inst_com_z_inst_n391,
         round_inst_S_4__sbox_inst_com_z_inst_n390,
         round_inst_S_5__sbox_inst_n6, round_inst_S_5__sbox_inst_n5,
         round_inst_S_5__sbox_inst_n4, round_inst_S_5__sbox_inst_n3,
         round_inst_S_5__sbox_inst_n2, round_inst_S_5__sbox_inst_n1,
         round_inst_S_5__sbox_inst_com_w_inst_n532,
         round_inst_S_5__sbox_inst_com_w_inst_n531,
         round_inst_S_5__sbox_inst_com_w_inst_n530,
         round_inst_S_5__sbox_inst_com_w_inst_n529,
         round_inst_S_5__sbox_inst_com_w_inst_n528,
         round_inst_S_5__sbox_inst_com_w_inst_n527,
         round_inst_S_5__sbox_inst_com_w_inst_n526,
         round_inst_S_5__sbox_inst_com_w_inst_n525,
         round_inst_S_5__sbox_inst_com_w_inst_n524,
         round_inst_S_5__sbox_inst_com_w_inst_n523,
         round_inst_S_5__sbox_inst_com_w_inst_n522,
         round_inst_S_5__sbox_inst_com_w_inst_n521,
         round_inst_S_5__sbox_inst_com_w_inst_n520,
         round_inst_S_5__sbox_inst_com_w_inst_n519,
         round_inst_S_5__sbox_inst_com_w_inst_n518,
         round_inst_S_5__sbox_inst_com_w_inst_n517,
         round_inst_S_5__sbox_inst_com_w_inst_n516,
         round_inst_S_5__sbox_inst_com_w_inst_n515,
         round_inst_S_5__sbox_inst_com_w_inst_n514,
         round_inst_S_5__sbox_inst_com_w_inst_n513,
         round_inst_S_5__sbox_inst_com_w_inst_n512,
         round_inst_S_5__sbox_inst_com_w_inst_n511,
         round_inst_S_5__sbox_inst_com_w_inst_n510,
         round_inst_S_5__sbox_inst_com_w_inst_n509,
         round_inst_S_5__sbox_inst_com_w_inst_n508,
         round_inst_S_5__sbox_inst_com_w_inst_n507,
         round_inst_S_5__sbox_inst_com_w_inst_n506,
         round_inst_S_5__sbox_inst_com_w_inst_n505,
         round_inst_S_5__sbox_inst_com_w_inst_n504,
         round_inst_S_5__sbox_inst_com_w_inst_n503,
         round_inst_S_5__sbox_inst_com_w_inst_n502,
         round_inst_S_5__sbox_inst_com_w_inst_n501,
         round_inst_S_5__sbox_inst_com_w_inst_n500,
         round_inst_S_5__sbox_inst_com_w_inst_n499,
         round_inst_S_5__sbox_inst_com_w_inst_n498,
         round_inst_S_5__sbox_inst_com_w_inst_n497,
         round_inst_S_5__sbox_inst_com_w_inst_n496,
         round_inst_S_5__sbox_inst_com_w_inst_n495,
         round_inst_S_5__sbox_inst_com_w_inst_n494,
         round_inst_S_5__sbox_inst_com_w_inst_n493,
         round_inst_S_5__sbox_inst_com_w_inst_n492,
         round_inst_S_5__sbox_inst_com_w_inst_n491,
         round_inst_S_5__sbox_inst_com_w_inst_n490,
         round_inst_S_5__sbox_inst_com_w_inst_n489,
         round_inst_S_5__sbox_inst_com_w_inst_n488,
         round_inst_S_5__sbox_inst_com_w_inst_n487,
         round_inst_S_5__sbox_inst_com_w_inst_n486,
         round_inst_S_5__sbox_inst_com_w_inst_n485,
         round_inst_S_5__sbox_inst_com_w_inst_n484,
         round_inst_S_5__sbox_inst_com_w_inst_n483,
         round_inst_S_5__sbox_inst_com_w_inst_n482,
         round_inst_S_5__sbox_inst_com_w_inst_n481,
         round_inst_S_5__sbox_inst_com_w_inst_n480,
         round_inst_S_5__sbox_inst_com_w_inst_n479,
         round_inst_S_5__sbox_inst_com_w_inst_n478,
         round_inst_S_5__sbox_inst_com_w_inst_n477,
         round_inst_S_5__sbox_inst_com_w_inst_n476,
         round_inst_S_5__sbox_inst_com_w_inst_n475,
         round_inst_S_5__sbox_inst_com_w_inst_n474,
         round_inst_S_5__sbox_inst_com_w_inst_n473,
         round_inst_S_5__sbox_inst_com_w_inst_n472,
         round_inst_S_5__sbox_inst_com_w_inst_n471,
         round_inst_S_5__sbox_inst_com_w_inst_n470,
         round_inst_S_5__sbox_inst_com_w_inst_n469,
         round_inst_S_5__sbox_inst_com_w_inst_n468,
         round_inst_S_5__sbox_inst_com_w_inst_n467,
         round_inst_S_5__sbox_inst_com_w_inst_n466,
         round_inst_S_5__sbox_inst_com_w_inst_n465,
         round_inst_S_5__sbox_inst_com_w_inst_n464,
         round_inst_S_5__sbox_inst_com_w_inst_n463,
         round_inst_S_5__sbox_inst_com_w_inst_n462,
         round_inst_S_5__sbox_inst_com_w_inst_n461,
         round_inst_S_5__sbox_inst_com_w_inst_n460,
         round_inst_S_5__sbox_inst_com_w_inst_n459,
         round_inst_S_5__sbox_inst_com_w_inst_n458,
         round_inst_S_5__sbox_inst_com_w_inst_n457,
         round_inst_S_5__sbox_inst_com_w_inst_n456,
         round_inst_S_5__sbox_inst_com_w_inst_n455,
         round_inst_S_5__sbox_inst_com_w_inst_n454,
         round_inst_S_5__sbox_inst_com_w_inst_n453,
         round_inst_S_5__sbox_inst_com_w_inst_n452,
         round_inst_S_5__sbox_inst_com_w_inst_n451,
         round_inst_S_5__sbox_inst_com_w_inst_n450,
         round_inst_S_5__sbox_inst_com_w_inst_n449,
         round_inst_S_5__sbox_inst_com_w_inst_n448,
         round_inst_S_5__sbox_inst_com_w_inst_n447,
         round_inst_S_5__sbox_inst_com_w_inst_n446,
         round_inst_S_5__sbox_inst_com_w_inst_n445,
         round_inst_S_5__sbox_inst_com_w_inst_n444,
         round_inst_S_5__sbox_inst_com_w_inst_n443,
         round_inst_S_5__sbox_inst_com_w_inst_n442,
         round_inst_S_5__sbox_inst_com_w_inst_n441,
         round_inst_S_5__sbox_inst_com_w_inst_n440,
         round_inst_S_5__sbox_inst_com_w_inst_n439,
         round_inst_S_5__sbox_inst_com_w_inst_n438,
         round_inst_S_5__sbox_inst_com_w_inst_n437,
         round_inst_S_5__sbox_inst_com_w_inst_n436,
         round_inst_S_5__sbox_inst_com_w_inst_n435,
         round_inst_S_5__sbox_inst_com_w_inst_n434,
         round_inst_S_5__sbox_inst_com_w_inst_n433,
         round_inst_S_5__sbox_inst_com_w_inst_n432,
         round_inst_S_5__sbox_inst_com_w_inst_n431,
         round_inst_S_5__sbox_inst_com_w_inst_n430,
         round_inst_S_5__sbox_inst_com_w_inst_n429,
         round_inst_S_5__sbox_inst_com_w_inst_n428,
         round_inst_S_5__sbox_inst_com_w_inst_n427,
         round_inst_S_5__sbox_inst_com_w_inst_n426,
         round_inst_S_5__sbox_inst_com_w_inst_n425,
         round_inst_S_5__sbox_inst_com_w_inst_n424,
         round_inst_S_5__sbox_inst_com_w_inst_n423,
         round_inst_S_5__sbox_inst_com_w_inst_n422,
         round_inst_S_5__sbox_inst_com_w_inst_n421,
         round_inst_S_5__sbox_inst_com_w_inst_n420,
         round_inst_S_5__sbox_inst_com_w_inst_n419,
         round_inst_S_5__sbox_inst_com_w_inst_n418,
         round_inst_S_5__sbox_inst_com_w_inst_n417,
         round_inst_S_5__sbox_inst_com_w_inst_n416,
         round_inst_S_5__sbox_inst_com_w_inst_n415,
         round_inst_S_5__sbox_inst_com_w_inst_n414,
         round_inst_S_5__sbox_inst_com_w_inst_n413,
         round_inst_S_5__sbox_inst_com_w_inst_n412,
         round_inst_S_5__sbox_inst_com_w_inst_n411,
         round_inst_S_5__sbox_inst_com_w_inst_n410,
         round_inst_S_5__sbox_inst_com_w_inst_n409,
         round_inst_S_5__sbox_inst_com_w_inst_n408,
         round_inst_S_5__sbox_inst_com_w_inst_n407,
         round_inst_S_5__sbox_inst_com_w_inst_n406,
         round_inst_S_5__sbox_inst_com_w_inst_n405,
         round_inst_S_5__sbox_inst_com_w_inst_n404,
         round_inst_S_5__sbox_inst_com_w_inst_n403,
         round_inst_S_5__sbox_inst_com_w_inst_n402,
         round_inst_S_5__sbox_inst_com_w_inst_n401,
         round_inst_S_5__sbox_inst_com_w_inst_n400,
         round_inst_S_5__sbox_inst_com_w_inst_n399,
         round_inst_S_5__sbox_inst_com_w_inst_n398,
         round_inst_S_5__sbox_inst_com_w_inst_n397,
         round_inst_S_5__sbox_inst_com_w_inst_n396,
         round_inst_S_5__sbox_inst_com_x_inst_n511,
         round_inst_S_5__sbox_inst_com_x_inst_n510,
         round_inst_S_5__sbox_inst_com_x_inst_n509,
         round_inst_S_5__sbox_inst_com_x_inst_n508,
         round_inst_S_5__sbox_inst_com_x_inst_n507,
         round_inst_S_5__sbox_inst_com_x_inst_n506,
         round_inst_S_5__sbox_inst_com_x_inst_n505,
         round_inst_S_5__sbox_inst_com_x_inst_n504,
         round_inst_S_5__sbox_inst_com_x_inst_n503,
         round_inst_S_5__sbox_inst_com_x_inst_n502,
         round_inst_S_5__sbox_inst_com_x_inst_n501,
         round_inst_S_5__sbox_inst_com_x_inst_n500,
         round_inst_S_5__sbox_inst_com_x_inst_n499,
         round_inst_S_5__sbox_inst_com_x_inst_n498,
         round_inst_S_5__sbox_inst_com_x_inst_n497,
         round_inst_S_5__sbox_inst_com_x_inst_n496,
         round_inst_S_5__sbox_inst_com_x_inst_n495,
         round_inst_S_5__sbox_inst_com_x_inst_n494,
         round_inst_S_5__sbox_inst_com_x_inst_n493,
         round_inst_S_5__sbox_inst_com_x_inst_n492,
         round_inst_S_5__sbox_inst_com_x_inst_n491,
         round_inst_S_5__sbox_inst_com_x_inst_n490,
         round_inst_S_5__sbox_inst_com_x_inst_n489,
         round_inst_S_5__sbox_inst_com_x_inst_n488,
         round_inst_S_5__sbox_inst_com_x_inst_n487,
         round_inst_S_5__sbox_inst_com_x_inst_n486,
         round_inst_S_5__sbox_inst_com_x_inst_n485,
         round_inst_S_5__sbox_inst_com_x_inst_n484,
         round_inst_S_5__sbox_inst_com_x_inst_n483,
         round_inst_S_5__sbox_inst_com_x_inst_n482,
         round_inst_S_5__sbox_inst_com_x_inst_n481,
         round_inst_S_5__sbox_inst_com_x_inst_n480,
         round_inst_S_5__sbox_inst_com_x_inst_n479,
         round_inst_S_5__sbox_inst_com_x_inst_n478,
         round_inst_S_5__sbox_inst_com_x_inst_n477,
         round_inst_S_5__sbox_inst_com_x_inst_n476,
         round_inst_S_5__sbox_inst_com_x_inst_n475,
         round_inst_S_5__sbox_inst_com_x_inst_n474,
         round_inst_S_5__sbox_inst_com_x_inst_n473,
         round_inst_S_5__sbox_inst_com_x_inst_n472,
         round_inst_S_5__sbox_inst_com_x_inst_n471,
         round_inst_S_5__sbox_inst_com_x_inst_n470,
         round_inst_S_5__sbox_inst_com_x_inst_n469,
         round_inst_S_5__sbox_inst_com_x_inst_n468,
         round_inst_S_5__sbox_inst_com_x_inst_n467,
         round_inst_S_5__sbox_inst_com_x_inst_n466,
         round_inst_S_5__sbox_inst_com_x_inst_n465,
         round_inst_S_5__sbox_inst_com_x_inst_n464,
         round_inst_S_5__sbox_inst_com_x_inst_n463,
         round_inst_S_5__sbox_inst_com_x_inst_n462,
         round_inst_S_5__sbox_inst_com_x_inst_n461,
         round_inst_S_5__sbox_inst_com_x_inst_n460,
         round_inst_S_5__sbox_inst_com_x_inst_n459,
         round_inst_S_5__sbox_inst_com_x_inst_n458,
         round_inst_S_5__sbox_inst_com_x_inst_n457,
         round_inst_S_5__sbox_inst_com_x_inst_n456,
         round_inst_S_5__sbox_inst_com_x_inst_n455,
         round_inst_S_5__sbox_inst_com_x_inst_n454,
         round_inst_S_5__sbox_inst_com_x_inst_n453,
         round_inst_S_5__sbox_inst_com_x_inst_n452,
         round_inst_S_5__sbox_inst_com_x_inst_n451,
         round_inst_S_5__sbox_inst_com_x_inst_n450,
         round_inst_S_5__sbox_inst_com_x_inst_n449,
         round_inst_S_5__sbox_inst_com_x_inst_n448,
         round_inst_S_5__sbox_inst_com_x_inst_n447,
         round_inst_S_5__sbox_inst_com_x_inst_n446,
         round_inst_S_5__sbox_inst_com_x_inst_n445,
         round_inst_S_5__sbox_inst_com_x_inst_n444,
         round_inst_S_5__sbox_inst_com_x_inst_n443,
         round_inst_S_5__sbox_inst_com_x_inst_n442,
         round_inst_S_5__sbox_inst_com_x_inst_n441,
         round_inst_S_5__sbox_inst_com_x_inst_n440,
         round_inst_S_5__sbox_inst_com_x_inst_n439,
         round_inst_S_5__sbox_inst_com_x_inst_n438,
         round_inst_S_5__sbox_inst_com_x_inst_n437,
         round_inst_S_5__sbox_inst_com_x_inst_n436,
         round_inst_S_5__sbox_inst_com_x_inst_n435,
         round_inst_S_5__sbox_inst_com_x_inst_n434,
         round_inst_S_5__sbox_inst_com_x_inst_n433,
         round_inst_S_5__sbox_inst_com_x_inst_n432,
         round_inst_S_5__sbox_inst_com_x_inst_n431,
         round_inst_S_5__sbox_inst_com_x_inst_n430,
         round_inst_S_5__sbox_inst_com_x_inst_n429,
         round_inst_S_5__sbox_inst_com_x_inst_n428,
         round_inst_S_5__sbox_inst_com_x_inst_n427,
         round_inst_S_5__sbox_inst_com_x_inst_n426,
         round_inst_S_5__sbox_inst_com_x_inst_n425,
         round_inst_S_5__sbox_inst_com_x_inst_n424,
         round_inst_S_5__sbox_inst_com_x_inst_n423,
         round_inst_S_5__sbox_inst_com_x_inst_n422,
         round_inst_S_5__sbox_inst_com_x_inst_n421,
         round_inst_S_5__sbox_inst_com_x_inst_n420,
         round_inst_S_5__sbox_inst_com_x_inst_n419,
         round_inst_S_5__sbox_inst_com_x_inst_n418,
         round_inst_S_5__sbox_inst_com_x_inst_n417,
         round_inst_S_5__sbox_inst_com_x_inst_n416,
         round_inst_S_5__sbox_inst_com_x_inst_n415,
         round_inst_S_5__sbox_inst_com_x_inst_n414,
         round_inst_S_5__sbox_inst_com_x_inst_n413,
         round_inst_S_5__sbox_inst_com_x_inst_n412,
         round_inst_S_5__sbox_inst_com_x_inst_n411,
         round_inst_S_5__sbox_inst_com_x_inst_n410,
         round_inst_S_5__sbox_inst_com_x_inst_n409,
         round_inst_S_5__sbox_inst_com_x_inst_n408,
         round_inst_S_5__sbox_inst_com_x_inst_n407,
         round_inst_S_5__sbox_inst_com_x_inst_n406,
         round_inst_S_5__sbox_inst_com_x_inst_n405,
         round_inst_S_5__sbox_inst_com_x_inst_n404,
         round_inst_S_5__sbox_inst_com_x_inst_n403,
         round_inst_S_5__sbox_inst_com_x_inst_n402,
         round_inst_S_5__sbox_inst_com_x_inst_n401,
         round_inst_S_5__sbox_inst_com_x_inst_n400,
         round_inst_S_5__sbox_inst_com_x_inst_n399,
         round_inst_S_5__sbox_inst_com_x_inst_n398,
         round_inst_S_5__sbox_inst_com_x_inst_n397,
         round_inst_S_5__sbox_inst_com_x_inst_n396,
         round_inst_S_5__sbox_inst_com_x_inst_n395,
         round_inst_S_5__sbox_inst_com_x_inst_n394,
         round_inst_S_5__sbox_inst_com_x_inst_n393,
         round_inst_S_5__sbox_inst_com_x_inst_n392,
         round_inst_S_5__sbox_inst_com_x_inst_n391,
         round_inst_S_5__sbox_inst_com_x_inst_n390,
         round_inst_S_5__sbox_inst_com_x_inst_n389,
         round_inst_S_5__sbox_inst_com_x_inst_n388,
         round_inst_S_5__sbox_inst_com_x_inst_n387,
         round_inst_S_5__sbox_inst_com_x_inst_n386,
         round_inst_S_5__sbox_inst_com_x_inst_n385,
         round_inst_S_5__sbox_inst_com_x_inst_n384,
         round_inst_S_5__sbox_inst_com_x_inst_n383,
         round_inst_S_5__sbox_inst_com_x_inst_n382,
         round_inst_S_5__sbox_inst_com_x_inst_n381,
         round_inst_S_5__sbox_inst_com_y_inst_n518,
         round_inst_S_5__sbox_inst_com_y_inst_n517,
         round_inst_S_5__sbox_inst_com_y_inst_n516,
         round_inst_S_5__sbox_inst_com_y_inst_n515,
         round_inst_S_5__sbox_inst_com_y_inst_n514,
         round_inst_S_5__sbox_inst_com_y_inst_n513,
         round_inst_S_5__sbox_inst_com_y_inst_n512,
         round_inst_S_5__sbox_inst_com_y_inst_n511,
         round_inst_S_5__sbox_inst_com_y_inst_n510,
         round_inst_S_5__sbox_inst_com_y_inst_n509,
         round_inst_S_5__sbox_inst_com_y_inst_n508,
         round_inst_S_5__sbox_inst_com_y_inst_n507,
         round_inst_S_5__sbox_inst_com_y_inst_n506,
         round_inst_S_5__sbox_inst_com_y_inst_n505,
         round_inst_S_5__sbox_inst_com_y_inst_n504,
         round_inst_S_5__sbox_inst_com_y_inst_n503,
         round_inst_S_5__sbox_inst_com_y_inst_n502,
         round_inst_S_5__sbox_inst_com_y_inst_n501,
         round_inst_S_5__sbox_inst_com_y_inst_n500,
         round_inst_S_5__sbox_inst_com_y_inst_n499,
         round_inst_S_5__sbox_inst_com_y_inst_n498,
         round_inst_S_5__sbox_inst_com_y_inst_n497,
         round_inst_S_5__sbox_inst_com_y_inst_n496,
         round_inst_S_5__sbox_inst_com_y_inst_n495,
         round_inst_S_5__sbox_inst_com_y_inst_n494,
         round_inst_S_5__sbox_inst_com_y_inst_n493,
         round_inst_S_5__sbox_inst_com_y_inst_n492,
         round_inst_S_5__sbox_inst_com_y_inst_n491,
         round_inst_S_5__sbox_inst_com_y_inst_n490,
         round_inst_S_5__sbox_inst_com_y_inst_n489,
         round_inst_S_5__sbox_inst_com_y_inst_n488,
         round_inst_S_5__sbox_inst_com_y_inst_n487,
         round_inst_S_5__sbox_inst_com_y_inst_n486,
         round_inst_S_5__sbox_inst_com_y_inst_n485,
         round_inst_S_5__sbox_inst_com_y_inst_n484,
         round_inst_S_5__sbox_inst_com_y_inst_n483,
         round_inst_S_5__sbox_inst_com_y_inst_n482,
         round_inst_S_5__sbox_inst_com_y_inst_n481,
         round_inst_S_5__sbox_inst_com_y_inst_n480,
         round_inst_S_5__sbox_inst_com_y_inst_n479,
         round_inst_S_5__sbox_inst_com_y_inst_n478,
         round_inst_S_5__sbox_inst_com_y_inst_n477,
         round_inst_S_5__sbox_inst_com_y_inst_n476,
         round_inst_S_5__sbox_inst_com_y_inst_n475,
         round_inst_S_5__sbox_inst_com_y_inst_n474,
         round_inst_S_5__sbox_inst_com_y_inst_n473,
         round_inst_S_5__sbox_inst_com_y_inst_n472,
         round_inst_S_5__sbox_inst_com_y_inst_n471,
         round_inst_S_5__sbox_inst_com_y_inst_n470,
         round_inst_S_5__sbox_inst_com_y_inst_n469,
         round_inst_S_5__sbox_inst_com_y_inst_n468,
         round_inst_S_5__sbox_inst_com_y_inst_n467,
         round_inst_S_5__sbox_inst_com_y_inst_n466,
         round_inst_S_5__sbox_inst_com_y_inst_n465,
         round_inst_S_5__sbox_inst_com_y_inst_n464,
         round_inst_S_5__sbox_inst_com_y_inst_n463,
         round_inst_S_5__sbox_inst_com_y_inst_n462,
         round_inst_S_5__sbox_inst_com_y_inst_n461,
         round_inst_S_5__sbox_inst_com_y_inst_n460,
         round_inst_S_5__sbox_inst_com_y_inst_n459,
         round_inst_S_5__sbox_inst_com_y_inst_n458,
         round_inst_S_5__sbox_inst_com_y_inst_n457,
         round_inst_S_5__sbox_inst_com_y_inst_n456,
         round_inst_S_5__sbox_inst_com_y_inst_n455,
         round_inst_S_5__sbox_inst_com_y_inst_n454,
         round_inst_S_5__sbox_inst_com_y_inst_n453,
         round_inst_S_5__sbox_inst_com_y_inst_n452,
         round_inst_S_5__sbox_inst_com_y_inst_n451,
         round_inst_S_5__sbox_inst_com_y_inst_n450,
         round_inst_S_5__sbox_inst_com_y_inst_n449,
         round_inst_S_5__sbox_inst_com_y_inst_n448,
         round_inst_S_5__sbox_inst_com_y_inst_n447,
         round_inst_S_5__sbox_inst_com_y_inst_n446,
         round_inst_S_5__sbox_inst_com_y_inst_n445,
         round_inst_S_5__sbox_inst_com_y_inst_n444,
         round_inst_S_5__sbox_inst_com_y_inst_n443,
         round_inst_S_5__sbox_inst_com_y_inst_n442,
         round_inst_S_5__sbox_inst_com_y_inst_n441,
         round_inst_S_5__sbox_inst_com_y_inst_n440,
         round_inst_S_5__sbox_inst_com_y_inst_n439,
         round_inst_S_5__sbox_inst_com_y_inst_n438,
         round_inst_S_5__sbox_inst_com_y_inst_n437,
         round_inst_S_5__sbox_inst_com_y_inst_n436,
         round_inst_S_5__sbox_inst_com_y_inst_n435,
         round_inst_S_5__sbox_inst_com_y_inst_n434,
         round_inst_S_5__sbox_inst_com_y_inst_n433,
         round_inst_S_5__sbox_inst_com_y_inst_n432,
         round_inst_S_5__sbox_inst_com_y_inst_n431,
         round_inst_S_5__sbox_inst_com_y_inst_n430,
         round_inst_S_5__sbox_inst_com_y_inst_n429,
         round_inst_S_5__sbox_inst_com_y_inst_n428,
         round_inst_S_5__sbox_inst_com_y_inst_n427,
         round_inst_S_5__sbox_inst_com_y_inst_n426,
         round_inst_S_5__sbox_inst_com_y_inst_n425,
         round_inst_S_5__sbox_inst_com_y_inst_n424,
         round_inst_S_5__sbox_inst_com_y_inst_n423,
         round_inst_S_5__sbox_inst_com_y_inst_n422,
         round_inst_S_5__sbox_inst_com_y_inst_n421,
         round_inst_S_5__sbox_inst_com_y_inst_n420,
         round_inst_S_5__sbox_inst_com_y_inst_n419,
         round_inst_S_5__sbox_inst_com_y_inst_n418,
         round_inst_S_5__sbox_inst_com_y_inst_n417,
         round_inst_S_5__sbox_inst_com_y_inst_n416,
         round_inst_S_5__sbox_inst_com_y_inst_n415,
         round_inst_S_5__sbox_inst_com_y_inst_n414,
         round_inst_S_5__sbox_inst_com_y_inst_n413,
         round_inst_S_5__sbox_inst_com_y_inst_n412,
         round_inst_S_5__sbox_inst_com_y_inst_n411,
         round_inst_S_5__sbox_inst_com_y_inst_n410,
         round_inst_S_5__sbox_inst_com_y_inst_n409,
         round_inst_S_5__sbox_inst_com_y_inst_n408,
         round_inst_S_5__sbox_inst_com_y_inst_n407,
         round_inst_S_5__sbox_inst_com_y_inst_n406,
         round_inst_S_5__sbox_inst_com_y_inst_n405,
         round_inst_S_5__sbox_inst_com_y_inst_n404,
         round_inst_S_5__sbox_inst_com_y_inst_n403,
         round_inst_S_5__sbox_inst_com_y_inst_n402,
         round_inst_S_5__sbox_inst_com_y_inst_n401,
         round_inst_S_5__sbox_inst_com_y_inst_n400,
         round_inst_S_5__sbox_inst_com_y_inst_n399,
         round_inst_S_5__sbox_inst_com_y_inst_n398,
         round_inst_S_5__sbox_inst_com_y_inst_n397,
         round_inst_S_5__sbox_inst_com_y_inst_n396,
         round_inst_S_5__sbox_inst_com_y_inst_n395,
         round_inst_S_5__sbox_inst_com_y_inst_n394,
         round_inst_S_5__sbox_inst_com_y_inst_n393,
         round_inst_S_5__sbox_inst_com_y_inst_n392,
         round_inst_S_5__sbox_inst_com_y_inst_n391,
         round_inst_S_5__sbox_inst_com_y_inst_n390,
         round_inst_S_5__sbox_inst_com_y_inst_n389,
         round_inst_S_5__sbox_inst_com_y_inst_n388,
         round_inst_S_5__sbox_inst_com_y_inst_n387,
         round_inst_S_5__sbox_inst_com_y_inst_n386,
         round_inst_S_5__sbox_inst_com_z_inst_n516,
         round_inst_S_5__sbox_inst_com_z_inst_n515,
         round_inst_S_5__sbox_inst_com_z_inst_n514,
         round_inst_S_5__sbox_inst_com_z_inst_n513,
         round_inst_S_5__sbox_inst_com_z_inst_n512,
         round_inst_S_5__sbox_inst_com_z_inst_n511,
         round_inst_S_5__sbox_inst_com_z_inst_n510,
         round_inst_S_5__sbox_inst_com_z_inst_n509,
         round_inst_S_5__sbox_inst_com_z_inst_n508,
         round_inst_S_5__sbox_inst_com_z_inst_n507,
         round_inst_S_5__sbox_inst_com_z_inst_n506,
         round_inst_S_5__sbox_inst_com_z_inst_n505,
         round_inst_S_5__sbox_inst_com_z_inst_n504,
         round_inst_S_5__sbox_inst_com_z_inst_n503,
         round_inst_S_5__sbox_inst_com_z_inst_n502,
         round_inst_S_5__sbox_inst_com_z_inst_n501,
         round_inst_S_5__sbox_inst_com_z_inst_n500,
         round_inst_S_5__sbox_inst_com_z_inst_n499,
         round_inst_S_5__sbox_inst_com_z_inst_n498,
         round_inst_S_5__sbox_inst_com_z_inst_n497,
         round_inst_S_5__sbox_inst_com_z_inst_n496,
         round_inst_S_5__sbox_inst_com_z_inst_n495,
         round_inst_S_5__sbox_inst_com_z_inst_n494,
         round_inst_S_5__sbox_inst_com_z_inst_n493,
         round_inst_S_5__sbox_inst_com_z_inst_n492,
         round_inst_S_5__sbox_inst_com_z_inst_n491,
         round_inst_S_5__sbox_inst_com_z_inst_n490,
         round_inst_S_5__sbox_inst_com_z_inst_n489,
         round_inst_S_5__sbox_inst_com_z_inst_n488,
         round_inst_S_5__sbox_inst_com_z_inst_n487,
         round_inst_S_5__sbox_inst_com_z_inst_n486,
         round_inst_S_5__sbox_inst_com_z_inst_n485,
         round_inst_S_5__sbox_inst_com_z_inst_n484,
         round_inst_S_5__sbox_inst_com_z_inst_n483,
         round_inst_S_5__sbox_inst_com_z_inst_n482,
         round_inst_S_5__sbox_inst_com_z_inst_n481,
         round_inst_S_5__sbox_inst_com_z_inst_n480,
         round_inst_S_5__sbox_inst_com_z_inst_n479,
         round_inst_S_5__sbox_inst_com_z_inst_n478,
         round_inst_S_5__sbox_inst_com_z_inst_n477,
         round_inst_S_5__sbox_inst_com_z_inst_n476,
         round_inst_S_5__sbox_inst_com_z_inst_n475,
         round_inst_S_5__sbox_inst_com_z_inst_n474,
         round_inst_S_5__sbox_inst_com_z_inst_n473,
         round_inst_S_5__sbox_inst_com_z_inst_n472,
         round_inst_S_5__sbox_inst_com_z_inst_n471,
         round_inst_S_5__sbox_inst_com_z_inst_n470,
         round_inst_S_5__sbox_inst_com_z_inst_n469,
         round_inst_S_5__sbox_inst_com_z_inst_n468,
         round_inst_S_5__sbox_inst_com_z_inst_n467,
         round_inst_S_5__sbox_inst_com_z_inst_n466,
         round_inst_S_5__sbox_inst_com_z_inst_n465,
         round_inst_S_5__sbox_inst_com_z_inst_n464,
         round_inst_S_5__sbox_inst_com_z_inst_n463,
         round_inst_S_5__sbox_inst_com_z_inst_n462,
         round_inst_S_5__sbox_inst_com_z_inst_n461,
         round_inst_S_5__sbox_inst_com_z_inst_n460,
         round_inst_S_5__sbox_inst_com_z_inst_n459,
         round_inst_S_5__sbox_inst_com_z_inst_n458,
         round_inst_S_5__sbox_inst_com_z_inst_n457,
         round_inst_S_5__sbox_inst_com_z_inst_n456,
         round_inst_S_5__sbox_inst_com_z_inst_n455,
         round_inst_S_5__sbox_inst_com_z_inst_n454,
         round_inst_S_5__sbox_inst_com_z_inst_n453,
         round_inst_S_5__sbox_inst_com_z_inst_n452,
         round_inst_S_5__sbox_inst_com_z_inst_n451,
         round_inst_S_5__sbox_inst_com_z_inst_n450,
         round_inst_S_5__sbox_inst_com_z_inst_n449,
         round_inst_S_5__sbox_inst_com_z_inst_n448,
         round_inst_S_5__sbox_inst_com_z_inst_n447,
         round_inst_S_5__sbox_inst_com_z_inst_n446,
         round_inst_S_5__sbox_inst_com_z_inst_n445,
         round_inst_S_5__sbox_inst_com_z_inst_n444,
         round_inst_S_5__sbox_inst_com_z_inst_n443,
         round_inst_S_5__sbox_inst_com_z_inst_n442,
         round_inst_S_5__sbox_inst_com_z_inst_n441,
         round_inst_S_5__sbox_inst_com_z_inst_n440,
         round_inst_S_5__sbox_inst_com_z_inst_n439,
         round_inst_S_5__sbox_inst_com_z_inst_n438,
         round_inst_S_5__sbox_inst_com_z_inst_n437,
         round_inst_S_5__sbox_inst_com_z_inst_n436,
         round_inst_S_5__sbox_inst_com_z_inst_n435,
         round_inst_S_5__sbox_inst_com_z_inst_n434,
         round_inst_S_5__sbox_inst_com_z_inst_n433,
         round_inst_S_5__sbox_inst_com_z_inst_n432,
         round_inst_S_5__sbox_inst_com_z_inst_n431,
         round_inst_S_5__sbox_inst_com_z_inst_n430,
         round_inst_S_5__sbox_inst_com_z_inst_n429,
         round_inst_S_5__sbox_inst_com_z_inst_n428,
         round_inst_S_5__sbox_inst_com_z_inst_n427,
         round_inst_S_5__sbox_inst_com_z_inst_n426,
         round_inst_S_5__sbox_inst_com_z_inst_n425,
         round_inst_S_5__sbox_inst_com_z_inst_n424,
         round_inst_S_5__sbox_inst_com_z_inst_n423,
         round_inst_S_5__sbox_inst_com_z_inst_n422,
         round_inst_S_5__sbox_inst_com_z_inst_n421,
         round_inst_S_5__sbox_inst_com_z_inst_n420,
         round_inst_S_5__sbox_inst_com_z_inst_n419,
         round_inst_S_5__sbox_inst_com_z_inst_n418,
         round_inst_S_5__sbox_inst_com_z_inst_n417,
         round_inst_S_5__sbox_inst_com_z_inst_n416,
         round_inst_S_5__sbox_inst_com_z_inst_n415,
         round_inst_S_5__sbox_inst_com_z_inst_n414,
         round_inst_S_5__sbox_inst_com_z_inst_n413,
         round_inst_S_5__sbox_inst_com_z_inst_n412,
         round_inst_S_5__sbox_inst_com_z_inst_n411,
         round_inst_S_5__sbox_inst_com_z_inst_n410,
         round_inst_S_5__sbox_inst_com_z_inst_n409,
         round_inst_S_5__sbox_inst_com_z_inst_n408,
         round_inst_S_5__sbox_inst_com_z_inst_n407,
         round_inst_S_5__sbox_inst_com_z_inst_n406,
         round_inst_S_5__sbox_inst_com_z_inst_n405,
         round_inst_S_5__sbox_inst_com_z_inst_n404,
         round_inst_S_5__sbox_inst_com_z_inst_n403,
         round_inst_S_5__sbox_inst_com_z_inst_n402,
         round_inst_S_5__sbox_inst_com_z_inst_n401,
         round_inst_S_5__sbox_inst_com_z_inst_n400,
         round_inst_S_5__sbox_inst_com_z_inst_n399,
         round_inst_S_5__sbox_inst_com_z_inst_n398,
         round_inst_S_5__sbox_inst_com_z_inst_n397,
         round_inst_S_5__sbox_inst_com_z_inst_n396,
         round_inst_S_5__sbox_inst_com_z_inst_n395,
         round_inst_S_5__sbox_inst_com_z_inst_n394,
         round_inst_S_5__sbox_inst_com_z_inst_n393,
         round_inst_S_5__sbox_inst_com_z_inst_n392,
         round_inst_S_5__sbox_inst_com_z_inst_n391,
         round_inst_S_5__sbox_inst_com_z_inst_n390,
         round_inst_S_6__sbox_inst_n6, round_inst_S_6__sbox_inst_n5,
         round_inst_S_6__sbox_inst_n4, round_inst_S_6__sbox_inst_n3,
         round_inst_S_6__sbox_inst_n2, round_inst_S_6__sbox_inst_n1,
         round_inst_S_6__sbox_inst_com_w_inst_n532,
         round_inst_S_6__sbox_inst_com_w_inst_n531,
         round_inst_S_6__sbox_inst_com_w_inst_n530,
         round_inst_S_6__sbox_inst_com_w_inst_n529,
         round_inst_S_6__sbox_inst_com_w_inst_n528,
         round_inst_S_6__sbox_inst_com_w_inst_n527,
         round_inst_S_6__sbox_inst_com_w_inst_n526,
         round_inst_S_6__sbox_inst_com_w_inst_n525,
         round_inst_S_6__sbox_inst_com_w_inst_n524,
         round_inst_S_6__sbox_inst_com_w_inst_n523,
         round_inst_S_6__sbox_inst_com_w_inst_n522,
         round_inst_S_6__sbox_inst_com_w_inst_n521,
         round_inst_S_6__sbox_inst_com_w_inst_n520,
         round_inst_S_6__sbox_inst_com_w_inst_n519,
         round_inst_S_6__sbox_inst_com_w_inst_n518,
         round_inst_S_6__sbox_inst_com_w_inst_n517,
         round_inst_S_6__sbox_inst_com_w_inst_n516,
         round_inst_S_6__sbox_inst_com_w_inst_n515,
         round_inst_S_6__sbox_inst_com_w_inst_n514,
         round_inst_S_6__sbox_inst_com_w_inst_n513,
         round_inst_S_6__sbox_inst_com_w_inst_n512,
         round_inst_S_6__sbox_inst_com_w_inst_n511,
         round_inst_S_6__sbox_inst_com_w_inst_n510,
         round_inst_S_6__sbox_inst_com_w_inst_n509,
         round_inst_S_6__sbox_inst_com_w_inst_n508,
         round_inst_S_6__sbox_inst_com_w_inst_n507,
         round_inst_S_6__sbox_inst_com_w_inst_n506,
         round_inst_S_6__sbox_inst_com_w_inst_n505,
         round_inst_S_6__sbox_inst_com_w_inst_n504,
         round_inst_S_6__sbox_inst_com_w_inst_n503,
         round_inst_S_6__sbox_inst_com_w_inst_n502,
         round_inst_S_6__sbox_inst_com_w_inst_n501,
         round_inst_S_6__sbox_inst_com_w_inst_n500,
         round_inst_S_6__sbox_inst_com_w_inst_n499,
         round_inst_S_6__sbox_inst_com_w_inst_n498,
         round_inst_S_6__sbox_inst_com_w_inst_n497,
         round_inst_S_6__sbox_inst_com_w_inst_n496,
         round_inst_S_6__sbox_inst_com_w_inst_n495,
         round_inst_S_6__sbox_inst_com_w_inst_n494,
         round_inst_S_6__sbox_inst_com_w_inst_n493,
         round_inst_S_6__sbox_inst_com_w_inst_n492,
         round_inst_S_6__sbox_inst_com_w_inst_n491,
         round_inst_S_6__sbox_inst_com_w_inst_n490,
         round_inst_S_6__sbox_inst_com_w_inst_n489,
         round_inst_S_6__sbox_inst_com_w_inst_n488,
         round_inst_S_6__sbox_inst_com_w_inst_n487,
         round_inst_S_6__sbox_inst_com_w_inst_n486,
         round_inst_S_6__sbox_inst_com_w_inst_n485,
         round_inst_S_6__sbox_inst_com_w_inst_n484,
         round_inst_S_6__sbox_inst_com_w_inst_n483,
         round_inst_S_6__sbox_inst_com_w_inst_n482,
         round_inst_S_6__sbox_inst_com_w_inst_n481,
         round_inst_S_6__sbox_inst_com_w_inst_n480,
         round_inst_S_6__sbox_inst_com_w_inst_n479,
         round_inst_S_6__sbox_inst_com_w_inst_n478,
         round_inst_S_6__sbox_inst_com_w_inst_n477,
         round_inst_S_6__sbox_inst_com_w_inst_n476,
         round_inst_S_6__sbox_inst_com_w_inst_n475,
         round_inst_S_6__sbox_inst_com_w_inst_n474,
         round_inst_S_6__sbox_inst_com_w_inst_n473,
         round_inst_S_6__sbox_inst_com_w_inst_n472,
         round_inst_S_6__sbox_inst_com_w_inst_n471,
         round_inst_S_6__sbox_inst_com_w_inst_n470,
         round_inst_S_6__sbox_inst_com_w_inst_n469,
         round_inst_S_6__sbox_inst_com_w_inst_n468,
         round_inst_S_6__sbox_inst_com_w_inst_n467,
         round_inst_S_6__sbox_inst_com_w_inst_n466,
         round_inst_S_6__sbox_inst_com_w_inst_n465,
         round_inst_S_6__sbox_inst_com_w_inst_n464,
         round_inst_S_6__sbox_inst_com_w_inst_n463,
         round_inst_S_6__sbox_inst_com_w_inst_n462,
         round_inst_S_6__sbox_inst_com_w_inst_n461,
         round_inst_S_6__sbox_inst_com_w_inst_n460,
         round_inst_S_6__sbox_inst_com_w_inst_n459,
         round_inst_S_6__sbox_inst_com_w_inst_n458,
         round_inst_S_6__sbox_inst_com_w_inst_n457,
         round_inst_S_6__sbox_inst_com_w_inst_n456,
         round_inst_S_6__sbox_inst_com_w_inst_n455,
         round_inst_S_6__sbox_inst_com_w_inst_n454,
         round_inst_S_6__sbox_inst_com_w_inst_n453,
         round_inst_S_6__sbox_inst_com_w_inst_n452,
         round_inst_S_6__sbox_inst_com_w_inst_n451,
         round_inst_S_6__sbox_inst_com_w_inst_n450,
         round_inst_S_6__sbox_inst_com_w_inst_n449,
         round_inst_S_6__sbox_inst_com_w_inst_n448,
         round_inst_S_6__sbox_inst_com_w_inst_n447,
         round_inst_S_6__sbox_inst_com_w_inst_n446,
         round_inst_S_6__sbox_inst_com_w_inst_n445,
         round_inst_S_6__sbox_inst_com_w_inst_n444,
         round_inst_S_6__sbox_inst_com_w_inst_n443,
         round_inst_S_6__sbox_inst_com_w_inst_n442,
         round_inst_S_6__sbox_inst_com_w_inst_n441,
         round_inst_S_6__sbox_inst_com_w_inst_n440,
         round_inst_S_6__sbox_inst_com_w_inst_n439,
         round_inst_S_6__sbox_inst_com_w_inst_n438,
         round_inst_S_6__sbox_inst_com_w_inst_n437,
         round_inst_S_6__sbox_inst_com_w_inst_n436,
         round_inst_S_6__sbox_inst_com_w_inst_n435,
         round_inst_S_6__sbox_inst_com_w_inst_n434,
         round_inst_S_6__sbox_inst_com_w_inst_n433,
         round_inst_S_6__sbox_inst_com_w_inst_n432,
         round_inst_S_6__sbox_inst_com_w_inst_n431,
         round_inst_S_6__sbox_inst_com_w_inst_n430,
         round_inst_S_6__sbox_inst_com_w_inst_n429,
         round_inst_S_6__sbox_inst_com_w_inst_n428,
         round_inst_S_6__sbox_inst_com_w_inst_n427,
         round_inst_S_6__sbox_inst_com_w_inst_n426,
         round_inst_S_6__sbox_inst_com_w_inst_n425,
         round_inst_S_6__sbox_inst_com_w_inst_n424,
         round_inst_S_6__sbox_inst_com_w_inst_n423,
         round_inst_S_6__sbox_inst_com_w_inst_n422,
         round_inst_S_6__sbox_inst_com_w_inst_n421,
         round_inst_S_6__sbox_inst_com_w_inst_n420,
         round_inst_S_6__sbox_inst_com_w_inst_n419,
         round_inst_S_6__sbox_inst_com_w_inst_n418,
         round_inst_S_6__sbox_inst_com_w_inst_n417,
         round_inst_S_6__sbox_inst_com_w_inst_n416,
         round_inst_S_6__sbox_inst_com_w_inst_n415,
         round_inst_S_6__sbox_inst_com_w_inst_n414,
         round_inst_S_6__sbox_inst_com_w_inst_n413,
         round_inst_S_6__sbox_inst_com_w_inst_n412,
         round_inst_S_6__sbox_inst_com_w_inst_n411,
         round_inst_S_6__sbox_inst_com_w_inst_n410,
         round_inst_S_6__sbox_inst_com_w_inst_n409,
         round_inst_S_6__sbox_inst_com_w_inst_n408,
         round_inst_S_6__sbox_inst_com_w_inst_n407,
         round_inst_S_6__sbox_inst_com_w_inst_n406,
         round_inst_S_6__sbox_inst_com_w_inst_n405,
         round_inst_S_6__sbox_inst_com_w_inst_n404,
         round_inst_S_6__sbox_inst_com_w_inst_n403,
         round_inst_S_6__sbox_inst_com_w_inst_n402,
         round_inst_S_6__sbox_inst_com_w_inst_n401,
         round_inst_S_6__sbox_inst_com_w_inst_n400,
         round_inst_S_6__sbox_inst_com_w_inst_n399,
         round_inst_S_6__sbox_inst_com_w_inst_n398,
         round_inst_S_6__sbox_inst_com_w_inst_n397,
         round_inst_S_6__sbox_inst_com_w_inst_n396,
         round_inst_S_6__sbox_inst_com_x_inst_n511,
         round_inst_S_6__sbox_inst_com_x_inst_n510,
         round_inst_S_6__sbox_inst_com_x_inst_n509,
         round_inst_S_6__sbox_inst_com_x_inst_n508,
         round_inst_S_6__sbox_inst_com_x_inst_n507,
         round_inst_S_6__sbox_inst_com_x_inst_n506,
         round_inst_S_6__sbox_inst_com_x_inst_n505,
         round_inst_S_6__sbox_inst_com_x_inst_n504,
         round_inst_S_6__sbox_inst_com_x_inst_n503,
         round_inst_S_6__sbox_inst_com_x_inst_n502,
         round_inst_S_6__sbox_inst_com_x_inst_n501,
         round_inst_S_6__sbox_inst_com_x_inst_n500,
         round_inst_S_6__sbox_inst_com_x_inst_n499,
         round_inst_S_6__sbox_inst_com_x_inst_n498,
         round_inst_S_6__sbox_inst_com_x_inst_n497,
         round_inst_S_6__sbox_inst_com_x_inst_n496,
         round_inst_S_6__sbox_inst_com_x_inst_n495,
         round_inst_S_6__sbox_inst_com_x_inst_n494,
         round_inst_S_6__sbox_inst_com_x_inst_n493,
         round_inst_S_6__sbox_inst_com_x_inst_n492,
         round_inst_S_6__sbox_inst_com_x_inst_n491,
         round_inst_S_6__sbox_inst_com_x_inst_n490,
         round_inst_S_6__sbox_inst_com_x_inst_n489,
         round_inst_S_6__sbox_inst_com_x_inst_n488,
         round_inst_S_6__sbox_inst_com_x_inst_n487,
         round_inst_S_6__sbox_inst_com_x_inst_n486,
         round_inst_S_6__sbox_inst_com_x_inst_n485,
         round_inst_S_6__sbox_inst_com_x_inst_n484,
         round_inst_S_6__sbox_inst_com_x_inst_n483,
         round_inst_S_6__sbox_inst_com_x_inst_n482,
         round_inst_S_6__sbox_inst_com_x_inst_n481,
         round_inst_S_6__sbox_inst_com_x_inst_n480,
         round_inst_S_6__sbox_inst_com_x_inst_n479,
         round_inst_S_6__sbox_inst_com_x_inst_n478,
         round_inst_S_6__sbox_inst_com_x_inst_n477,
         round_inst_S_6__sbox_inst_com_x_inst_n476,
         round_inst_S_6__sbox_inst_com_x_inst_n475,
         round_inst_S_6__sbox_inst_com_x_inst_n474,
         round_inst_S_6__sbox_inst_com_x_inst_n473,
         round_inst_S_6__sbox_inst_com_x_inst_n472,
         round_inst_S_6__sbox_inst_com_x_inst_n471,
         round_inst_S_6__sbox_inst_com_x_inst_n470,
         round_inst_S_6__sbox_inst_com_x_inst_n469,
         round_inst_S_6__sbox_inst_com_x_inst_n468,
         round_inst_S_6__sbox_inst_com_x_inst_n467,
         round_inst_S_6__sbox_inst_com_x_inst_n466,
         round_inst_S_6__sbox_inst_com_x_inst_n465,
         round_inst_S_6__sbox_inst_com_x_inst_n464,
         round_inst_S_6__sbox_inst_com_x_inst_n463,
         round_inst_S_6__sbox_inst_com_x_inst_n462,
         round_inst_S_6__sbox_inst_com_x_inst_n461,
         round_inst_S_6__sbox_inst_com_x_inst_n460,
         round_inst_S_6__sbox_inst_com_x_inst_n459,
         round_inst_S_6__sbox_inst_com_x_inst_n458,
         round_inst_S_6__sbox_inst_com_x_inst_n457,
         round_inst_S_6__sbox_inst_com_x_inst_n456,
         round_inst_S_6__sbox_inst_com_x_inst_n455,
         round_inst_S_6__sbox_inst_com_x_inst_n454,
         round_inst_S_6__sbox_inst_com_x_inst_n453,
         round_inst_S_6__sbox_inst_com_x_inst_n452,
         round_inst_S_6__sbox_inst_com_x_inst_n451,
         round_inst_S_6__sbox_inst_com_x_inst_n450,
         round_inst_S_6__sbox_inst_com_x_inst_n449,
         round_inst_S_6__sbox_inst_com_x_inst_n448,
         round_inst_S_6__sbox_inst_com_x_inst_n447,
         round_inst_S_6__sbox_inst_com_x_inst_n446,
         round_inst_S_6__sbox_inst_com_x_inst_n445,
         round_inst_S_6__sbox_inst_com_x_inst_n444,
         round_inst_S_6__sbox_inst_com_x_inst_n443,
         round_inst_S_6__sbox_inst_com_x_inst_n442,
         round_inst_S_6__sbox_inst_com_x_inst_n441,
         round_inst_S_6__sbox_inst_com_x_inst_n440,
         round_inst_S_6__sbox_inst_com_x_inst_n439,
         round_inst_S_6__sbox_inst_com_x_inst_n438,
         round_inst_S_6__sbox_inst_com_x_inst_n437,
         round_inst_S_6__sbox_inst_com_x_inst_n436,
         round_inst_S_6__sbox_inst_com_x_inst_n435,
         round_inst_S_6__sbox_inst_com_x_inst_n434,
         round_inst_S_6__sbox_inst_com_x_inst_n433,
         round_inst_S_6__sbox_inst_com_x_inst_n432,
         round_inst_S_6__sbox_inst_com_x_inst_n431,
         round_inst_S_6__sbox_inst_com_x_inst_n430,
         round_inst_S_6__sbox_inst_com_x_inst_n429,
         round_inst_S_6__sbox_inst_com_x_inst_n428,
         round_inst_S_6__sbox_inst_com_x_inst_n427,
         round_inst_S_6__sbox_inst_com_x_inst_n426,
         round_inst_S_6__sbox_inst_com_x_inst_n425,
         round_inst_S_6__sbox_inst_com_x_inst_n424,
         round_inst_S_6__sbox_inst_com_x_inst_n423,
         round_inst_S_6__sbox_inst_com_x_inst_n422,
         round_inst_S_6__sbox_inst_com_x_inst_n421,
         round_inst_S_6__sbox_inst_com_x_inst_n420,
         round_inst_S_6__sbox_inst_com_x_inst_n419,
         round_inst_S_6__sbox_inst_com_x_inst_n418,
         round_inst_S_6__sbox_inst_com_x_inst_n417,
         round_inst_S_6__sbox_inst_com_x_inst_n416,
         round_inst_S_6__sbox_inst_com_x_inst_n415,
         round_inst_S_6__sbox_inst_com_x_inst_n414,
         round_inst_S_6__sbox_inst_com_x_inst_n413,
         round_inst_S_6__sbox_inst_com_x_inst_n412,
         round_inst_S_6__sbox_inst_com_x_inst_n411,
         round_inst_S_6__sbox_inst_com_x_inst_n410,
         round_inst_S_6__sbox_inst_com_x_inst_n409,
         round_inst_S_6__sbox_inst_com_x_inst_n408,
         round_inst_S_6__sbox_inst_com_x_inst_n407,
         round_inst_S_6__sbox_inst_com_x_inst_n406,
         round_inst_S_6__sbox_inst_com_x_inst_n405,
         round_inst_S_6__sbox_inst_com_x_inst_n404,
         round_inst_S_6__sbox_inst_com_x_inst_n403,
         round_inst_S_6__sbox_inst_com_x_inst_n402,
         round_inst_S_6__sbox_inst_com_x_inst_n401,
         round_inst_S_6__sbox_inst_com_x_inst_n400,
         round_inst_S_6__sbox_inst_com_x_inst_n399,
         round_inst_S_6__sbox_inst_com_x_inst_n398,
         round_inst_S_6__sbox_inst_com_x_inst_n397,
         round_inst_S_6__sbox_inst_com_x_inst_n396,
         round_inst_S_6__sbox_inst_com_x_inst_n395,
         round_inst_S_6__sbox_inst_com_x_inst_n394,
         round_inst_S_6__sbox_inst_com_x_inst_n393,
         round_inst_S_6__sbox_inst_com_x_inst_n392,
         round_inst_S_6__sbox_inst_com_x_inst_n391,
         round_inst_S_6__sbox_inst_com_x_inst_n390,
         round_inst_S_6__sbox_inst_com_x_inst_n389,
         round_inst_S_6__sbox_inst_com_x_inst_n388,
         round_inst_S_6__sbox_inst_com_x_inst_n387,
         round_inst_S_6__sbox_inst_com_x_inst_n386,
         round_inst_S_6__sbox_inst_com_x_inst_n385,
         round_inst_S_6__sbox_inst_com_x_inst_n384,
         round_inst_S_6__sbox_inst_com_x_inst_n383,
         round_inst_S_6__sbox_inst_com_x_inst_n382,
         round_inst_S_6__sbox_inst_com_x_inst_n381,
         round_inst_S_6__sbox_inst_com_y_inst_n518,
         round_inst_S_6__sbox_inst_com_y_inst_n517,
         round_inst_S_6__sbox_inst_com_y_inst_n516,
         round_inst_S_6__sbox_inst_com_y_inst_n515,
         round_inst_S_6__sbox_inst_com_y_inst_n514,
         round_inst_S_6__sbox_inst_com_y_inst_n513,
         round_inst_S_6__sbox_inst_com_y_inst_n512,
         round_inst_S_6__sbox_inst_com_y_inst_n511,
         round_inst_S_6__sbox_inst_com_y_inst_n510,
         round_inst_S_6__sbox_inst_com_y_inst_n509,
         round_inst_S_6__sbox_inst_com_y_inst_n508,
         round_inst_S_6__sbox_inst_com_y_inst_n507,
         round_inst_S_6__sbox_inst_com_y_inst_n506,
         round_inst_S_6__sbox_inst_com_y_inst_n505,
         round_inst_S_6__sbox_inst_com_y_inst_n504,
         round_inst_S_6__sbox_inst_com_y_inst_n503,
         round_inst_S_6__sbox_inst_com_y_inst_n502,
         round_inst_S_6__sbox_inst_com_y_inst_n501,
         round_inst_S_6__sbox_inst_com_y_inst_n500,
         round_inst_S_6__sbox_inst_com_y_inst_n499,
         round_inst_S_6__sbox_inst_com_y_inst_n498,
         round_inst_S_6__sbox_inst_com_y_inst_n497,
         round_inst_S_6__sbox_inst_com_y_inst_n496,
         round_inst_S_6__sbox_inst_com_y_inst_n495,
         round_inst_S_6__sbox_inst_com_y_inst_n494,
         round_inst_S_6__sbox_inst_com_y_inst_n493,
         round_inst_S_6__sbox_inst_com_y_inst_n492,
         round_inst_S_6__sbox_inst_com_y_inst_n491,
         round_inst_S_6__sbox_inst_com_y_inst_n490,
         round_inst_S_6__sbox_inst_com_y_inst_n489,
         round_inst_S_6__sbox_inst_com_y_inst_n488,
         round_inst_S_6__sbox_inst_com_y_inst_n487,
         round_inst_S_6__sbox_inst_com_y_inst_n486,
         round_inst_S_6__sbox_inst_com_y_inst_n485,
         round_inst_S_6__sbox_inst_com_y_inst_n484,
         round_inst_S_6__sbox_inst_com_y_inst_n483,
         round_inst_S_6__sbox_inst_com_y_inst_n482,
         round_inst_S_6__sbox_inst_com_y_inst_n481,
         round_inst_S_6__sbox_inst_com_y_inst_n480,
         round_inst_S_6__sbox_inst_com_y_inst_n479,
         round_inst_S_6__sbox_inst_com_y_inst_n478,
         round_inst_S_6__sbox_inst_com_y_inst_n477,
         round_inst_S_6__sbox_inst_com_y_inst_n476,
         round_inst_S_6__sbox_inst_com_y_inst_n475,
         round_inst_S_6__sbox_inst_com_y_inst_n474,
         round_inst_S_6__sbox_inst_com_y_inst_n473,
         round_inst_S_6__sbox_inst_com_y_inst_n472,
         round_inst_S_6__sbox_inst_com_y_inst_n471,
         round_inst_S_6__sbox_inst_com_y_inst_n470,
         round_inst_S_6__sbox_inst_com_y_inst_n469,
         round_inst_S_6__sbox_inst_com_y_inst_n468,
         round_inst_S_6__sbox_inst_com_y_inst_n467,
         round_inst_S_6__sbox_inst_com_y_inst_n466,
         round_inst_S_6__sbox_inst_com_y_inst_n465,
         round_inst_S_6__sbox_inst_com_y_inst_n464,
         round_inst_S_6__sbox_inst_com_y_inst_n463,
         round_inst_S_6__sbox_inst_com_y_inst_n462,
         round_inst_S_6__sbox_inst_com_y_inst_n461,
         round_inst_S_6__sbox_inst_com_y_inst_n460,
         round_inst_S_6__sbox_inst_com_y_inst_n459,
         round_inst_S_6__sbox_inst_com_y_inst_n458,
         round_inst_S_6__sbox_inst_com_y_inst_n457,
         round_inst_S_6__sbox_inst_com_y_inst_n456,
         round_inst_S_6__sbox_inst_com_y_inst_n455,
         round_inst_S_6__sbox_inst_com_y_inst_n454,
         round_inst_S_6__sbox_inst_com_y_inst_n453,
         round_inst_S_6__sbox_inst_com_y_inst_n452,
         round_inst_S_6__sbox_inst_com_y_inst_n451,
         round_inst_S_6__sbox_inst_com_y_inst_n450,
         round_inst_S_6__sbox_inst_com_y_inst_n449,
         round_inst_S_6__sbox_inst_com_y_inst_n448,
         round_inst_S_6__sbox_inst_com_y_inst_n447,
         round_inst_S_6__sbox_inst_com_y_inst_n446,
         round_inst_S_6__sbox_inst_com_y_inst_n445,
         round_inst_S_6__sbox_inst_com_y_inst_n444,
         round_inst_S_6__sbox_inst_com_y_inst_n443,
         round_inst_S_6__sbox_inst_com_y_inst_n442,
         round_inst_S_6__sbox_inst_com_y_inst_n441,
         round_inst_S_6__sbox_inst_com_y_inst_n440,
         round_inst_S_6__sbox_inst_com_y_inst_n439,
         round_inst_S_6__sbox_inst_com_y_inst_n438,
         round_inst_S_6__sbox_inst_com_y_inst_n437,
         round_inst_S_6__sbox_inst_com_y_inst_n436,
         round_inst_S_6__sbox_inst_com_y_inst_n435,
         round_inst_S_6__sbox_inst_com_y_inst_n434,
         round_inst_S_6__sbox_inst_com_y_inst_n433,
         round_inst_S_6__sbox_inst_com_y_inst_n432,
         round_inst_S_6__sbox_inst_com_y_inst_n431,
         round_inst_S_6__sbox_inst_com_y_inst_n430,
         round_inst_S_6__sbox_inst_com_y_inst_n429,
         round_inst_S_6__sbox_inst_com_y_inst_n428,
         round_inst_S_6__sbox_inst_com_y_inst_n427,
         round_inst_S_6__sbox_inst_com_y_inst_n426,
         round_inst_S_6__sbox_inst_com_y_inst_n425,
         round_inst_S_6__sbox_inst_com_y_inst_n424,
         round_inst_S_6__sbox_inst_com_y_inst_n423,
         round_inst_S_6__sbox_inst_com_y_inst_n422,
         round_inst_S_6__sbox_inst_com_y_inst_n421,
         round_inst_S_6__sbox_inst_com_y_inst_n420,
         round_inst_S_6__sbox_inst_com_y_inst_n419,
         round_inst_S_6__sbox_inst_com_y_inst_n418,
         round_inst_S_6__sbox_inst_com_y_inst_n417,
         round_inst_S_6__sbox_inst_com_y_inst_n416,
         round_inst_S_6__sbox_inst_com_y_inst_n415,
         round_inst_S_6__sbox_inst_com_y_inst_n414,
         round_inst_S_6__sbox_inst_com_y_inst_n413,
         round_inst_S_6__sbox_inst_com_y_inst_n412,
         round_inst_S_6__sbox_inst_com_y_inst_n411,
         round_inst_S_6__sbox_inst_com_y_inst_n410,
         round_inst_S_6__sbox_inst_com_y_inst_n409,
         round_inst_S_6__sbox_inst_com_y_inst_n408,
         round_inst_S_6__sbox_inst_com_y_inst_n407,
         round_inst_S_6__sbox_inst_com_y_inst_n406,
         round_inst_S_6__sbox_inst_com_y_inst_n405,
         round_inst_S_6__sbox_inst_com_y_inst_n404,
         round_inst_S_6__sbox_inst_com_y_inst_n403,
         round_inst_S_6__sbox_inst_com_y_inst_n402,
         round_inst_S_6__sbox_inst_com_y_inst_n401,
         round_inst_S_6__sbox_inst_com_y_inst_n400,
         round_inst_S_6__sbox_inst_com_y_inst_n399,
         round_inst_S_6__sbox_inst_com_y_inst_n398,
         round_inst_S_6__sbox_inst_com_y_inst_n397,
         round_inst_S_6__sbox_inst_com_y_inst_n396,
         round_inst_S_6__sbox_inst_com_y_inst_n395,
         round_inst_S_6__sbox_inst_com_y_inst_n394,
         round_inst_S_6__sbox_inst_com_y_inst_n393,
         round_inst_S_6__sbox_inst_com_y_inst_n392,
         round_inst_S_6__sbox_inst_com_y_inst_n391,
         round_inst_S_6__sbox_inst_com_y_inst_n390,
         round_inst_S_6__sbox_inst_com_y_inst_n389,
         round_inst_S_6__sbox_inst_com_y_inst_n388,
         round_inst_S_6__sbox_inst_com_y_inst_n387,
         round_inst_S_6__sbox_inst_com_y_inst_n386,
         round_inst_S_6__sbox_inst_com_z_inst_n516,
         round_inst_S_6__sbox_inst_com_z_inst_n515,
         round_inst_S_6__sbox_inst_com_z_inst_n514,
         round_inst_S_6__sbox_inst_com_z_inst_n513,
         round_inst_S_6__sbox_inst_com_z_inst_n512,
         round_inst_S_6__sbox_inst_com_z_inst_n511,
         round_inst_S_6__sbox_inst_com_z_inst_n510,
         round_inst_S_6__sbox_inst_com_z_inst_n509,
         round_inst_S_6__sbox_inst_com_z_inst_n508,
         round_inst_S_6__sbox_inst_com_z_inst_n507,
         round_inst_S_6__sbox_inst_com_z_inst_n506,
         round_inst_S_6__sbox_inst_com_z_inst_n505,
         round_inst_S_6__sbox_inst_com_z_inst_n504,
         round_inst_S_6__sbox_inst_com_z_inst_n503,
         round_inst_S_6__sbox_inst_com_z_inst_n502,
         round_inst_S_6__sbox_inst_com_z_inst_n501,
         round_inst_S_6__sbox_inst_com_z_inst_n500,
         round_inst_S_6__sbox_inst_com_z_inst_n499,
         round_inst_S_6__sbox_inst_com_z_inst_n498,
         round_inst_S_6__sbox_inst_com_z_inst_n497,
         round_inst_S_6__sbox_inst_com_z_inst_n496,
         round_inst_S_6__sbox_inst_com_z_inst_n495,
         round_inst_S_6__sbox_inst_com_z_inst_n494,
         round_inst_S_6__sbox_inst_com_z_inst_n493,
         round_inst_S_6__sbox_inst_com_z_inst_n492,
         round_inst_S_6__sbox_inst_com_z_inst_n491,
         round_inst_S_6__sbox_inst_com_z_inst_n490,
         round_inst_S_6__sbox_inst_com_z_inst_n489,
         round_inst_S_6__sbox_inst_com_z_inst_n488,
         round_inst_S_6__sbox_inst_com_z_inst_n487,
         round_inst_S_6__sbox_inst_com_z_inst_n486,
         round_inst_S_6__sbox_inst_com_z_inst_n485,
         round_inst_S_6__sbox_inst_com_z_inst_n484,
         round_inst_S_6__sbox_inst_com_z_inst_n483,
         round_inst_S_6__sbox_inst_com_z_inst_n482,
         round_inst_S_6__sbox_inst_com_z_inst_n481,
         round_inst_S_6__sbox_inst_com_z_inst_n480,
         round_inst_S_6__sbox_inst_com_z_inst_n479,
         round_inst_S_6__sbox_inst_com_z_inst_n478,
         round_inst_S_6__sbox_inst_com_z_inst_n477,
         round_inst_S_6__sbox_inst_com_z_inst_n476,
         round_inst_S_6__sbox_inst_com_z_inst_n475,
         round_inst_S_6__sbox_inst_com_z_inst_n474,
         round_inst_S_6__sbox_inst_com_z_inst_n473,
         round_inst_S_6__sbox_inst_com_z_inst_n472,
         round_inst_S_6__sbox_inst_com_z_inst_n471,
         round_inst_S_6__sbox_inst_com_z_inst_n470,
         round_inst_S_6__sbox_inst_com_z_inst_n469,
         round_inst_S_6__sbox_inst_com_z_inst_n468,
         round_inst_S_6__sbox_inst_com_z_inst_n467,
         round_inst_S_6__sbox_inst_com_z_inst_n466,
         round_inst_S_6__sbox_inst_com_z_inst_n465,
         round_inst_S_6__sbox_inst_com_z_inst_n464,
         round_inst_S_6__sbox_inst_com_z_inst_n463,
         round_inst_S_6__sbox_inst_com_z_inst_n462,
         round_inst_S_6__sbox_inst_com_z_inst_n461,
         round_inst_S_6__sbox_inst_com_z_inst_n460,
         round_inst_S_6__sbox_inst_com_z_inst_n459,
         round_inst_S_6__sbox_inst_com_z_inst_n458,
         round_inst_S_6__sbox_inst_com_z_inst_n457,
         round_inst_S_6__sbox_inst_com_z_inst_n456,
         round_inst_S_6__sbox_inst_com_z_inst_n455,
         round_inst_S_6__sbox_inst_com_z_inst_n454,
         round_inst_S_6__sbox_inst_com_z_inst_n453,
         round_inst_S_6__sbox_inst_com_z_inst_n452,
         round_inst_S_6__sbox_inst_com_z_inst_n451,
         round_inst_S_6__sbox_inst_com_z_inst_n450,
         round_inst_S_6__sbox_inst_com_z_inst_n449,
         round_inst_S_6__sbox_inst_com_z_inst_n448,
         round_inst_S_6__sbox_inst_com_z_inst_n447,
         round_inst_S_6__sbox_inst_com_z_inst_n446,
         round_inst_S_6__sbox_inst_com_z_inst_n445,
         round_inst_S_6__sbox_inst_com_z_inst_n444,
         round_inst_S_6__sbox_inst_com_z_inst_n443,
         round_inst_S_6__sbox_inst_com_z_inst_n442,
         round_inst_S_6__sbox_inst_com_z_inst_n441,
         round_inst_S_6__sbox_inst_com_z_inst_n440,
         round_inst_S_6__sbox_inst_com_z_inst_n439,
         round_inst_S_6__sbox_inst_com_z_inst_n438,
         round_inst_S_6__sbox_inst_com_z_inst_n437,
         round_inst_S_6__sbox_inst_com_z_inst_n436,
         round_inst_S_6__sbox_inst_com_z_inst_n435,
         round_inst_S_6__sbox_inst_com_z_inst_n434,
         round_inst_S_6__sbox_inst_com_z_inst_n433,
         round_inst_S_6__sbox_inst_com_z_inst_n432,
         round_inst_S_6__sbox_inst_com_z_inst_n431,
         round_inst_S_6__sbox_inst_com_z_inst_n430,
         round_inst_S_6__sbox_inst_com_z_inst_n429,
         round_inst_S_6__sbox_inst_com_z_inst_n428,
         round_inst_S_6__sbox_inst_com_z_inst_n427,
         round_inst_S_6__sbox_inst_com_z_inst_n426,
         round_inst_S_6__sbox_inst_com_z_inst_n425,
         round_inst_S_6__sbox_inst_com_z_inst_n424,
         round_inst_S_6__sbox_inst_com_z_inst_n423,
         round_inst_S_6__sbox_inst_com_z_inst_n422,
         round_inst_S_6__sbox_inst_com_z_inst_n421,
         round_inst_S_6__sbox_inst_com_z_inst_n420,
         round_inst_S_6__sbox_inst_com_z_inst_n419,
         round_inst_S_6__sbox_inst_com_z_inst_n418,
         round_inst_S_6__sbox_inst_com_z_inst_n417,
         round_inst_S_6__sbox_inst_com_z_inst_n416,
         round_inst_S_6__sbox_inst_com_z_inst_n415,
         round_inst_S_6__sbox_inst_com_z_inst_n414,
         round_inst_S_6__sbox_inst_com_z_inst_n413,
         round_inst_S_6__sbox_inst_com_z_inst_n412,
         round_inst_S_6__sbox_inst_com_z_inst_n411,
         round_inst_S_6__sbox_inst_com_z_inst_n410,
         round_inst_S_6__sbox_inst_com_z_inst_n409,
         round_inst_S_6__sbox_inst_com_z_inst_n408,
         round_inst_S_6__sbox_inst_com_z_inst_n407,
         round_inst_S_6__sbox_inst_com_z_inst_n406,
         round_inst_S_6__sbox_inst_com_z_inst_n405,
         round_inst_S_6__sbox_inst_com_z_inst_n404,
         round_inst_S_6__sbox_inst_com_z_inst_n403,
         round_inst_S_6__sbox_inst_com_z_inst_n402,
         round_inst_S_6__sbox_inst_com_z_inst_n401,
         round_inst_S_6__sbox_inst_com_z_inst_n400,
         round_inst_S_6__sbox_inst_com_z_inst_n399,
         round_inst_S_6__sbox_inst_com_z_inst_n398,
         round_inst_S_6__sbox_inst_com_z_inst_n397,
         round_inst_S_6__sbox_inst_com_z_inst_n396,
         round_inst_S_6__sbox_inst_com_z_inst_n395,
         round_inst_S_6__sbox_inst_com_z_inst_n394,
         round_inst_S_6__sbox_inst_com_z_inst_n393,
         round_inst_S_6__sbox_inst_com_z_inst_n392,
         round_inst_S_6__sbox_inst_com_z_inst_n391,
         round_inst_S_6__sbox_inst_com_z_inst_n390,
         round_inst_S_7__sbox_inst_n6, round_inst_S_7__sbox_inst_n5,
         round_inst_S_7__sbox_inst_n4, round_inst_S_7__sbox_inst_n3,
         round_inst_S_7__sbox_inst_n2, round_inst_S_7__sbox_inst_n1,
         round_inst_S_7__sbox_inst_com_w_inst_n532,
         round_inst_S_7__sbox_inst_com_w_inst_n531,
         round_inst_S_7__sbox_inst_com_w_inst_n530,
         round_inst_S_7__sbox_inst_com_w_inst_n529,
         round_inst_S_7__sbox_inst_com_w_inst_n528,
         round_inst_S_7__sbox_inst_com_w_inst_n527,
         round_inst_S_7__sbox_inst_com_w_inst_n526,
         round_inst_S_7__sbox_inst_com_w_inst_n525,
         round_inst_S_7__sbox_inst_com_w_inst_n524,
         round_inst_S_7__sbox_inst_com_w_inst_n523,
         round_inst_S_7__sbox_inst_com_w_inst_n522,
         round_inst_S_7__sbox_inst_com_w_inst_n521,
         round_inst_S_7__sbox_inst_com_w_inst_n520,
         round_inst_S_7__sbox_inst_com_w_inst_n519,
         round_inst_S_7__sbox_inst_com_w_inst_n518,
         round_inst_S_7__sbox_inst_com_w_inst_n517,
         round_inst_S_7__sbox_inst_com_w_inst_n516,
         round_inst_S_7__sbox_inst_com_w_inst_n515,
         round_inst_S_7__sbox_inst_com_w_inst_n514,
         round_inst_S_7__sbox_inst_com_w_inst_n513,
         round_inst_S_7__sbox_inst_com_w_inst_n512,
         round_inst_S_7__sbox_inst_com_w_inst_n511,
         round_inst_S_7__sbox_inst_com_w_inst_n510,
         round_inst_S_7__sbox_inst_com_w_inst_n509,
         round_inst_S_7__sbox_inst_com_w_inst_n508,
         round_inst_S_7__sbox_inst_com_w_inst_n507,
         round_inst_S_7__sbox_inst_com_w_inst_n506,
         round_inst_S_7__sbox_inst_com_w_inst_n505,
         round_inst_S_7__sbox_inst_com_w_inst_n504,
         round_inst_S_7__sbox_inst_com_w_inst_n503,
         round_inst_S_7__sbox_inst_com_w_inst_n502,
         round_inst_S_7__sbox_inst_com_w_inst_n501,
         round_inst_S_7__sbox_inst_com_w_inst_n500,
         round_inst_S_7__sbox_inst_com_w_inst_n499,
         round_inst_S_7__sbox_inst_com_w_inst_n498,
         round_inst_S_7__sbox_inst_com_w_inst_n497,
         round_inst_S_7__sbox_inst_com_w_inst_n496,
         round_inst_S_7__sbox_inst_com_w_inst_n495,
         round_inst_S_7__sbox_inst_com_w_inst_n494,
         round_inst_S_7__sbox_inst_com_w_inst_n493,
         round_inst_S_7__sbox_inst_com_w_inst_n492,
         round_inst_S_7__sbox_inst_com_w_inst_n491,
         round_inst_S_7__sbox_inst_com_w_inst_n490,
         round_inst_S_7__sbox_inst_com_w_inst_n489,
         round_inst_S_7__sbox_inst_com_w_inst_n488,
         round_inst_S_7__sbox_inst_com_w_inst_n487,
         round_inst_S_7__sbox_inst_com_w_inst_n486,
         round_inst_S_7__sbox_inst_com_w_inst_n485,
         round_inst_S_7__sbox_inst_com_w_inst_n484,
         round_inst_S_7__sbox_inst_com_w_inst_n483,
         round_inst_S_7__sbox_inst_com_w_inst_n482,
         round_inst_S_7__sbox_inst_com_w_inst_n481,
         round_inst_S_7__sbox_inst_com_w_inst_n480,
         round_inst_S_7__sbox_inst_com_w_inst_n479,
         round_inst_S_7__sbox_inst_com_w_inst_n478,
         round_inst_S_7__sbox_inst_com_w_inst_n477,
         round_inst_S_7__sbox_inst_com_w_inst_n476,
         round_inst_S_7__sbox_inst_com_w_inst_n475,
         round_inst_S_7__sbox_inst_com_w_inst_n474,
         round_inst_S_7__sbox_inst_com_w_inst_n473,
         round_inst_S_7__sbox_inst_com_w_inst_n472,
         round_inst_S_7__sbox_inst_com_w_inst_n471,
         round_inst_S_7__sbox_inst_com_w_inst_n470,
         round_inst_S_7__sbox_inst_com_w_inst_n469,
         round_inst_S_7__sbox_inst_com_w_inst_n468,
         round_inst_S_7__sbox_inst_com_w_inst_n467,
         round_inst_S_7__sbox_inst_com_w_inst_n466,
         round_inst_S_7__sbox_inst_com_w_inst_n465,
         round_inst_S_7__sbox_inst_com_w_inst_n464,
         round_inst_S_7__sbox_inst_com_w_inst_n463,
         round_inst_S_7__sbox_inst_com_w_inst_n462,
         round_inst_S_7__sbox_inst_com_w_inst_n461,
         round_inst_S_7__sbox_inst_com_w_inst_n460,
         round_inst_S_7__sbox_inst_com_w_inst_n459,
         round_inst_S_7__sbox_inst_com_w_inst_n458,
         round_inst_S_7__sbox_inst_com_w_inst_n457,
         round_inst_S_7__sbox_inst_com_w_inst_n456,
         round_inst_S_7__sbox_inst_com_w_inst_n455,
         round_inst_S_7__sbox_inst_com_w_inst_n454,
         round_inst_S_7__sbox_inst_com_w_inst_n453,
         round_inst_S_7__sbox_inst_com_w_inst_n452,
         round_inst_S_7__sbox_inst_com_w_inst_n451,
         round_inst_S_7__sbox_inst_com_w_inst_n450,
         round_inst_S_7__sbox_inst_com_w_inst_n449,
         round_inst_S_7__sbox_inst_com_w_inst_n448,
         round_inst_S_7__sbox_inst_com_w_inst_n447,
         round_inst_S_7__sbox_inst_com_w_inst_n446,
         round_inst_S_7__sbox_inst_com_w_inst_n445,
         round_inst_S_7__sbox_inst_com_w_inst_n444,
         round_inst_S_7__sbox_inst_com_w_inst_n443,
         round_inst_S_7__sbox_inst_com_w_inst_n442,
         round_inst_S_7__sbox_inst_com_w_inst_n441,
         round_inst_S_7__sbox_inst_com_w_inst_n440,
         round_inst_S_7__sbox_inst_com_w_inst_n439,
         round_inst_S_7__sbox_inst_com_w_inst_n438,
         round_inst_S_7__sbox_inst_com_w_inst_n437,
         round_inst_S_7__sbox_inst_com_w_inst_n436,
         round_inst_S_7__sbox_inst_com_w_inst_n435,
         round_inst_S_7__sbox_inst_com_w_inst_n434,
         round_inst_S_7__sbox_inst_com_w_inst_n433,
         round_inst_S_7__sbox_inst_com_w_inst_n432,
         round_inst_S_7__sbox_inst_com_w_inst_n431,
         round_inst_S_7__sbox_inst_com_w_inst_n430,
         round_inst_S_7__sbox_inst_com_w_inst_n429,
         round_inst_S_7__sbox_inst_com_w_inst_n428,
         round_inst_S_7__sbox_inst_com_w_inst_n427,
         round_inst_S_7__sbox_inst_com_w_inst_n426,
         round_inst_S_7__sbox_inst_com_w_inst_n425,
         round_inst_S_7__sbox_inst_com_w_inst_n424,
         round_inst_S_7__sbox_inst_com_w_inst_n423,
         round_inst_S_7__sbox_inst_com_w_inst_n422,
         round_inst_S_7__sbox_inst_com_w_inst_n421,
         round_inst_S_7__sbox_inst_com_w_inst_n420,
         round_inst_S_7__sbox_inst_com_w_inst_n419,
         round_inst_S_7__sbox_inst_com_w_inst_n418,
         round_inst_S_7__sbox_inst_com_w_inst_n417,
         round_inst_S_7__sbox_inst_com_w_inst_n416,
         round_inst_S_7__sbox_inst_com_w_inst_n415,
         round_inst_S_7__sbox_inst_com_w_inst_n414,
         round_inst_S_7__sbox_inst_com_w_inst_n413,
         round_inst_S_7__sbox_inst_com_w_inst_n412,
         round_inst_S_7__sbox_inst_com_w_inst_n411,
         round_inst_S_7__sbox_inst_com_w_inst_n410,
         round_inst_S_7__sbox_inst_com_w_inst_n409,
         round_inst_S_7__sbox_inst_com_w_inst_n408,
         round_inst_S_7__sbox_inst_com_w_inst_n407,
         round_inst_S_7__sbox_inst_com_w_inst_n406,
         round_inst_S_7__sbox_inst_com_w_inst_n405,
         round_inst_S_7__sbox_inst_com_w_inst_n404,
         round_inst_S_7__sbox_inst_com_w_inst_n403,
         round_inst_S_7__sbox_inst_com_w_inst_n402,
         round_inst_S_7__sbox_inst_com_w_inst_n401,
         round_inst_S_7__sbox_inst_com_w_inst_n400,
         round_inst_S_7__sbox_inst_com_w_inst_n399,
         round_inst_S_7__sbox_inst_com_w_inst_n398,
         round_inst_S_7__sbox_inst_com_w_inst_n397,
         round_inst_S_7__sbox_inst_com_w_inst_n396,
         round_inst_S_7__sbox_inst_com_x_inst_n511,
         round_inst_S_7__sbox_inst_com_x_inst_n510,
         round_inst_S_7__sbox_inst_com_x_inst_n509,
         round_inst_S_7__sbox_inst_com_x_inst_n508,
         round_inst_S_7__sbox_inst_com_x_inst_n507,
         round_inst_S_7__sbox_inst_com_x_inst_n506,
         round_inst_S_7__sbox_inst_com_x_inst_n505,
         round_inst_S_7__sbox_inst_com_x_inst_n504,
         round_inst_S_7__sbox_inst_com_x_inst_n503,
         round_inst_S_7__sbox_inst_com_x_inst_n502,
         round_inst_S_7__sbox_inst_com_x_inst_n501,
         round_inst_S_7__sbox_inst_com_x_inst_n500,
         round_inst_S_7__sbox_inst_com_x_inst_n499,
         round_inst_S_7__sbox_inst_com_x_inst_n498,
         round_inst_S_7__sbox_inst_com_x_inst_n497,
         round_inst_S_7__sbox_inst_com_x_inst_n496,
         round_inst_S_7__sbox_inst_com_x_inst_n495,
         round_inst_S_7__sbox_inst_com_x_inst_n494,
         round_inst_S_7__sbox_inst_com_x_inst_n493,
         round_inst_S_7__sbox_inst_com_x_inst_n492,
         round_inst_S_7__sbox_inst_com_x_inst_n491,
         round_inst_S_7__sbox_inst_com_x_inst_n490,
         round_inst_S_7__sbox_inst_com_x_inst_n489,
         round_inst_S_7__sbox_inst_com_x_inst_n488,
         round_inst_S_7__sbox_inst_com_x_inst_n487,
         round_inst_S_7__sbox_inst_com_x_inst_n486,
         round_inst_S_7__sbox_inst_com_x_inst_n485,
         round_inst_S_7__sbox_inst_com_x_inst_n484,
         round_inst_S_7__sbox_inst_com_x_inst_n483,
         round_inst_S_7__sbox_inst_com_x_inst_n482,
         round_inst_S_7__sbox_inst_com_x_inst_n481,
         round_inst_S_7__sbox_inst_com_x_inst_n480,
         round_inst_S_7__sbox_inst_com_x_inst_n479,
         round_inst_S_7__sbox_inst_com_x_inst_n478,
         round_inst_S_7__sbox_inst_com_x_inst_n477,
         round_inst_S_7__sbox_inst_com_x_inst_n476,
         round_inst_S_7__sbox_inst_com_x_inst_n475,
         round_inst_S_7__sbox_inst_com_x_inst_n474,
         round_inst_S_7__sbox_inst_com_x_inst_n473,
         round_inst_S_7__sbox_inst_com_x_inst_n472,
         round_inst_S_7__sbox_inst_com_x_inst_n471,
         round_inst_S_7__sbox_inst_com_x_inst_n470,
         round_inst_S_7__sbox_inst_com_x_inst_n469,
         round_inst_S_7__sbox_inst_com_x_inst_n468,
         round_inst_S_7__sbox_inst_com_x_inst_n467,
         round_inst_S_7__sbox_inst_com_x_inst_n466,
         round_inst_S_7__sbox_inst_com_x_inst_n465,
         round_inst_S_7__sbox_inst_com_x_inst_n464,
         round_inst_S_7__sbox_inst_com_x_inst_n463,
         round_inst_S_7__sbox_inst_com_x_inst_n462,
         round_inst_S_7__sbox_inst_com_x_inst_n461,
         round_inst_S_7__sbox_inst_com_x_inst_n460,
         round_inst_S_7__sbox_inst_com_x_inst_n459,
         round_inst_S_7__sbox_inst_com_x_inst_n458,
         round_inst_S_7__sbox_inst_com_x_inst_n457,
         round_inst_S_7__sbox_inst_com_x_inst_n456,
         round_inst_S_7__sbox_inst_com_x_inst_n455,
         round_inst_S_7__sbox_inst_com_x_inst_n454,
         round_inst_S_7__sbox_inst_com_x_inst_n453,
         round_inst_S_7__sbox_inst_com_x_inst_n452,
         round_inst_S_7__sbox_inst_com_x_inst_n451,
         round_inst_S_7__sbox_inst_com_x_inst_n450,
         round_inst_S_7__sbox_inst_com_x_inst_n449,
         round_inst_S_7__sbox_inst_com_x_inst_n448,
         round_inst_S_7__sbox_inst_com_x_inst_n447,
         round_inst_S_7__sbox_inst_com_x_inst_n446,
         round_inst_S_7__sbox_inst_com_x_inst_n445,
         round_inst_S_7__sbox_inst_com_x_inst_n444,
         round_inst_S_7__sbox_inst_com_x_inst_n443,
         round_inst_S_7__sbox_inst_com_x_inst_n442,
         round_inst_S_7__sbox_inst_com_x_inst_n441,
         round_inst_S_7__sbox_inst_com_x_inst_n440,
         round_inst_S_7__sbox_inst_com_x_inst_n439,
         round_inst_S_7__sbox_inst_com_x_inst_n438,
         round_inst_S_7__sbox_inst_com_x_inst_n437,
         round_inst_S_7__sbox_inst_com_x_inst_n436,
         round_inst_S_7__sbox_inst_com_x_inst_n435,
         round_inst_S_7__sbox_inst_com_x_inst_n434,
         round_inst_S_7__sbox_inst_com_x_inst_n433,
         round_inst_S_7__sbox_inst_com_x_inst_n432,
         round_inst_S_7__sbox_inst_com_x_inst_n431,
         round_inst_S_7__sbox_inst_com_x_inst_n430,
         round_inst_S_7__sbox_inst_com_x_inst_n429,
         round_inst_S_7__sbox_inst_com_x_inst_n428,
         round_inst_S_7__sbox_inst_com_x_inst_n427,
         round_inst_S_7__sbox_inst_com_x_inst_n426,
         round_inst_S_7__sbox_inst_com_x_inst_n425,
         round_inst_S_7__sbox_inst_com_x_inst_n424,
         round_inst_S_7__sbox_inst_com_x_inst_n423,
         round_inst_S_7__sbox_inst_com_x_inst_n422,
         round_inst_S_7__sbox_inst_com_x_inst_n421,
         round_inst_S_7__sbox_inst_com_x_inst_n420,
         round_inst_S_7__sbox_inst_com_x_inst_n419,
         round_inst_S_7__sbox_inst_com_x_inst_n418,
         round_inst_S_7__sbox_inst_com_x_inst_n417,
         round_inst_S_7__sbox_inst_com_x_inst_n416,
         round_inst_S_7__sbox_inst_com_x_inst_n415,
         round_inst_S_7__sbox_inst_com_x_inst_n414,
         round_inst_S_7__sbox_inst_com_x_inst_n413,
         round_inst_S_7__sbox_inst_com_x_inst_n412,
         round_inst_S_7__sbox_inst_com_x_inst_n411,
         round_inst_S_7__sbox_inst_com_x_inst_n410,
         round_inst_S_7__sbox_inst_com_x_inst_n409,
         round_inst_S_7__sbox_inst_com_x_inst_n408,
         round_inst_S_7__sbox_inst_com_x_inst_n407,
         round_inst_S_7__sbox_inst_com_x_inst_n406,
         round_inst_S_7__sbox_inst_com_x_inst_n405,
         round_inst_S_7__sbox_inst_com_x_inst_n404,
         round_inst_S_7__sbox_inst_com_x_inst_n403,
         round_inst_S_7__sbox_inst_com_x_inst_n402,
         round_inst_S_7__sbox_inst_com_x_inst_n401,
         round_inst_S_7__sbox_inst_com_x_inst_n400,
         round_inst_S_7__sbox_inst_com_x_inst_n399,
         round_inst_S_7__sbox_inst_com_x_inst_n398,
         round_inst_S_7__sbox_inst_com_x_inst_n397,
         round_inst_S_7__sbox_inst_com_x_inst_n396,
         round_inst_S_7__sbox_inst_com_x_inst_n395,
         round_inst_S_7__sbox_inst_com_x_inst_n394,
         round_inst_S_7__sbox_inst_com_x_inst_n393,
         round_inst_S_7__sbox_inst_com_x_inst_n392,
         round_inst_S_7__sbox_inst_com_x_inst_n391,
         round_inst_S_7__sbox_inst_com_x_inst_n390,
         round_inst_S_7__sbox_inst_com_x_inst_n389,
         round_inst_S_7__sbox_inst_com_x_inst_n388,
         round_inst_S_7__sbox_inst_com_x_inst_n387,
         round_inst_S_7__sbox_inst_com_x_inst_n386,
         round_inst_S_7__sbox_inst_com_x_inst_n385,
         round_inst_S_7__sbox_inst_com_x_inst_n384,
         round_inst_S_7__sbox_inst_com_x_inst_n383,
         round_inst_S_7__sbox_inst_com_x_inst_n382,
         round_inst_S_7__sbox_inst_com_x_inst_n381,
         round_inst_S_7__sbox_inst_com_y_inst_n518,
         round_inst_S_7__sbox_inst_com_y_inst_n517,
         round_inst_S_7__sbox_inst_com_y_inst_n516,
         round_inst_S_7__sbox_inst_com_y_inst_n515,
         round_inst_S_7__sbox_inst_com_y_inst_n514,
         round_inst_S_7__sbox_inst_com_y_inst_n513,
         round_inst_S_7__sbox_inst_com_y_inst_n512,
         round_inst_S_7__sbox_inst_com_y_inst_n511,
         round_inst_S_7__sbox_inst_com_y_inst_n510,
         round_inst_S_7__sbox_inst_com_y_inst_n509,
         round_inst_S_7__sbox_inst_com_y_inst_n508,
         round_inst_S_7__sbox_inst_com_y_inst_n507,
         round_inst_S_7__sbox_inst_com_y_inst_n506,
         round_inst_S_7__sbox_inst_com_y_inst_n505,
         round_inst_S_7__sbox_inst_com_y_inst_n504,
         round_inst_S_7__sbox_inst_com_y_inst_n503,
         round_inst_S_7__sbox_inst_com_y_inst_n502,
         round_inst_S_7__sbox_inst_com_y_inst_n501,
         round_inst_S_7__sbox_inst_com_y_inst_n500,
         round_inst_S_7__sbox_inst_com_y_inst_n499,
         round_inst_S_7__sbox_inst_com_y_inst_n498,
         round_inst_S_7__sbox_inst_com_y_inst_n497,
         round_inst_S_7__sbox_inst_com_y_inst_n496,
         round_inst_S_7__sbox_inst_com_y_inst_n495,
         round_inst_S_7__sbox_inst_com_y_inst_n494,
         round_inst_S_7__sbox_inst_com_y_inst_n493,
         round_inst_S_7__sbox_inst_com_y_inst_n492,
         round_inst_S_7__sbox_inst_com_y_inst_n491,
         round_inst_S_7__sbox_inst_com_y_inst_n490,
         round_inst_S_7__sbox_inst_com_y_inst_n489,
         round_inst_S_7__sbox_inst_com_y_inst_n488,
         round_inst_S_7__sbox_inst_com_y_inst_n487,
         round_inst_S_7__sbox_inst_com_y_inst_n486,
         round_inst_S_7__sbox_inst_com_y_inst_n485,
         round_inst_S_7__sbox_inst_com_y_inst_n484,
         round_inst_S_7__sbox_inst_com_y_inst_n483,
         round_inst_S_7__sbox_inst_com_y_inst_n482,
         round_inst_S_7__sbox_inst_com_y_inst_n481,
         round_inst_S_7__sbox_inst_com_y_inst_n480,
         round_inst_S_7__sbox_inst_com_y_inst_n479,
         round_inst_S_7__sbox_inst_com_y_inst_n478,
         round_inst_S_7__sbox_inst_com_y_inst_n477,
         round_inst_S_7__sbox_inst_com_y_inst_n476,
         round_inst_S_7__sbox_inst_com_y_inst_n475,
         round_inst_S_7__sbox_inst_com_y_inst_n474,
         round_inst_S_7__sbox_inst_com_y_inst_n473,
         round_inst_S_7__sbox_inst_com_y_inst_n472,
         round_inst_S_7__sbox_inst_com_y_inst_n471,
         round_inst_S_7__sbox_inst_com_y_inst_n470,
         round_inst_S_7__sbox_inst_com_y_inst_n469,
         round_inst_S_7__sbox_inst_com_y_inst_n468,
         round_inst_S_7__sbox_inst_com_y_inst_n467,
         round_inst_S_7__sbox_inst_com_y_inst_n466,
         round_inst_S_7__sbox_inst_com_y_inst_n465,
         round_inst_S_7__sbox_inst_com_y_inst_n464,
         round_inst_S_7__sbox_inst_com_y_inst_n463,
         round_inst_S_7__sbox_inst_com_y_inst_n462,
         round_inst_S_7__sbox_inst_com_y_inst_n461,
         round_inst_S_7__sbox_inst_com_y_inst_n460,
         round_inst_S_7__sbox_inst_com_y_inst_n459,
         round_inst_S_7__sbox_inst_com_y_inst_n458,
         round_inst_S_7__sbox_inst_com_y_inst_n457,
         round_inst_S_7__sbox_inst_com_y_inst_n456,
         round_inst_S_7__sbox_inst_com_y_inst_n455,
         round_inst_S_7__sbox_inst_com_y_inst_n454,
         round_inst_S_7__sbox_inst_com_y_inst_n453,
         round_inst_S_7__sbox_inst_com_y_inst_n452,
         round_inst_S_7__sbox_inst_com_y_inst_n451,
         round_inst_S_7__sbox_inst_com_y_inst_n450,
         round_inst_S_7__sbox_inst_com_y_inst_n449,
         round_inst_S_7__sbox_inst_com_y_inst_n448,
         round_inst_S_7__sbox_inst_com_y_inst_n447,
         round_inst_S_7__sbox_inst_com_y_inst_n446,
         round_inst_S_7__sbox_inst_com_y_inst_n445,
         round_inst_S_7__sbox_inst_com_y_inst_n444,
         round_inst_S_7__sbox_inst_com_y_inst_n443,
         round_inst_S_7__sbox_inst_com_y_inst_n442,
         round_inst_S_7__sbox_inst_com_y_inst_n441,
         round_inst_S_7__sbox_inst_com_y_inst_n440,
         round_inst_S_7__sbox_inst_com_y_inst_n439,
         round_inst_S_7__sbox_inst_com_y_inst_n438,
         round_inst_S_7__sbox_inst_com_y_inst_n437,
         round_inst_S_7__sbox_inst_com_y_inst_n436,
         round_inst_S_7__sbox_inst_com_y_inst_n435,
         round_inst_S_7__sbox_inst_com_y_inst_n434,
         round_inst_S_7__sbox_inst_com_y_inst_n433,
         round_inst_S_7__sbox_inst_com_y_inst_n432,
         round_inst_S_7__sbox_inst_com_y_inst_n431,
         round_inst_S_7__sbox_inst_com_y_inst_n430,
         round_inst_S_7__sbox_inst_com_y_inst_n429,
         round_inst_S_7__sbox_inst_com_y_inst_n428,
         round_inst_S_7__sbox_inst_com_y_inst_n427,
         round_inst_S_7__sbox_inst_com_y_inst_n426,
         round_inst_S_7__sbox_inst_com_y_inst_n425,
         round_inst_S_7__sbox_inst_com_y_inst_n424,
         round_inst_S_7__sbox_inst_com_y_inst_n423,
         round_inst_S_7__sbox_inst_com_y_inst_n422,
         round_inst_S_7__sbox_inst_com_y_inst_n421,
         round_inst_S_7__sbox_inst_com_y_inst_n420,
         round_inst_S_7__sbox_inst_com_y_inst_n419,
         round_inst_S_7__sbox_inst_com_y_inst_n418,
         round_inst_S_7__sbox_inst_com_y_inst_n417,
         round_inst_S_7__sbox_inst_com_y_inst_n416,
         round_inst_S_7__sbox_inst_com_y_inst_n415,
         round_inst_S_7__sbox_inst_com_y_inst_n414,
         round_inst_S_7__sbox_inst_com_y_inst_n413,
         round_inst_S_7__sbox_inst_com_y_inst_n412,
         round_inst_S_7__sbox_inst_com_y_inst_n411,
         round_inst_S_7__sbox_inst_com_y_inst_n410,
         round_inst_S_7__sbox_inst_com_y_inst_n409,
         round_inst_S_7__sbox_inst_com_y_inst_n408,
         round_inst_S_7__sbox_inst_com_y_inst_n407,
         round_inst_S_7__sbox_inst_com_y_inst_n406,
         round_inst_S_7__sbox_inst_com_y_inst_n405,
         round_inst_S_7__sbox_inst_com_y_inst_n404,
         round_inst_S_7__sbox_inst_com_y_inst_n403,
         round_inst_S_7__sbox_inst_com_y_inst_n402,
         round_inst_S_7__sbox_inst_com_y_inst_n401,
         round_inst_S_7__sbox_inst_com_y_inst_n400,
         round_inst_S_7__sbox_inst_com_y_inst_n399,
         round_inst_S_7__sbox_inst_com_y_inst_n398,
         round_inst_S_7__sbox_inst_com_y_inst_n397,
         round_inst_S_7__sbox_inst_com_y_inst_n396,
         round_inst_S_7__sbox_inst_com_y_inst_n395,
         round_inst_S_7__sbox_inst_com_y_inst_n394,
         round_inst_S_7__sbox_inst_com_y_inst_n393,
         round_inst_S_7__sbox_inst_com_y_inst_n392,
         round_inst_S_7__sbox_inst_com_y_inst_n391,
         round_inst_S_7__sbox_inst_com_y_inst_n390,
         round_inst_S_7__sbox_inst_com_y_inst_n389,
         round_inst_S_7__sbox_inst_com_y_inst_n388,
         round_inst_S_7__sbox_inst_com_y_inst_n387,
         round_inst_S_7__sbox_inst_com_y_inst_n386,
         round_inst_S_7__sbox_inst_com_z_inst_n516,
         round_inst_S_7__sbox_inst_com_z_inst_n515,
         round_inst_S_7__sbox_inst_com_z_inst_n514,
         round_inst_S_7__sbox_inst_com_z_inst_n513,
         round_inst_S_7__sbox_inst_com_z_inst_n512,
         round_inst_S_7__sbox_inst_com_z_inst_n511,
         round_inst_S_7__sbox_inst_com_z_inst_n510,
         round_inst_S_7__sbox_inst_com_z_inst_n509,
         round_inst_S_7__sbox_inst_com_z_inst_n508,
         round_inst_S_7__sbox_inst_com_z_inst_n507,
         round_inst_S_7__sbox_inst_com_z_inst_n506,
         round_inst_S_7__sbox_inst_com_z_inst_n505,
         round_inst_S_7__sbox_inst_com_z_inst_n504,
         round_inst_S_7__sbox_inst_com_z_inst_n503,
         round_inst_S_7__sbox_inst_com_z_inst_n502,
         round_inst_S_7__sbox_inst_com_z_inst_n501,
         round_inst_S_7__sbox_inst_com_z_inst_n500,
         round_inst_S_7__sbox_inst_com_z_inst_n499,
         round_inst_S_7__sbox_inst_com_z_inst_n498,
         round_inst_S_7__sbox_inst_com_z_inst_n497,
         round_inst_S_7__sbox_inst_com_z_inst_n496,
         round_inst_S_7__sbox_inst_com_z_inst_n495,
         round_inst_S_7__sbox_inst_com_z_inst_n494,
         round_inst_S_7__sbox_inst_com_z_inst_n493,
         round_inst_S_7__sbox_inst_com_z_inst_n492,
         round_inst_S_7__sbox_inst_com_z_inst_n491,
         round_inst_S_7__sbox_inst_com_z_inst_n490,
         round_inst_S_7__sbox_inst_com_z_inst_n489,
         round_inst_S_7__sbox_inst_com_z_inst_n488,
         round_inst_S_7__sbox_inst_com_z_inst_n487,
         round_inst_S_7__sbox_inst_com_z_inst_n486,
         round_inst_S_7__sbox_inst_com_z_inst_n485,
         round_inst_S_7__sbox_inst_com_z_inst_n484,
         round_inst_S_7__sbox_inst_com_z_inst_n483,
         round_inst_S_7__sbox_inst_com_z_inst_n482,
         round_inst_S_7__sbox_inst_com_z_inst_n481,
         round_inst_S_7__sbox_inst_com_z_inst_n480,
         round_inst_S_7__sbox_inst_com_z_inst_n479,
         round_inst_S_7__sbox_inst_com_z_inst_n478,
         round_inst_S_7__sbox_inst_com_z_inst_n477,
         round_inst_S_7__sbox_inst_com_z_inst_n476,
         round_inst_S_7__sbox_inst_com_z_inst_n475,
         round_inst_S_7__sbox_inst_com_z_inst_n474,
         round_inst_S_7__sbox_inst_com_z_inst_n473,
         round_inst_S_7__sbox_inst_com_z_inst_n472,
         round_inst_S_7__sbox_inst_com_z_inst_n471,
         round_inst_S_7__sbox_inst_com_z_inst_n470,
         round_inst_S_7__sbox_inst_com_z_inst_n469,
         round_inst_S_7__sbox_inst_com_z_inst_n468,
         round_inst_S_7__sbox_inst_com_z_inst_n467,
         round_inst_S_7__sbox_inst_com_z_inst_n466,
         round_inst_S_7__sbox_inst_com_z_inst_n465,
         round_inst_S_7__sbox_inst_com_z_inst_n464,
         round_inst_S_7__sbox_inst_com_z_inst_n463,
         round_inst_S_7__sbox_inst_com_z_inst_n462,
         round_inst_S_7__sbox_inst_com_z_inst_n461,
         round_inst_S_7__sbox_inst_com_z_inst_n460,
         round_inst_S_7__sbox_inst_com_z_inst_n459,
         round_inst_S_7__sbox_inst_com_z_inst_n458,
         round_inst_S_7__sbox_inst_com_z_inst_n457,
         round_inst_S_7__sbox_inst_com_z_inst_n456,
         round_inst_S_7__sbox_inst_com_z_inst_n455,
         round_inst_S_7__sbox_inst_com_z_inst_n454,
         round_inst_S_7__sbox_inst_com_z_inst_n453,
         round_inst_S_7__sbox_inst_com_z_inst_n452,
         round_inst_S_7__sbox_inst_com_z_inst_n451,
         round_inst_S_7__sbox_inst_com_z_inst_n450,
         round_inst_S_7__sbox_inst_com_z_inst_n449,
         round_inst_S_7__sbox_inst_com_z_inst_n448,
         round_inst_S_7__sbox_inst_com_z_inst_n447,
         round_inst_S_7__sbox_inst_com_z_inst_n446,
         round_inst_S_7__sbox_inst_com_z_inst_n445,
         round_inst_S_7__sbox_inst_com_z_inst_n444,
         round_inst_S_7__sbox_inst_com_z_inst_n443,
         round_inst_S_7__sbox_inst_com_z_inst_n442,
         round_inst_S_7__sbox_inst_com_z_inst_n441,
         round_inst_S_7__sbox_inst_com_z_inst_n440,
         round_inst_S_7__sbox_inst_com_z_inst_n439,
         round_inst_S_7__sbox_inst_com_z_inst_n438,
         round_inst_S_7__sbox_inst_com_z_inst_n437,
         round_inst_S_7__sbox_inst_com_z_inst_n436,
         round_inst_S_7__sbox_inst_com_z_inst_n435,
         round_inst_S_7__sbox_inst_com_z_inst_n434,
         round_inst_S_7__sbox_inst_com_z_inst_n433,
         round_inst_S_7__sbox_inst_com_z_inst_n432,
         round_inst_S_7__sbox_inst_com_z_inst_n431,
         round_inst_S_7__sbox_inst_com_z_inst_n430,
         round_inst_S_7__sbox_inst_com_z_inst_n429,
         round_inst_S_7__sbox_inst_com_z_inst_n428,
         round_inst_S_7__sbox_inst_com_z_inst_n427,
         round_inst_S_7__sbox_inst_com_z_inst_n426,
         round_inst_S_7__sbox_inst_com_z_inst_n425,
         round_inst_S_7__sbox_inst_com_z_inst_n424,
         round_inst_S_7__sbox_inst_com_z_inst_n423,
         round_inst_S_7__sbox_inst_com_z_inst_n422,
         round_inst_S_7__sbox_inst_com_z_inst_n421,
         round_inst_S_7__sbox_inst_com_z_inst_n420,
         round_inst_S_7__sbox_inst_com_z_inst_n419,
         round_inst_S_7__sbox_inst_com_z_inst_n418,
         round_inst_S_7__sbox_inst_com_z_inst_n417,
         round_inst_S_7__sbox_inst_com_z_inst_n416,
         round_inst_S_7__sbox_inst_com_z_inst_n415,
         round_inst_S_7__sbox_inst_com_z_inst_n414,
         round_inst_S_7__sbox_inst_com_z_inst_n413,
         round_inst_S_7__sbox_inst_com_z_inst_n412,
         round_inst_S_7__sbox_inst_com_z_inst_n411,
         round_inst_S_7__sbox_inst_com_z_inst_n410,
         round_inst_S_7__sbox_inst_com_z_inst_n409,
         round_inst_S_7__sbox_inst_com_z_inst_n408,
         round_inst_S_7__sbox_inst_com_z_inst_n407,
         round_inst_S_7__sbox_inst_com_z_inst_n406,
         round_inst_S_7__sbox_inst_com_z_inst_n405,
         round_inst_S_7__sbox_inst_com_z_inst_n404,
         round_inst_S_7__sbox_inst_com_z_inst_n403,
         round_inst_S_7__sbox_inst_com_z_inst_n402,
         round_inst_S_7__sbox_inst_com_z_inst_n401,
         round_inst_S_7__sbox_inst_com_z_inst_n400,
         round_inst_S_7__sbox_inst_com_z_inst_n399,
         round_inst_S_7__sbox_inst_com_z_inst_n398,
         round_inst_S_7__sbox_inst_com_z_inst_n397,
         round_inst_S_7__sbox_inst_com_z_inst_n396,
         round_inst_S_7__sbox_inst_com_z_inst_n395,
         round_inst_S_7__sbox_inst_com_z_inst_n394,
         round_inst_S_7__sbox_inst_com_z_inst_n393,
         round_inst_S_7__sbox_inst_com_z_inst_n392,
         round_inst_S_7__sbox_inst_com_z_inst_n391,
         round_inst_S_7__sbox_inst_com_z_inst_n390,
         round_inst_S_8__sbox_inst_n6, round_inst_S_8__sbox_inst_n5,
         round_inst_S_8__sbox_inst_n4, round_inst_S_8__sbox_inst_n3,
         round_inst_S_8__sbox_inst_n2, round_inst_S_8__sbox_inst_n1,
         round_inst_S_8__sbox_inst_com_w_inst_n529,
         round_inst_S_8__sbox_inst_com_w_inst_n528,
         round_inst_S_8__sbox_inst_com_w_inst_n527,
         round_inst_S_8__sbox_inst_com_w_inst_n526,
         round_inst_S_8__sbox_inst_com_w_inst_n525,
         round_inst_S_8__sbox_inst_com_w_inst_n524,
         round_inst_S_8__sbox_inst_com_w_inst_n523,
         round_inst_S_8__sbox_inst_com_w_inst_n522,
         round_inst_S_8__sbox_inst_com_w_inst_n521,
         round_inst_S_8__sbox_inst_com_w_inst_n520,
         round_inst_S_8__sbox_inst_com_w_inst_n519,
         round_inst_S_8__sbox_inst_com_w_inst_n518,
         round_inst_S_8__sbox_inst_com_w_inst_n517,
         round_inst_S_8__sbox_inst_com_w_inst_n516,
         round_inst_S_8__sbox_inst_com_w_inst_n515,
         round_inst_S_8__sbox_inst_com_w_inst_n514,
         round_inst_S_8__sbox_inst_com_w_inst_n513,
         round_inst_S_8__sbox_inst_com_w_inst_n512,
         round_inst_S_8__sbox_inst_com_w_inst_n511,
         round_inst_S_8__sbox_inst_com_w_inst_n510,
         round_inst_S_8__sbox_inst_com_w_inst_n509,
         round_inst_S_8__sbox_inst_com_w_inst_n508,
         round_inst_S_8__sbox_inst_com_w_inst_n507,
         round_inst_S_8__sbox_inst_com_w_inst_n506,
         round_inst_S_8__sbox_inst_com_w_inst_n505,
         round_inst_S_8__sbox_inst_com_w_inst_n504,
         round_inst_S_8__sbox_inst_com_w_inst_n503,
         round_inst_S_8__sbox_inst_com_w_inst_n502,
         round_inst_S_8__sbox_inst_com_w_inst_n501,
         round_inst_S_8__sbox_inst_com_w_inst_n500,
         round_inst_S_8__sbox_inst_com_w_inst_n499,
         round_inst_S_8__sbox_inst_com_w_inst_n498,
         round_inst_S_8__sbox_inst_com_w_inst_n497,
         round_inst_S_8__sbox_inst_com_w_inst_n496,
         round_inst_S_8__sbox_inst_com_w_inst_n495,
         round_inst_S_8__sbox_inst_com_w_inst_n494,
         round_inst_S_8__sbox_inst_com_w_inst_n493,
         round_inst_S_8__sbox_inst_com_w_inst_n492,
         round_inst_S_8__sbox_inst_com_w_inst_n491,
         round_inst_S_8__sbox_inst_com_w_inst_n490,
         round_inst_S_8__sbox_inst_com_w_inst_n489,
         round_inst_S_8__sbox_inst_com_w_inst_n488,
         round_inst_S_8__sbox_inst_com_w_inst_n487,
         round_inst_S_8__sbox_inst_com_w_inst_n486,
         round_inst_S_8__sbox_inst_com_w_inst_n485,
         round_inst_S_8__sbox_inst_com_w_inst_n484,
         round_inst_S_8__sbox_inst_com_w_inst_n483,
         round_inst_S_8__sbox_inst_com_w_inst_n482,
         round_inst_S_8__sbox_inst_com_w_inst_n481,
         round_inst_S_8__sbox_inst_com_w_inst_n480,
         round_inst_S_8__sbox_inst_com_w_inst_n479,
         round_inst_S_8__sbox_inst_com_w_inst_n478,
         round_inst_S_8__sbox_inst_com_w_inst_n477,
         round_inst_S_8__sbox_inst_com_w_inst_n476,
         round_inst_S_8__sbox_inst_com_w_inst_n475,
         round_inst_S_8__sbox_inst_com_w_inst_n474,
         round_inst_S_8__sbox_inst_com_w_inst_n473,
         round_inst_S_8__sbox_inst_com_w_inst_n472,
         round_inst_S_8__sbox_inst_com_w_inst_n471,
         round_inst_S_8__sbox_inst_com_w_inst_n470,
         round_inst_S_8__sbox_inst_com_w_inst_n469,
         round_inst_S_8__sbox_inst_com_w_inst_n468,
         round_inst_S_8__sbox_inst_com_w_inst_n467,
         round_inst_S_8__sbox_inst_com_w_inst_n466,
         round_inst_S_8__sbox_inst_com_w_inst_n465,
         round_inst_S_8__sbox_inst_com_w_inst_n464,
         round_inst_S_8__sbox_inst_com_w_inst_n463,
         round_inst_S_8__sbox_inst_com_w_inst_n462,
         round_inst_S_8__sbox_inst_com_w_inst_n461,
         round_inst_S_8__sbox_inst_com_w_inst_n460,
         round_inst_S_8__sbox_inst_com_w_inst_n459,
         round_inst_S_8__sbox_inst_com_w_inst_n458,
         round_inst_S_8__sbox_inst_com_w_inst_n457,
         round_inst_S_8__sbox_inst_com_w_inst_n456,
         round_inst_S_8__sbox_inst_com_w_inst_n455,
         round_inst_S_8__sbox_inst_com_w_inst_n454,
         round_inst_S_8__sbox_inst_com_w_inst_n453,
         round_inst_S_8__sbox_inst_com_w_inst_n452,
         round_inst_S_8__sbox_inst_com_w_inst_n451,
         round_inst_S_8__sbox_inst_com_w_inst_n450,
         round_inst_S_8__sbox_inst_com_w_inst_n449,
         round_inst_S_8__sbox_inst_com_w_inst_n448,
         round_inst_S_8__sbox_inst_com_w_inst_n447,
         round_inst_S_8__sbox_inst_com_w_inst_n446,
         round_inst_S_8__sbox_inst_com_w_inst_n445,
         round_inst_S_8__sbox_inst_com_w_inst_n444,
         round_inst_S_8__sbox_inst_com_w_inst_n443,
         round_inst_S_8__sbox_inst_com_w_inst_n442,
         round_inst_S_8__sbox_inst_com_w_inst_n441,
         round_inst_S_8__sbox_inst_com_w_inst_n440,
         round_inst_S_8__sbox_inst_com_w_inst_n439,
         round_inst_S_8__sbox_inst_com_w_inst_n438,
         round_inst_S_8__sbox_inst_com_w_inst_n437,
         round_inst_S_8__sbox_inst_com_w_inst_n436,
         round_inst_S_8__sbox_inst_com_w_inst_n435,
         round_inst_S_8__sbox_inst_com_w_inst_n434,
         round_inst_S_8__sbox_inst_com_w_inst_n433,
         round_inst_S_8__sbox_inst_com_w_inst_n432,
         round_inst_S_8__sbox_inst_com_w_inst_n431,
         round_inst_S_8__sbox_inst_com_w_inst_n430,
         round_inst_S_8__sbox_inst_com_w_inst_n429,
         round_inst_S_8__sbox_inst_com_w_inst_n428,
         round_inst_S_8__sbox_inst_com_w_inst_n427,
         round_inst_S_8__sbox_inst_com_w_inst_n426,
         round_inst_S_8__sbox_inst_com_w_inst_n425,
         round_inst_S_8__sbox_inst_com_w_inst_n424,
         round_inst_S_8__sbox_inst_com_w_inst_n423,
         round_inst_S_8__sbox_inst_com_w_inst_n422,
         round_inst_S_8__sbox_inst_com_w_inst_n421,
         round_inst_S_8__sbox_inst_com_w_inst_n420,
         round_inst_S_8__sbox_inst_com_w_inst_n419,
         round_inst_S_8__sbox_inst_com_w_inst_n418,
         round_inst_S_8__sbox_inst_com_w_inst_n417,
         round_inst_S_8__sbox_inst_com_w_inst_n416,
         round_inst_S_8__sbox_inst_com_w_inst_n415,
         round_inst_S_8__sbox_inst_com_w_inst_n414,
         round_inst_S_8__sbox_inst_com_w_inst_n413,
         round_inst_S_8__sbox_inst_com_w_inst_n412,
         round_inst_S_8__sbox_inst_com_w_inst_n411,
         round_inst_S_8__sbox_inst_com_w_inst_n410,
         round_inst_S_8__sbox_inst_com_w_inst_n409,
         round_inst_S_8__sbox_inst_com_w_inst_n408,
         round_inst_S_8__sbox_inst_com_w_inst_n407,
         round_inst_S_8__sbox_inst_com_w_inst_n406,
         round_inst_S_8__sbox_inst_com_w_inst_n405,
         round_inst_S_8__sbox_inst_com_w_inst_n404,
         round_inst_S_8__sbox_inst_com_w_inst_n403,
         round_inst_S_8__sbox_inst_com_w_inst_n402,
         round_inst_S_8__sbox_inst_com_w_inst_n401,
         round_inst_S_8__sbox_inst_com_w_inst_n400,
         round_inst_S_8__sbox_inst_com_w_inst_n399,
         round_inst_S_8__sbox_inst_com_w_inst_n398,
         round_inst_S_8__sbox_inst_com_w_inst_n397,
         round_inst_S_8__sbox_inst_com_w_inst_n396,
         round_inst_S_8__sbox_inst_com_x_inst_n512,
         round_inst_S_8__sbox_inst_com_x_inst_n511,
         round_inst_S_8__sbox_inst_com_x_inst_n510,
         round_inst_S_8__sbox_inst_com_x_inst_n509,
         round_inst_S_8__sbox_inst_com_x_inst_n508,
         round_inst_S_8__sbox_inst_com_x_inst_n507,
         round_inst_S_8__sbox_inst_com_x_inst_n506,
         round_inst_S_8__sbox_inst_com_x_inst_n505,
         round_inst_S_8__sbox_inst_com_x_inst_n504,
         round_inst_S_8__sbox_inst_com_x_inst_n503,
         round_inst_S_8__sbox_inst_com_x_inst_n502,
         round_inst_S_8__sbox_inst_com_x_inst_n501,
         round_inst_S_8__sbox_inst_com_x_inst_n500,
         round_inst_S_8__sbox_inst_com_x_inst_n499,
         round_inst_S_8__sbox_inst_com_x_inst_n498,
         round_inst_S_8__sbox_inst_com_x_inst_n497,
         round_inst_S_8__sbox_inst_com_x_inst_n496,
         round_inst_S_8__sbox_inst_com_x_inst_n495,
         round_inst_S_8__sbox_inst_com_x_inst_n494,
         round_inst_S_8__sbox_inst_com_x_inst_n493,
         round_inst_S_8__sbox_inst_com_x_inst_n492,
         round_inst_S_8__sbox_inst_com_x_inst_n491,
         round_inst_S_8__sbox_inst_com_x_inst_n490,
         round_inst_S_8__sbox_inst_com_x_inst_n489,
         round_inst_S_8__sbox_inst_com_x_inst_n488,
         round_inst_S_8__sbox_inst_com_x_inst_n487,
         round_inst_S_8__sbox_inst_com_x_inst_n486,
         round_inst_S_8__sbox_inst_com_x_inst_n485,
         round_inst_S_8__sbox_inst_com_x_inst_n484,
         round_inst_S_8__sbox_inst_com_x_inst_n483,
         round_inst_S_8__sbox_inst_com_x_inst_n482,
         round_inst_S_8__sbox_inst_com_x_inst_n481,
         round_inst_S_8__sbox_inst_com_x_inst_n480,
         round_inst_S_8__sbox_inst_com_x_inst_n479,
         round_inst_S_8__sbox_inst_com_x_inst_n478,
         round_inst_S_8__sbox_inst_com_x_inst_n477,
         round_inst_S_8__sbox_inst_com_x_inst_n476,
         round_inst_S_8__sbox_inst_com_x_inst_n475,
         round_inst_S_8__sbox_inst_com_x_inst_n474,
         round_inst_S_8__sbox_inst_com_x_inst_n473,
         round_inst_S_8__sbox_inst_com_x_inst_n472,
         round_inst_S_8__sbox_inst_com_x_inst_n471,
         round_inst_S_8__sbox_inst_com_x_inst_n470,
         round_inst_S_8__sbox_inst_com_x_inst_n469,
         round_inst_S_8__sbox_inst_com_x_inst_n468,
         round_inst_S_8__sbox_inst_com_x_inst_n467,
         round_inst_S_8__sbox_inst_com_x_inst_n466,
         round_inst_S_8__sbox_inst_com_x_inst_n465,
         round_inst_S_8__sbox_inst_com_x_inst_n464,
         round_inst_S_8__sbox_inst_com_x_inst_n463,
         round_inst_S_8__sbox_inst_com_x_inst_n462,
         round_inst_S_8__sbox_inst_com_x_inst_n461,
         round_inst_S_8__sbox_inst_com_x_inst_n460,
         round_inst_S_8__sbox_inst_com_x_inst_n459,
         round_inst_S_8__sbox_inst_com_x_inst_n458,
         round_inst_S_8__sbox_inst_com_x_inst_n457,
         round_inst_S_8__sbox_inst_com_x_inst_n456,
         round_inst_S_8__sbox_inst_com_x_inst_n455,
         round_inst_S_8__sbox_inst_com_x_inst_n454,
         round_inst_S_8__sbox_inst_com_x_inst_n453,
         round_inst_S_8__sbox_inst_com_x_inst_n452,
         round_inst_S_8__sbox_inst_com_x_inst_n451,
         round_inst_S_8__sbox_inst_com_x_inst_n450,
         round_inst_S_8__sbox_inst_com_x_inst_n449,
         round_inst_S_8__sbox_inst_com_x_inst_n448,
         round_inst_S_8__sbox_inst_com_x_inst_n447,
         round_inst_S_8__sbox_inst_com_x_inst_n446,
         round_inst_S_8__sbox_inst_com_x_inst_n445,
         round_inst_S_8__sbox_inst_com_x_inst_n444,
         round_inst_S_8__sbox_inst_com_x_inst_n443,
         round_inst_S_8__sbox_inst_com_x_inst_n442,
         round_inst_S_8__sbox_inst_com_x_inst_n441,
         round_inst_S_8__sbox_inst_com_x_inst_n440,
         round_inst_S_8__sbox_inst_com_x_inst_n439,
         round_inst_S_8__sbox_inst_com_x_inst_n438,
         round_inst_S_8__sbox_inst_com_x_inst_n437,
         round_inst_S_8__sbox_inst_com_x_inst_n436,
         round_inst_S_8__sbox_inst_com_x_inst_n435,
         round_inst_S_8__sbox_inst_com_x_inst_n434,
         round_inst_S_8__sbox_inst_com_x_inst_n433,
         round_inst_S_8__sbox_inst_com_x_inst_n432,
         round_inst_S_8__sbox_inst_com_x_inst_n431,
         round_inst_S_8__sbox_inst_com_x_inst_n430,
         round_inst_S_8__sbox_inst_com_x_inst_n429,
         round_inst_S_8__sbox_inst_com_x_inst_n428,
         round_inst_S_8__sbox_inst_com_x_inst_n427,
         round_inst_S_8__sbox_inst_com_x_inst_n426,
         round_inst_S_8__sbox_inst_com_x_inst_n425,
         round_inst_S_8__sbox_inst_com_x_inst_n424,
         round_inst_S_8__sbox_inst_com_x_inst_n423,
         round_inst_S_8__sbox_inst_com_x_inst_n422,
         round_inst_S_8__sbox_inst_com_x_inst_n421,
         round_inst_S_8__sbox_inst_com_x_inst_n420,
         round_inst_S_8__sbox_inst_com_x_inst_n419,
         round_inst_S_8__sbox_inst_com_x_inst_n418,
         round_inst_S_8__sbox_inst_com_x_inst_n417,
         round_inst_S_8__sbox_inst_com_x_inst_n416,
         round_inst_S_8__sbox_inst_com_x_inst_n415,
         round_inst_S_8__sbox_inst_com_x_inst_n414,
         round_inst_S_8__sbox_inst_com_x_inst_n413,
         round_inst_S_8__sbox_inst_com_x_inst_n412,
         round_inst_S_8__sbox_inst_com_x_inst_n411,
         round_inst_S_8__sbox_inst_com_x_inst_n410,
         round_inst_S_8__sbox_inst_com_x_inst_n409,
         round_inst_S_8__sbox_inst_com_x_inst_n408,
         round_inst_S_8__sbox_inst_com_x_inst_n407,
         round_inst_S_8__sbox_inst_com_x_inst_n406,
         round_inst_S_8__sbox_inst_com_x_inst_n405,
         round_inst_S_8__sbox_inst_com_x_inst_n404,
         round_inst_S_8__sbox_inst_com_x_inst_n403,
         round_inst_S_8__sbox_inst_com_x_inst_n402,
         round_inst_S_8__sbox_inst_com_x_inst_n401,
         round_inst_S_8__sbox_inst_com_x_inst_n400,
         round_inst_S_8__sbox_inst_com_x_inst_n399,
         round_inst_S_8__sbox_inst_com_x_inst_n398,
         round_inst_S_8__sbox_inst_com_x_inst_n397,
         round_inst_S_8__sbox_inst_com_x_inst_n396,
         round_inst_S_8__sbox_inst_com_x_inst_n395,
         round_inst_S_8__sbox_inst_com_x_inst_n394,
         round_inst_S_8__sbox_inst_com_x_inst_n393,
         round_inst_S_8__sbox_inst_com_x_inst_n392,
         round_inst_S_8__sbox_inst_com_x_inst_n391,
         round_inst_S_8__sbox_inst_com_x_inst_n390,
         round_inst_S_8__sbox_inst_com_x_inst_n389,
         round_inst_S_8__sbox_inst_com_x_inst_n388,
         round_inst_S_8__sbox_inst_com_x_inst_n387,
         round_inst_S_8__sbox_inst_com_x_inst_n386,
         round_inst_S_8__sbox_inst_com_x_inst_n385,
         round_inst_S_8__sbox_inst_com_x_inst_n384,
         round_inst_S_8__sbox_inst_com_x_inst_n383,
         round_inst_S_8__sbox_inst_com_x_inst_n382,
         round_inst_S_8__sbox_inst_com_x_inst_n381,
         round_inst_S_8__sbox_inst_com_y_inst_n519,
         round_inst_S_8__sbox_inst_com_y_inst_n518,
         round_inst_S_8__sbox_inst_com_y_inst_n517,
         round_inst_S_8__sbox_inst_com_y_inst_n516,
         round_inst_S_8__sbox_inst_com_y_inst_n515,
         round_inst_S_8__sbox_inst_com_y_inst_n514,
         round_inst_S_8__sbox_inst_com_y_inst_n513,
         round_inst_S_8__sbox_inst_com_y_inst_n512,
         round_inst_S_8__sbox_inst_com_y_inst_n511,
         round_inst_S_8__sbox_inst_com_y_inst_n510,
         round_inst_S_8__sbox_inst_com_y_inst_n509,
         round_inst_S_8__sbox_inst_com_y_inst_n508,
         round_inst_S_8__sbox_inst_com_y_inst_n507,
         round_inst_S_8__sbox_inst_com_y_inst_n506,
         round_inst_S_8__sbox_inst_com_y_inst_n505,
         round_inst_S_8__sbox_inst_com_y_inst_n504,
         round_inst_S_8__sbox_inst_com_y_inst_n503,
         round_inst_S_8__sbox_inst_com_y_inst_n502,
         round_inst_S_8__sbox_inst_com_y_inst_n501,
         round_inst_S_8__sbox_inst_com_y_inst_n500,
         round_inst_S_8__sbox_inst_com_y_inst_n499,
         round_inst_S_8__sbox_inst_com_y_inst_n498,
         round_inst_S_8__sbox_inst_com_y_inst_n497,
         round_inst_S_8__sbox_inst_com_y_inst_n496,
         round_inst_S_8__sbox_inst_com_y_inst_n495,
         round_inst_S_8__sbox_inst_com_y_inst_n494,
         round_inst_S_8__sbox_inst_com_y_inst_n493,
         round_inst_S_8__sbox_inst_com_y_inst_n492,
         round_inst_S_8__sbox_inst_com_y_inst_n491,
         round_inst_S_8__sbox_inst_com_y_inst_n490,
         round_inst_S_8__sbox_inst_com_y_inst_n489,
         round_inst_S_8__sbox_inst_com_y_inst_n488,
         round_inst_S_8__sbox_inst_com_y_inst_n487,
         round_inst_S_8__sbox_inst_com_y_inst_n486,
         round_inst_S_8__sbox_inst_com_y_inst_n485,
         round_inst_S_8__sbox_inst_com_y_inst_n484,
         round_inst_S_8__sbox_inst_com_y_inst_n483,
         round_inst_S_8__sbox_inst_com_y_inst_n482,
         round_inst_S_8__sbox_inst_com_y_inst_n481,
         round_inst_S_8__sbox_inst_com_y_inst_n480,
         round_inst_S_8__sbox_inst_com_y_inst_n479,
         round_inst_S_8__sbox_inst_com_y_inst_n478,
         round_inst_S_8__sbox_inst_com_y_inst_n477,
         round_inst_S_8__sbox_inst_com_y_inst_n476,
         round_inst_S_8__sbox_inst_com_y_inst_n475,
         round_inst_S_8__sbox_inst_com_y_inst_n474,
         round_inst_S_8__sbox_inst_com_y_inst_n473,
         round_inst_S_8__sbox_inst_com_y_inst_n472,
         round_inst_S_8__sbox_inst_com_y_inst_n471,
         round_inst_S_8__sbox_inst_com_y_inst_n470,
         round_inst_S_8__sbox_inst_com_y_inst_n469,
         round_inst_S_8__sbox_inst_com_y_inst_n468,
         round_inst_S_8__sbox_inst_com_y_inst_n467,
         round_inst_S_8__sbox_inst_com_y_inst_n466,
         round_inst_S_8__sbox_inst_com_y_inst_n465,
         round_inst_S_8__sbox_inst_com_y_inst_n464,
         round_inst_S_8__sbox_inst_com_y_inst_n463,
         round_inst_S_8__sbox_inst_com_y_inst_n462,
         round_inst_S_8__sbox_inst_com_y_inst_n461,
         round_inst_S_8__sbox_inst_com_y_inst_n460,
         round_inst_S_8__sbox_inst_com_y_inst_n459,
         round_inst_S_8__sbox_inst_com_y_inst_n458,
         round_inst_S_8__sbox_inst_com_y_inst_n457,
         round_inst_S_8__sbox_inst_com_y_inst_n456,
         round_inst_S_8__sbox_inst_com_y_inst_n455,
         round_inst_S_8__sbox_inst_com_y_inst_n454,
         round_inst_S_8__sbox_inst_com_y_inst_n453,
         round_inst_S_8__sbox_inst_com_y_inst_n452,
         round_inst_S_8__sbox_inst_com_y_inst_n451,
         round_inst_S_8__sbox_inst_com_y_inst_n450,
         round_inst_S_8__sbox_inst_com_y_inst_n449,
         round_inst_S_8__sbox_inst_com_y_inst_n448,
         round_inst_S_8__sbox_inst_com_y_inst_n447,
         round_inst_S_8__sbox_inst_com_y_inst_n446,
         round_inst_S_8__sbox_inst_com_y_inst_n445,
         round_inst_S_8__sbox_inst_com_y_inst_n444,
         round_inst_S_8__sbox_inst_com_y_inst_n443,
         round_inst_S_8__sbox_inst_com_y_inst_n442,
         round_inst_S_8__sbox_inst_com_y_inst_n441,
         round_inst_S_8__sbox_inst_com_y_inst_n440,
         round_inst_S_8__sbox_inst_com_y_inst_n439,
         round_inst_S_8__sbox_inst_com_y_inst_n438,
         round_inst_S_8__sbox_inst_com_y_inst_n437,
         round_inst_S_8__sbox_inst_com_y_inst_n436,
         round_inst_S_8__sbox_inst_com_y_inst_n435,
         round_inst_S_8__sbox_inst_com_y_inst_n434,
         round_inst_S_8__sbox_inst_com_y_inst_n433,
         round_inst_S_8__sbox_inst_com_y_inst_n432,
         round_inst_S_8__sbox_inst_com_y_inst_n431,
         round_inst_S_8__sbox_inst_com_y_inst_n430,
         round_inst_S_8__sbox_inst_com_y_inst_n429,
         round_inst_S_8__sbox_inst_com_y_inst_n428,
         round_inst_S_8__sbox_inst_com_y_inst_n427,
         round_inst_S_8__sbox_inst_com_y_inst_n426,
         round_inst_S_8__sbox_inst_com_y_inst_n425,
         round_inst_S_8__sbox_inst_com_y_inst_n424,
         round_inst_S_8__sbox_inst_com_y_inst_n423,
         round_inst_S_8__sbox_inst_com_y_inst_n422,
         round_inst_S_8__sbox_inst_com_y_inst_n421,
         round_inst_S_8__sbox_inst_com_y_inst_n420,
         round_inst_S_8__sbox_inst_com_y_inst_n419,
         round_inst_S_8__sbox_inst_com_y_inst_n418,
         round_inst_S_8__sbox_inst_com_y_inst_n417,
         round_inst_S_8__sbox_inst_com_y_inst_n416,
         round_inst_S_8__sbox_inst_com_y_inst_n415,
         round_inst_S_8__sbox_inst_com_y_inst_n414,
         round_inst_S_8__sbox_inst_com_y_inst_n413,
         round_inst_S_8__sbox_inst_com_y_inst_n412,
         round_inst_S_8__sbox_inst_com_y_inst_n411,
         round_inst_S_8__sbox_inst_com_y_inst_n410,
         round_inst_S_8__sbox_inst_com_y_inst_n409,
         round_inst_S_8__sbox_inst_com_y_inst_n408,
         round_inst_S_8__sbox_inst_com_y_inst_n407,
         round_inst_S_8__sbox_inst_com_y_inst_n406,
         round_inst_S_8__sbox_inst_com_y_inst_n405,
         round_inst_S_8__sbox_inst_com_y_inst_n404,
         round_inst_S_8__sbox_inst_com_y_inst_n403,
         round_inst_S_8__sbox_inst_com_y_inst_n402,
         round_inst_S_8__sbox_inst_com_y_inst_n401,
         round_inst_S_8__sbox_inst_com_y_inst_n400,
         round_inst_S_8__sbox_inst_com_y_inst_n399,
         round_inst_S_8__sbox_inst_com_y_inst_n398,
         round_inst_S_8__sbox_inst_com_y_inst_n397,
         round_inst_S_8__sbox_inst_com_y_inst_n396,
         round_inst_S_8__sbox_inst_com_y_inst_n395,
         round_inst_S_8__sbox_inst_com_y_inst_n394,
         round_inst_S_8__sbox_inst_com_y_inst_n393,
         round_inst_S_8__sbox_inst_com_y_inst_n392,
         round_inst_S_8__sbox_inst_com_y_inst_n391,
         round_inst_S_8__sbox_inst_com_y_inst_n390,
         round_inst_S_8__sbox_inst_com_y_inst_n389,
         round_inst_S_8__sbox_inst_com_y_inst_n388,
         round_inst_S_8__sbox_inst_com_y_inst_n387,
         round_inst_S_8__sbox_inst_com_y_inst_n386,
         round_inst_S_8__sbox_inst_com_z_inst_n517,
         round_inst_S_8__sbox_inst_com_z_inst_n516,
         round_inst_S_8__sbox_inst_com_z_inst_n515,
         round_inst_S_8__sbox_inst_com_z_inst_n514,
         round_inst_S_8__sbox_inst_com_z_inst_n513,
         round_inst_S_8__sbox_inst_com_z_inst_n512,
         round_inst_S_8__sbox_inst_com_z_inst_n511,
         round_inst_S_8__sbox_inst_com_z_inst_n510,
         round_inst_S_8__sbox_inst_com_z_inst_n509,
         round_inst_S_8__sbox_inst_com_z_inst_n508,
         round_inst_S_8__sbox_inst_com_z_inst_n507,
         round_inst_S_8__sbox_inst_com_z_inst_n506,
         round_inst_S_8__sbox_inst_com_z_inst_n505,
         round_inst_S_8__sbox_inst_com_z_inst_n504,
         round_inst_S_8__sbox_inst_com_z_inst_n503,
         round_inst_S_8__sbox_inst_com_z_inst_n502,
         round_inst_S_8__sbox_inst_com_z_inst_n501,
         round_inst_S_8__sbox_inst_com_z_inst_n500,
         round_inst_S_8__sbox_inst_com_z_inst_n499,
         round_inst_S_8__sbox_inst_com_z_inst_n498,
         round_inst_S_8__sbox_inst_com_z_inst_n497,
         round_inst_S_8__sbox_inst_com_z_inst_n496,
         round_inst_S_8__sbox_inst_com_z_inst_n495,
         round_inst_S_8__sbox_inst_com_z_inst_n494,
         round_inst_S_8__sbox_inst_com_z_inst_n493,
         round_inst_S_8__sbox_inst_com_z_inst_n492,
         round_inst_S_8__sbox_inst_com_z_inst_n491,
         round_inst_S_8__sbox_inst_com_z_inst_n490,
         round_inst_S_8__sbox_inst_com_z_inst_n489,
         round_inst_S_8__sbox_inst_com_z_inst_n488,
         round_inst_S_8__sbox_inst_com_z_inst_n487,
         round_inst_S_8__sbox_inst_com_z_inst_n486,
         round_inst_S_8__sbox_inst_com_z_inst_n485,
         round_inst_S_8__sbox_inst_com_z_inst_n484,
         round_inst_S_8__sbox_inst_com_z_inst_n483,
         round_inst_S_8__sbox_inst_com_z_inst_n482,
         round_inst_S_8__sbox_inst_com_z_inst_n481,
         round_inst_S_8__sbox_inst_com_z_inst_n480,
         round_inst_S_8__sbox_inst_com_z_inst_n479,
         round_inst_S_8__sbox_inst_com_z_inst_n478,
         round_inst_S_8__sbox_inst_com_z_inst_n477,
         round_inst_S_8__sbox_inst_com_z_inst_n476,
         round_inst_S_8__sbox_inst_com_z_inst_n475,
         round_inst_S_8__sbox_inst_com_z_inst_n474,
         round_inst_S_8__sbox_inst_com_z_inst_n473,
         round_inst_S_8__sbox_inst_com_z_inst_n472,
         round_inst_S_8__sbox_inst_com_z_inst_n471,
         round_inst_S_8__sbox_inst_com_z_inst_n470,
         round_inst_S_8__sbox_inst_com_z_inst_n469,
         round_inst_S_8__sbox_inst_com_z_inst_n468,
         round_inst_S_8__sbox_inst_com_z_inst_n467,
         round_inst_S_8__sbox_inst_com_z_inst_n466,
         round_inst_S_8__sbox_inst_com_z_inst_n465,
         round_inst_S_8__sbox_inst_com_z_inst_n464,
         round_inst_S_8__sbox_inst_com_z_inst_n463,
         round_inst_S_8__sbox_inst_com_z_inst_n462,
         round_inst_S_8__sbox_inst_com_z_inst_n461,
         round_inst_S_8__sbox_inst_com_z_inst_n460,
         round_inst_S_8__sbox_inst_com_z_inst_n459,
         round_inst_S_8__sbox_inst_com_z_inst_n458,
         round_inst_S_8__sbox_inst_com_z_inst_n457,
         round_inst_S_8__sbox_inst_com_z_inst_n456,
         round_inst_S_8__sbox_inst_com_z_inst_n455,
         round_inst_S_8__sbox_inst_com_z_inst_n454,
         round_inst_S_8__sbox_inst_com_z_inst_n453,
         round_inst_S_8__sbox_inst_com_z_inst_n452,
         round_inst_S_8__sbox_inst_com_z_inst_n451,
         round_inst_S_8__sbox_inst_com_z_inst_n450,
         round_inst_S_8__sbox_inst_com_z_inst_n449,
         round_inst_S_8__sbox_inst_com_z_inst_n448,
         round_inst_S_8__sbox_inst_com_z_inst_n447,
         round_inst_S_8__sbox_inst_com_z_inst_n446,
         round_inst_S_8__sbox_inst_com_z_inst_n445,
         round_inst_S_8__sbox_inst_com_z_inst_n444,
         round_inst_S_8__sbox_inst_com_z_inst_n443,
         round_inst_S_8__sbox_inst_com_z_inst_n442,
         round_inst_S_8__sbox_inst_com_z_inst_n441,
         round_inst_S_8__sbox_inst_com_z_inst_n440,
         round_inst_S_8__sbox_inst_com_z_inst_n439,
         round_inst_S_8__sbox_inst_com_z_inst_n438,
         round_inst_S_8__sbox_inst_com_z_inst_n437,
         round_inst_S_8__sbox_inst_com_z_inst_n436,
         round_inst_S_8__sbox_inst_com_z_inst_n435,
         round_inst_S_8__sbox_inst_com_z_inst_n434,
         round_inst_S_8__sbox_inst_com_z_inst_n433,
         round_inst_S_8__sbox_inst_com_z_inst_n432,
         round_inst_S_8__sbox_inst_com_z_inst_n431,
         round_inst_S_8__sbox_inst_com_z_inst_n430,
         round_inst_S_8__sbox_inst_com_z_inst_n429,
         round_inst_S_8__sbox_inst_com_z_inst_n428,
         round_inst_S_8__sbox_inst_com_z_inst_n427,
         round_inst_S_8__sbox_inst_com_z_inst_n426,
         round_inst_S_8__sbox_inst_com_z_inst_n425,
         round_inst_S_8__sbox_inst_com_z_inst_n424,
         round_inst_S_8__sbox_inst_com_z_inst_n423,
         round_inst_S_8__sbox_inst_com_z_inst_n422,
         round_inst_S_8__sbox_inst_com_z_inst_n421,
         round_inst_S_8__sbox_inst_com_z_inst_n420,
         round_inst_S_8__sbox_inst_com_z_inst_n419,
         round_inst_S_8__sbox_inst_com_z_inst_n418,
         round_inst_S_8__sbox_inst_com_z_inst_n417,
         round_inst_S_8__sbox_inst_com_z_inst_n416,
         round_inst_S_8__sbox_inst_com_z_inst_n415,
         round_inst_S_8__sbox_inst_com_z_inst_n414,
         round_inst_S_8__sbox_inst_com_z_inst_n413,
         round_inst_S_8__sbox_inst_com_z_inst_n412,
         round_inst_S_8__sbox_inst_com_z_inst_n411,
         round_inst_S_8__sbox_inst_com_z_inst_n410,
         round_inst_S_8__sbox_inst_com_z_inst_n409,
         round_inst_S_8__sbox_inst_com_z_inst_n408,
         round_inst_S_8__sbox_inst_com_z_inst_n407,
         round_inst_S_8__sbox_inst_com_z_inst_n406,
         round_inst_S_8__sbox_inst_com_z_inst_n405,
         round_inst_S_8__sbox_inst_com_z_inst_n404,
         round_inst_S_8__sbox_inst_com_z_inst_n403,
         round_inst_S_8__sbox_inst_com_z_inst_n402,
         round_inst_S_8__sbox_inst_com_z_inst_n401,
         round_inst_S_8__sbox_inst_com_z_inst_n400,
         round_inst_S_8__sbox_inst_com_z_inst_n399,
         round_inst_S_8__sbox_inst_com_z_inst_n398,
         round_inst_S_8__sbox_inst_com_z_inst_n397,
         round_inst_S_8__sbox_inst_com_z_inst_n396,
         round_inst_S_8__sbox_inst_com_z_inst_n395,
         round_inst_S_8__sbox_inst_com_z_inst_n394,
         round_inst_S_8__sbox_inst_com_z_inst_n393,
         round_inst_S_8__sbox_inst_com_z_inst_n392,
         round_inst_S_8__sbox_inst_com_z_inst_n391,
         round_inst_S_8__sbox_inst_com_z_inst_n390,
         round_inst_S_9__sbox_inst_n10, round_inst_S_9__sbox_inst_n9,
         round_inst_S_9__sbox_inst_n8, round_inst_S_9__sbox_inst_n7,
         round_inst_S_9__sbox_inst_n6, round_inst_S_9__sbox_inst_n5,
         round_inst_S_9__sbox_inst_n4, round_inst_S_9__sbox_inst_n3,
         round_inst_S_9__sbox_inst_n2, round_inst_S_9__sbox_inst_n1,
         round_inst_S_9__sbox_inst_com_w_inst_n532,
         round_inst_S_9__sbox_inst_com_w_inst_n531,
         round_inst_S_9__sbox_inst_com_w_inst_n530,
         round_inst_S_9__sbox_inst_com_w_inst_n529,
         round_inst_S_9__sbox_inst_com_w_inst_n528,
         round_inst_S_9__sbox_inst_com_w_inst_n527,
         round_inst_S_9__sbox_inst_com_w_inst_n526,
         round_inst_S_9__sbox_inst_com_w_inst_n525,
         round_inst_S_9__sbox_inst_com_w_inst_n524,
         round_inst_S_9__sbox_inst_com_w_inst_n523,
         round_inst_S_9__sbox_inst_com_w_inst_n522,
         round_inst_S_9__sbox_inst_com_w_inst_n521,
         round_inst_S_9__sbox_inst_com_w_inst_n520,
         round_inst_S_9__sbox_inst_com_w_inst_n519,
         round_inst_S_9__sbox_inst_com_w_inst_n518,
         round_inst_S_9__sbox_inst_com_w_inst_n517,
         round_inst_S_9__sbox_inst_com_w_inst_n516,
         round_inst_S_9__sbox_inst_com_w_inst_n515,
         round_inst_S_9__sbox_inst_com_w_inst_n514,
         round_inst_S_9__sbox_inst_com_w_inst_n513,
         round_inst_S_9__sbox_inst_com_w_inst_n512,
         round_inst_S_9__sbox_inst_com_w_inst_n511,
         round_inst_S_9__sbox_inst_com_w_inst_n510,
         round_inst_S_9__sbox_inst_com_w_inst_n509,
         round_inst_S_9__sbox_inst_com_w_inst_n508,
         round_inst_S_9__sbox_inst_com_w_inst_n507,
         round_inst_S_9__sbox_inst_com_w_inst_n506,
         round_inst_S_9__sbox_inst_com_w_inst_n505,
         round_inst_S_9__sbox_inst_com_w_inst_n504,
         round_inst_S_9__sbox_inst_com_w_inst_n503,
         round_inst_S_9__sbox_inst_com_w_inst_n502,
         round_inst_S_9__sbox_inst_com_w_inst_n501,
         round_inst_S_9__sbox_inst_com_w_inst_n500,
         round_inst_S_9__sbox_inst_com_w_inst_n499,
         round_inst_S_9__sbox_inst_com_w_inst_n498,
         round_inst_S_9__sbox_inst_com_w_inst_n497,
         round_inst_S_9__sbox_inst_com_w_inst_n496,
         round_inst_S_9__sbox_inst_com_w_inst_n495,
         round_inst_S_9__sbox_inst_com_w_inst_n494,
         round_inst_S_9__sbox_inst_com_w_inst_n493,
         round_inst_S_9__sbox_inst_com_w_inst_n492,
         round_inst_S_9__sbox_inst_com_w_inst_n491,
         round_inst_S_9__sbox_inst_com_w_inst_n490,
         round_inst_S_9__sbox_inst_com_w_inst_n489,
         round_inst_S_9__sbox_inst_com_w_inst_n488,
         round_inst_S_9__sbox_inst_com_w_inst_n487,
         round_inst_S_9__sbox_inst_com_w_inst_n486,
         round_inst_S_9__sbox_inst_com_w_inst_n485,
         round_inst_S_9__sbox_inst_com_w_inst_n484,
         round_inst_S_9__sbox_inst_com_w_inst_n483,
         round_inst_S_9__sbox_inst_com_w_inst_n482,
         round_inst_S_9__sbox_inst_com_w_inst_n481,
         round_inst_S_9__sbox_inst_com_w_inst_n480,
         round_inst_S_9__sbox_inst_com_w_inst_n479,
         round_inst_S_9__sbox_inst_com_w_inst_n478,
         round_inst_S_9__sbox_inst_com_w_inst_n477,
         round_inst_S_9__sbox_inst_com_w_inst_n476,
         round_inst_S_9__sbox_inst_com_w_inst_n475,
         round_inst_S_9__sbox_inst_com_w_inst_n474,
         round_inst_S_9__sbox_inst_com_w_inst_n473,
         round_inst_S_9__sbox_inst_com_w_inst_n472,
         round_inst_S_9__sbox_inst_com_w_inst_n471,
         round_inst_S_9__sbox_inst_com_w_inst_n470,
         round_inst_S_9__sbox_inst_com_w_inst_n469,
         round_inst_S_9__sbox_inst_com_w_inst_n468,
         round_inst_S_9__sbox_inst_com_w_inst_n467,
         round_inst_S_9__sbox_inst_com_w_inst_n466,
         round_inst_S_9__sbox_inst_com_w_inst_n465,
         round_inst_S_9__sbox_inst_com_w_inst_n464,
         round_inst_S_9__sbox_inst_com_w_inst_n463,
         round_inst_S_9__sbox_inst_com_w_inst_n462,
         round_inst_S_9__sbox_inst_com_w_inst_n461,
         round_inst_S_9__sbox_inst_com_w_inst_n460,
         round_inst_S_9__sbox_inst_com_w_inst_n459,
         round_inst_S_9__sbox_inst_com_w_inst_n458,
         round_inst_S_9__sbox_inst_com_w_inst_n457,
         round_inst_S_9__sbox_inst_com_w_inst_n456,
         round_inst_S_9__sbox_inst_com_w_inst_n455,
         round_inst_S_9__sbox_inst_com_w_inst_n454,
         round_inst_S_9__sbox_inst_com_w_inst_n453,
         round_inst_S_9__sbox_inst_com_w_inst_n452,
         round_inst_S_9__sbox_inst_com_w_inst_n451,
         round_inst_S_9__sbox_inst_com_w_inst_n450,
         round_inst_S_9__sbox_inst_com_w_inst_n449,
         round_inst_S_9__sbox_inst_com_w_inst_n448,
         round_inst_S_9__sbox_inst_com_w_inst_n447,
         round_inst_S_9__sbox_inst_com_w_inst_n446,
         round_inst_S_9__sbox_inst_com_w_inst_n445,
         round_inst_S_9__sbox_inst_com_w_inst_n444,
         round_inst_S_9__sbox_inst_com_w_inst_n443,
         round_inst_S_9__sbox_inst_com_w_inst_n442,
         round_inst_S_9__sbox_inst_com_w_inst_n441,
         round_inst_S_9__sbox_inst_com_w_inst_n440,
         round_inst_S_9__sbox_inst_com_w_inst_n439,
         round_inst_S_9__sbox_inst_com_w_inst_n438,
         round_inst_S_9__sbox_inst_com_w_inst_n437,
         round_inst_S_9__sbox_inst_com_w_inst_n436,
         round_inst_S_9__sbox_inst_com_w_inst_n435,
         round_inst_S_9__sbox_inst_com_w_inst_n434,
         round_inst_S_9__sbox_inst_com_w_inst_n433,
         round_inst_S_9__sbox_inst_com_w_inst_n432,
         round_inst_S_9__sbox_inst_com_w_inst_n431,
         round_inst_S_9__sbox_inst_com_w_inst_n430,
         round_inst_S_9__sbox_inst_com_w_inst_n429,
         round_inst_S_9__sbox_inst_com_w_inst_n428,
         round_inst_S_9__sbox_inst_com_w_inst_n427,
         round_inst_S_9__sbox_inst_com_w_inst_n426,
         round_inst_S_9__sbox_inst_com_w_inst_n425,
         round_inst_S_9__sbox_inst_com_w_inst_n424,
         round_inst_S_9__sbox_inst_com_w_inst_n423,
         round_inst_S_9__sbox_inst_com_w_inst_n422,
         round_inst_S_9__sbox_inst_com_w_inst_n421,
         round_inst_S_9__sbox_inst_com_w_inst_n420,
         round_inst_S_9__sbox_inst_com_w_inst_n419,
         round_inst_S_9__sbox_inst_com_w_inst_n418,
         round_inst_S_9__sbox_inst_com_w_inst_n417,
         round_inst_S_9__sbox_inst_com_w_inst_n416,
         round_inst_S_9__sbox_inst_com_w_inst_n415,
         round_inst_S_9__sbox_inst_com_w_inst_n414,
         round_inst_S_9__sbox_inst_com_w_inst_n413,
         round_inst_S_9__sbox_inst_com_w_inst_n412,
         round_inst_S_9__sbox_inst_com_w_inst_n411,
         round_inst_S_9__sbox_inst_com_w_inst_n410,
         round_inst_S_9__sbox_inst_com_w_inst_n409,
         round_inst_S_9__sbox_inst_com_w_inst_n408,
         round_inst_S_9__sbox_inst_com_w_inst_n407,
         round_inst_S_9__sbox_inst_com_w_inst_n406,
         round_inst_S_9__sbox_inst_com_w_inst_n405,
         round_inst_S_9__sbox_inst_com_w_inst_n404,
         round_inst_S_9__sbox_inst_com_w_inst_n403,
         round_inst_S_9__sbox_inst_com_w_inst_n402,
         round_inst_S_9__sbox_inst_com_w_inst_n401,
         round_inst_S_9__sbox_inst_com_w_inst_n400,
         round_inst_S_9__sbox_inst_com_w_inst_n399,
         round_inst_S_9__sbox_inst_com_w_inst_n398,
         round_inst_S_9__sbox_inst_com_w_inst_n397,
         round_inst_S_9__sbox_inst_com_w_inst_n396,
         round_inst_S_9__sbox_inst_com_x_inst_n511,
         round_inst_S_9__sbox_inst_com_x_inst_n510,
         round_inst_S_9__sbox_inst_com_x_inst_n509,
         round_inst_S_9__sbox_inst_com_x_inst_n508,
         round_inst_S_9__sbox_inst_com_x_inst_n507,
         round_inst_S_9__sbox_inst_com_x_inst_n506,
         round_inst_S_9__sbox_inst_com_x_inst_n505,
         round_inst_S_9__sbox_inst_com_x_inst_n504,
         round_inst_S_9__sbox_inst_com_x_inst_n503,
         round_inst_S_9__sbox_inst_com_x_inst_n502,
         round_inst_S_9__sbox_inst_com_x_inst_n501,
         round_inst_S_9__sbox_inst_com_x_inst_n500,
         round_inst_S_9__sbox_inst_com_x_inst_n499,
         round_inst_S_9__sbox_inst_com_x_inst_n498,
         round_inst_S_9__sbox_inst_com_x_inst_n497,
         round_inst_S_9__sbox_inst_com_x_inst_n496,
         round_inst_S_9__sbox_inst_com_x_inst_n495,
         round_inst_S_9__sbox_inst_com_x_inst_n494,
         round_inst_S_9__sbox_inst_com_x_inst_n493,
         round_inst_S_9__sbox_inst_com_x_inst_n492,
         round_inst_S_9__sbox_inst_com_x_inst_n491,
         round_inst_S_9__sbox_inst_com_x_inst_n490,
         round_inst_S_9__sbox_inst_com_x_inst_n489,
         round_inst_S_9__sbox_inst_com_x_inst_n488,
         round_inst_S_9__sbox_inst_com_x_inst_n487,
         round_inst_S_9__sbox_inst_com_x_inst_n486,
         round_inst_S_9__sbox_inst_com_x_inst_n485,
         round_inst_S_9__sbox_inst_com_x_inst_n484,
         round_inst_S_9__sbox_inst_com_x_inst_n483,
         round_inst_S_9__sbox_inst_com_x_inst_n482,
         round_inst_S_9__sbox_inst_com_x_inst_n481,
         round_inst_S_9__sbox_inst_com_x_inst_n480,
         round_inst_S_9__sbox_inst_com_x_inst_n479,
         round_inst_S_9__sbox_inst_com_x_inst_n478,
         round_inst_S_9__sbox_inst_com_x_inst_n477,
         round_inst_S_9__sbox_inst_com_x_inst_n476,
         round_inst_S_9__sbox_inst_com_x_inst_n475,
         round_inst_S_9__sbox_inst_com_x_inst_n474,
         round_inst_S_9__sbox_inst_com_x_inst_n473,
         round_inst_S_9__sbox_inst_com_x_inst_n472,
         round_inst_S_9__sbox_inst_com_x_inst_n471,
         round_inst_S_9__sbox_inst_com_x_inst_n470,
         round_inst_S_9__sbox_inst_com_x_inst_n469,
         round_inst_S_9__sbox_inst_com_x_inst_n468,
         round_inst_S_9__sbox_inst_com_x_inst_n467,
         round_inst_S_9__sbox_inst_com_x_inst_n466,
         round_inst_S_9__sbox_inst_com_x_inst_n465,
         round_inst_S_9__sbox_inst_com_x_inst_n464,
         round_inst_S_9__sbox_inst_com_x_inst_n463,
         round_inst_S_9__sbox_inst_com_x_inst_n462,
         round_inst_S_9__sbox_inst_com_x_inst_n461,
         round_inst_S_9__sbox_inst_com_x_inst_n460,
         round_inst_S_9__sbox_inst_com_x_inst_n459,
         round_inst_S_9__sbox_inst_com_x_inst_n458,
         round_inst_S_9__sbox_inst_com_x_inst_n457,
         round_inst_S_9__sbox_inst_com_x_inst_n456,
         round_inst_S_9__sbox_inst_com_x_inst_n455,
         round_inst_S_9__sbox_inst_com_x_inst_n454,
         round_inst_S_9__sbox_inst_com_x_inst_n453,
         round_inst_S_9__sbox_inst_com_x_inst_n452,
         round_inst_S_9__sbox_inst_com_x_inst_n451,
         round_inst_S_9__sbox_inst_com_x_inst_n450,
         round_inst_S_9__sbox_inst_com_x_inst_n449,
         round_inst_S_9__sbox_inst_com_x_inst_n448,
         round_inst_S_9__sbox_inst_com_x_inst_n447,
         round_inst_S_9__sbox_inst_com_x_inst_n446,
         round_inst_S_9__sbox_inst_com_x_inst_n445,
         round_inst_S_9__sbox_inst_com_x_inst_n444,
         round_inst_S_9__sbox_inst_com_x_inst_n443,
         round_inst_S_9__sbox_inst_com_x_inst_n442,
         round_inst_S_9__sbox_inst_com_x_inst_n441,
         round_inst_S_9__sbox_inst_com_x_inst_n440,
         round_inst_S_9__sbox_inst_com_x_inst_n439,
         round_inst_S_9__sbox_inst_com_x_inst_n438,
         round_inst_S_9__sbox_inst_com_x_inst_n437,
         round_inst_S_9__sbox_inst_com_x_inst_n436,
         round_inst_S_9__sbox_inst_com_x_inst_n435,
         round_inst_S_9__sbox_inst_com_x_inst_n434,
         round_inst_S_9__sbox_inst_com_x_inst_n433,
         round_inst_S_9__sbox_inst_com_x_inst_n432,
         round_inst_S_9__sbox_inst_com_x_inst_n431,
         round_inst_S_9__sbox_inst_com_x_inst_n430,
         round_inst_S_9__sbox_inst_com_x_inst_n429,
         round_inst_S_9__sbox_inst_com_x_inst_n428,
         round_inst_S_9__sbox_inst_com_x_inst_n427,
         round_inst_S_9__sbox_inst_com_x_inst_n426,
         round_inst_S_9__sbox_inst_com_x_inst_n425,
         round_inst_S_9__sbox_inst_com_x_inst_n424,
         round_inst_S_9__sbox_inst_com_x_inst_n423,
         round_inst_S_9__sbox_inst_com_x_inst_n422,
         round_inst_S_9__sbox_inst_com_x_inst_n421,
         round_inst_S_9__sbox_inst_com_x_inst_n420,
         round_inst_S_9__sbox_inst_com_x_inst_n419,
         round_inst_S_9__sbox_inst_com_x_inst_n418,
         round_inst_S_9__sbox_inst_com_x_inst_n417,
         round_inst_S_9__sbox_inst_com_x_inst_n416,
         round_inst_S_9__sbox_inst_com_x_inst_n415,
         round_inst_S_9__sbox_inst_com_x_inst_n414,
         round_inst_S_9__sbox_inst_com_x_inst_n413,
         round_inst_S_9__sbox_inst_com_x_inst_n412,
         round_inst_S_9__sbox_inst_com_x_inst_n411,
         round_inst_S_9__sbox_inst_com_x_inst_n410,
         round_inst_S_9__sbox_inst_com_x_inst_n409,
         round_inst_S_9__sbox_inst_com_x_inst_n408,
         round_inst_S_9__sbox_inst_com_x_inst_n407,
         round_inst_S_9__sbox_inst_com_x_inst_n406,
         round_inst_S_9__sbox_inst_com_x_inst_n405,
         round_inst_S_9__sbox_inst_com_x_inst_n404,
         round_inst_S_9__sbox_inst_com_x_inst_n403,
         round_inst_S_9__sbox_inst_com_x_inst_n402,
         round_inst_S_9__sbox_inst_com_x_inst_n401,
         round_inst_S_9__sbox_inst_com_x_inst_n400,
         round_inst_S_9__sbox_inst_com_x_inst_n399,
         round_inst_S_9__sbox_inst_com_x_inst_n398,
         round_inst_S_9__sbox_inst_com_x_inst_n397,
         round_inst_S_9__sbox_inst_com_x_inst_n396,
         round_inst_S_9__sbox_inst_com_x_inst_n395,
         round_inst_S_9__sbox_inst_com_x_inst_n394,
         round_inst_S_9__sbox_inst_com_x_inst_n393,
         round_inst_S_9__sbox_inst_com_x_inst_n392,
         round_inst_S_9__sbox_inst_com_x_inst_n391,
         round_inst_S_9__sbox_inst_com_x_inst_n390,
         round_inst_S_9__sbox_inst_com_x_inst_n389,
         round_inst_S_9__sbox_inst_com_x_inst_n388,
         round_inst_S_9__sbox_inst_com_x_inst_n387,
         round_inst_S_9__sbox_inst_com_x_inst_n386,
         round_inst_S_9__sbox_inst_com_x_inst_n385,
         round_inst_S_9__sbox_inst_com_x_inst_n384,
         round_inst_S_9__sbox_inst_com_x_inst_n383,
         round_inst_S_9__sbox_inst_com_x_inst_n382,
         round_inst_S_9__sbox_inst_com_x_inst_n381,
         round_inst_S_9__sbox_inst_com_y_inst_n518,
         round_inst_S_9__sbox_inst_com_y_inst_n517,
         round_inst_S_9__sbox_inst_com_y_inst_n516,
         round_inst_S_9__sbox_inst_com_y_inst_n515,
         round_inst_S_9__sbox_inst_com_y_inst_n514,
         round_inst_S_9__sbox_inst_com_y_inst_n513,
         round_inst_S_9__sbox_inst_com_y_inst_n512,
         round_inst_S_9__sbox_inst_com_y_inst_n511,
         round_inst_S_9__sbox_inst_com_y_inst_n510,
         round_inst_S_9__sbox_inst_com_y_inst_n509,
         round_inst_S_9__sbox_inst_com_y_inst_n508,
         round_inst_S_9__sbox_inst_com_y_inst_n507,
         round_inst_S_9__sbox_inst_com_y_inst_n506,
         round_inst_S_9__sbox_inst_com_y_inst_n505,
         round_inst_S_9__sbox_inst_com_y_inst_n504,
         round_inst_S_9__sbox_inst_com_y_inst_n503,
         round_inst_S_9__sbox_inst_com_y_inst_n502,
         round_inst_S_9__sbox_inst_com_y_inst_n501,
         round_inst_S_9__sbox_inst_com_y_inst_n500,
         round_inst_S_9__sbox_inst_com_y_inst_n499,
         round_inst_S_9__sbox_inst_com_y_inst_n498,
         round_inst_S_9__sbox_inst_com_y_inst_n497,
         round_inst_S_9__sbox_inst_com_y_inst_n496,
         round_inst_S_9__sbox_inst_com_y_inst_n495,
         round_inst_S_9__sbox_inst_com_y_inst_n494,
         round_inst_S_9__sbox_inst_com_y_inst_n493,
         round_inst_S_9__sbox_inst_com_y_inst_n492,
         round_inst_S_9__sbox_inst_com_y_inst_n491,
         round_inst_S_9__sbox_inst_com_y_inst_n490,
         round_inst_S_9__sbox_inst_com_y_inst_n489,
         round_inst_S_9__sbox_inst_com_y_inst_n488,
         round_inst_S_9__sbox_inst_com_y_inst_n487,
         round_inst_S_9__sbox_inst_com_y_inst_n486,
         round_inst_S_9__sbox_inst_com_y_inst_n485,
         round_inst_S_9__sbox_inst_com_y_inst_n484,
         round_inst_S_9__sbox_inst_com_y_inst_n483,
         round_inst_S_9__sbox_inst_com_y_inst_n482,
         round_inst_S_9__sbox_inst_com_y_inst_n481,
         round_inst_S_9__sbox_inst_com_y_inst_n480,
         round_inst_S_9__sbox_inst_com_y_inst_n479,
         round_inst_S_9__sbox_inst_com_y_inst_n478,
         round_inst_S_9__sbox_inst_com_y_inst_n477,
         round_inst_S_9__sbox_inst_com_y_inst_n476,
         round_inst_S_9__sbox_inst_com_y_inst_n475,
         round_inst_S_9__sbox_inst_com_y_inst_n474,
         round_inst_S_9__sbox_inst_com_y_inst_n473,
         round_inst_S_9__sbox_inst_com_y_inst_n472,
         round_inst_S_9__sbox_inst_com_y_inst_n471,
         round_inst_S_9__sbox_inst_com_y_inst_n470,
         round_inst_S_9__sbox_inst_com_y_inst_n469,
         round_inst_S_9__sbox_inst_com_y_inst_n468,
         round_inst_S_9__sbox_inst_com_y_inst_n467,
         round_inst_S_9__sbox_inst_com_y_inst_n466,
         round_inst_S_9__sbox_inst_com_y_inst_n465,
         round_inst_S_9__sbox_inst_com_y_inst_n464,
         round_inst_S_9__sbox_inst_com_y_inst_n463,
         round_inst_S_9__sbox_inst_com_y_inst_n462,
         round_inst_S_9__sbox_inst_com_y_inst_n461,
         round_inst_S_9__sbox_inst_com_y_inst_n460,
         round_inst_S_9__sbox_inst_com_y_inst_n459,
         round_inst_S_9__sbox_inst_com_y_inst_n458,
         round_inst_S_9__sbox_inst_com_y_inst_n457,
         round_inst_S_9__sbox_inst_com_y_inst_n456,
         round_inst_S_9__sbox_inst_com_y_inst_n455,
         round_inst_S_9__sbox_inst_com_y_inst_n454,
         round_inst_S_9__sbox_inst_com_y_inst_n453,
         round_inst_S_9__sbox_inst_com_y_inst_n452,
         round_inst_S_9__sbox_inst_com_y_inst_n451,
         round_inst_S_9__sbox_inst_com_y_inst_n450,
         round_inst_S_9__sbox_inst_com_y_inst_n449,
         round_inst_S_9__sbox_inst_com_y_inst_n448,
         round_inst_S_9__sbox_inst_com_y_inst_n447,
         round_inst_S_9__sbox_inst_com_y_inst_n446,
         round_inst_S_9__sbox_inst_com_y_inst_n445,
         round_inst_S_9__sbox_inst_com_y_inst_n444,
         round_inst_S_9__sbox_inst_com_y_inst_n443,
         round_inst_S_9__sbox_inst_com_y_inst_n442,
         round_inst_S_9__sbox_inst_com_y_inst_n441,
         round_inst_S_9__sbox_inst_com_y_inst_n440,
         round_inst_S_9__sbox_inst_com_y_inst_n439,
         round_inst_S_9__sbox_inst_com_y_inst_n438,
         round_inst_S_9__sbox_inst_com_y_inst_n437,
         round_inst_S_9__sbox_inst_com_y_inst_n436,
         round_inst_S_9__sbox_inst_com_y_inst_n435,
         round_inst_S_9__sbox_inst_com_y_inst_n434,
         round_inst_S_9__sbox_inst_com_y_inst_n433,
         round_inst_S_9__sbox_inst_com_y_inst_n432,
         round_inst_S_9__sbox_inst_com_y_inst_n431,
         round_inst_S_9__sbox_inst_com_y_inst_n430,
         round_inst_S_9__sbox_inst_com_y_inst_n429,
         round_inst_S_9__sbox_inst_com_y_inst_n428,
         round_inst_S_9__sbox_inst_com_y_inst_n427,
         round_inst_S_9__sbox_inst_com_y_inst_n426,
         round_inst_S_9__sbox_inst_com_y_inst_n425,
         round_inst_S_9__sbox_inst_com_y_inst_n424,
         round_inst_S_9__sbox_inst_com_y_inst_n423,
         round_inst_S_9__sbox_inst_com_y_inst_n422,
         round_inst_S_9__sbox_inst_com_y_inst_n421,
         round_inst_S_9__sbox_inst_com_y_inst_n420,
         round_inst_S_9__sbox_inst_com_y_inst_n419,
         round_inst_S_9__sbox_inst_com_y_inst_n418,
         round_inst_S_9__sbox_inst_com_y_inst_n417,
         round_inst_S_9__sbox_inst_com_y_inst_n416,
         round_inst_S_9__sbox_inst_com_y_inst_n415,
         round_inst_S_9__sbox_inst_com_y_inst_n414,
         round_inst_S_9__sbox_inst_com_y_inst_n413,
         round_inst_S_9__sbox_inst_com_y_inst_n412,
         round_inst_S_9__sbox_inst_com_y_inst_n411,
         round_inst_S_9__sbox_inst_com_y_inst_n410,
         round_inst_S_9__sbox_inst_com_y_inst_n409,
         round_inst_S_9__sbox_inst_com_y_inst_n408,
         round_inst_S_9__sbox_inst_com_y_inst_n407,
         round_inst_S_9__sbox_inst_com_y_inst_n406,
         round_inst_S_9__sbox_inst_com_y_inst_n405,
         round_inst_S_9__sbox_inst_com_y_inst_n404,
         round_inst_S_9__sbox_inst_com_y_inst_n403,
         round_inst_S_9__sbox_inst_com_y_inst_n402,
         round_inst_S_9__sbox_inst_com_y_inst_n401,
         round_inst_S_9__sbox_inst_com_y_inst_n400,
         round_inst_S_9__sbox_inst_com_y_inst_n399,
         round_inst_S_9__sbox_inst_com_y_inst_n398,
         round_inst_S_9__sbox_inst_com_y_inst_n397,
         round_inst_S_9__sbox_inst_com_y_inst_n396,
         round_inst_S_9__sbox_inst_com_y_inst_n395,
         round_inst_S_9__sbox_inst_com_y_inst_n394,
         round_inst_S_9__sbox_inst_com_y_inst_n393,
         round_inst_S_9__sbox_inst_com_y_inst_n392,
         round_inst_S_9__sbox_inst_com_y_inst_n391,
         round_inst_S_9__sbox_inst_com_y_inst_n390,
         round_inst_S_9__sbox_inst_com_y_inst_n389,
         round_inst_S_9__sbox_inst_com_y_inst_n388,
         round_inst_S_9__sbox_inst_com_y_inst_n387,
         round_inst_S_9__sbox_inst_com_y_inst_n386,
         round_inst_S_9__sbox_inst_com_z_inst_n516,
         round_inst_S_9__sbox_inst_com_z_inst_n515,
         round_inst_S_9__sbox_inst_com_z_inst_n514,
         round_inst_S_9__sbox_inst_com_z_inst_n513,
         round_inst_S_9__sbox_inst_com_z_inst_n512,
         round_inst_S_9__sbox_inst_com_z_inst_n511,
         round_inst_S_9__sbox_inst_com_z_inst_n510,
         round_inst_S_9__sbox_inst_com_z_inst_n509,
         round_inst_S_9__sbox_inst_com_z_inst_n508,
         round_inst_S_9__sbox_inst_com_z_inst_n507,
         round_inst_S_9__sbox_inst_com_z_inst_n506,
         round_inst_S_9__sbox_inst_com_z_inst_n505,
         round_inst_S_9__sbox_inst_com_z_inst_n504,
         round_inst_S_9__sbox_inst_com_z_inst_n503,
         round_inst_S_9__sbox_inst_com_z_inst_n502,
         round_inst_S_9__sbox_inst_com_z_inst_n501,
         round_inst_S_9__sbox_inst_com_z_inst_n500,
         round_inst_S_9__sbox_inst_com_z_inst_n499,
         round_inst_S_9__sbox_inst_com_z_inst_n498,
         round_inst_S_9__sbox_inst_com_z_inst_n497,
         round_inst_S_9__sbox_inst_com_z_inst_n496,
         round_inst_S_9__sbox_inst_com_z_inst_n495,
         round_inst_S_9__sbox_inst_com_z_inst_n494,
         round_inst_S_9__sbox_inst_com_z_inst_n493,
         round_inst_S_9__sbox_inst_com_z_inst_n492,
         round_inst_S_9__sbox_inst_com_z_inst_n491,
         round_inst_S_9__sbox_inst_com_z_inst_n490,
         round_inst_S_9__sbox_inst_com_z_inst_n489,
         round_inst_S_9__sbox_inst_com_z_inst_n488,
         round_inst_S_9__sbox_inst_com_z_inst_n487,
         round_inst_S_9__sbox_inst_com_z_inst_n486,
         round_inst_S_9__sbox_inst_com_z_inst_n485,
         round_inst_S_9__sbox_inst_com_z_inst_n484,
         round_inst_S_9__sbox_inst_com_z_inst_n483,
         round_inst_S_9__sbox_inst_com_z_inst_n482,
         round_inst_S_9__sbox_inst_com_z_inst_n481,
         round_inst_S_9__sbox_inst_com_z_inst_n480,
         round_inst_S_9__sbox_inst_com_z_inst_n479,
         round_inst_S_9__sbox_inst_com_z_inst_n478,
         round_inst_S_9__sbox_inst_com_z_inst_n477,
         round_inst_S_9__sbox_inst_com_z_inst_n476,
         round_inst_S_9__sbox_inst_com_z_inst_n475,
         round_inst_S_9__sbox_inst_com_z_inst_n474,
         round_inst_S_9__sbox_inst_com_z_inst_n473,
         round_inst_S_9__sbox_inst_com_z_inst_n472,
         round_inst_S_9__sbox_inst_com_z_inst_n471,
         round_inst_S_9__sbox_inst_com_z_inst_n470,
         round_inst_S_9__sbox_inst_com_z_inst_n469,
         round_inst_S_9__sbox_inst_com_z_inst_n468,
         round_inst_S_9__sbox_inst_com_z_inst_n467,
         round_inst_S_9__sbox_inst_com_z_inst_n466,
         round_inst_S_9__sbox_inst_com_z_inst_n465,
         round_inst_S_9__sbox_inst_com_z_inst_n464,
         round_inst_S_9__sbox_inst_com_z_inst_n463,
         round_inst_S_9__sbox_inst_com_z_inst_n462,
         round_inst_S_9__sbox_inst_com_z_inst_n461,
         round_inst_S_9__sbox_inst_com_z_inst_n460,
         round_inst_S_9__sbox_inst_com_z_inst_n459,
         round_inst_S_9__sbox_inst_com_z_inst_n458,
         round_inst_S_9__sbox_inst_com_z_inst_n457,
         round_inst_S_9__sbox_inst_com_z_inst_n456,
         round_inst_S_9__sbox_inst_com_z_inst_n455,
         round_inst_S_9__sbox_inst_com_z_inst_n454,
         round_inst_S_9__sbox_inst_com_z_inst_n453,
         round_inst_S_9__sbox_inst_com_z_inst_n452,
         round_inst_S_9__sbox_inst_com_z_inst_n451,
         round_inst_S_9__sbox_inst_com_z_inst_n450,
         round_inst_S_9__sbox_inst_com_z_inst_n449,
         round_inst_S_9__sbox_inst_com_z_inst_n448,
         round_inst_S_9__sbox_inst_com_z_inst_n447,
         round_inst_S_9__sbox_inst_com_z_inst_n446,
         round_inst_S_9__sbox_inst_com_z_inst_n445,
         round_inst_S_9__sbox_inst_com_z_inst_n444,
         round_inst_S_9__sbox_inst_com_z_inst_n443,
         round_inst_S_9__sbox_inst_com_z_inst_n442,
         round_inst_S_9__sbox_inst_com_z_inst_n441,
         round_inst_S_9__sbox_inst_com_z_inst_n440,
         round_inst_S_9__sbox_inst_com_z_inst_n439,
         round_inst_S_9__sbox_inst_com_z_inst_n438,
         round_inst_S_9__sbox_inst_com_z_inst_n437,
         round_inst_S_9__sbox_inst_com_z_inst_n436,
         round_inst_S_9__sbox_inst_com_z_inst_n435,
         round_inst_S_9__sbox_inst_com_z_inst_n434,
         round_inst_S_9__sbox_inst_com_z_inst_n433,
         round_inst_S_9__sbox_inst_com_z_inst_n432,
         round_inst_S_9__sbox_inst_com_z_inst_n431,
         round_inst_S_9__sbox_inst_com_z_inst_n430,
         round_inst_S_9__sbox_inst_com_z_inst_n429,
         round_inst_S_9__sbox_inst_com_z_inst_n428,
         round_inst_S_9__sbox_inst_com_z_inst_n427,
         round_inst_S_9__sbox_inst_com_z_inst_n426,
         round_inst_S_9__sbox_inst_com_z_inst_n425,
         round_inst_S_9__sbox_inst_com_z_inst_n424,
         round_inst_S_9__sbox_inst_com_z_inst_n423,
         round_inst_S_9__sbox_inst_com_z_inst_n422,
         round_inst_S_9__sbox_inst_com_z_inst_n421,
         round_inst_S_9__sbox_inst_com_z_inst_n420,
         round_inst_S_9__sbox_inst_com_z_inst_n419,
         round_inst_S_9__sbox_inst_com_z_inst_n418,
         round_inst_S_9__sbox_inst_com_z_inst_n417,
         round_inst_S_9__sbox_inst_com_z_inst_n416,
         round_inst_S_9__sbox_inst_com_z_inst_n415,
         round_inst_S_9__sbox_inst_com_z_inst_n414,
         round_inst_S_9__sbox_inst_com_z_inst_n413,
         round_inst_S_9__sbox_inst_com_z_inst_n412,
         round_inst_S_9__sbox_inst_com_z_inst_n411,
         round_inst_S_9__sbox_inst_com_z_inst_n410,
         round_inst_S_9__sbox_inst_com_z_inst_n409,
         round_inst_S_9__sbox_inst_com_z_inst_n408,
         round_inst_S_9__sbox_inst_com_z_inst_n407,
         round_inst_S_9__sbox_inst_com_z_inst_n406,
         round_inst_S_9__sbox_inst_com_z_inst_n405,
         round_inst_S_9__sbox_inst_com_z_inst_n404,
         round_inst_S_9__sbox_inst_com_z_inst_n403,
         round_inst_S_9__sbox_inst_com_z_inst_n402,
         round_inst_S_9__sbox_inst_com_z_inst_n401,
         round_inst_S_9__sbox_inst_com_z_inst_n400,
         round_inst_S_9__sbox_inst_com_z_inst_n399,
         round_inst_S_9__sbox_inst_com_z_inst_n398,
         round_inst_S_9__sbox_inst_com_z_inst_n397,
         round_inst_S_9__sbox_inst_com_z_inst_n396,
         round_inst_S_9__sbox_inst_com_z_inst_n395,
         round_inst_S_9__sbox_inst_com_z_inst_n394,
         round_inst_S_9__sbox_inst_com_z_inst_n393,
         round_inst_S_9__sbox_inst_com_z_inst_n392,
         round_inst_S_9__sbox_inst_com_z_inst_n391,
         round_inst_S_9__sbox_inst_com_z_inst_n390,
         round_inst_S_9__sbox_inst_com_z_inst_n389,
         round_inst_S_10__sbox_inst_n6, round_inst_S_10__sbox_inst_n5,
         round_inst_S_10__sbox_inst_n4, round_inst_S_10__sbox_inst_n3,
         round_inst_S_10__sbox_inst_n2, round_inst_S_10__sbox_inst_n1,
         round_inst_S_10__sbox_inst_com_w_inst_n532,
         round_inst_S_10__sbox_inst_com_w_inst_n531,
         round_inst_S_10__sbox_inst_com_w_inst_n530,
         round_inst_S_10__sbox_inst_com_w_inst_n529,
         round_inst_S_10__sbox_inst_com_w_inst_n528,
         round_inst_S_10__sbox_inst_com_w_inst_n527,
         round_inst_S_10__sbox_inst_com_w_inst_n526,
         round_inst_S_10__sbox_inst_com_w_inst_n525,
         round_inst_S_10__sbox_inst_com_w_inst_n524,
         round_inst_S_10__sbox_inst_com_w_inst_n523,
         round_inst_S_10__sbox_inst_com_w_inst_n522,
         round_inst_S_10__sbox_inst_com_w_inst_n521,
         round_inst_S_10__sbox_inst_com_w_inst_n520,
         round_inst_S_10__sbox_inst_com_w_inst_n519,
         round_inst_S_10__sbox_inst_com_w_inst_n518,
         round_inst_S_10__sbox_inst_com_w_inst_n517,
         round_inst_S_10__sbox_inst_com_w_inst_n516,
         round_inst_S_10__sbox_inst_com_w_inst_n515,
         round_inst_S_10__sbox_inst_com_w_inst_n514,
         round_inst_S_10__sbox_inst_com_w_inst_n513,
         round_inst_S_10__sbox_inst_com_w_inst_n512,
         round_inst_S_10__sbox_inst_com_w_inst_n511,
         round_inst_S_10__sbox_inst_com_w_inst_n510,
         round_inst_S_10__sbox_inst_com_w_inst_n509,
         round_inst_S_10__sbox_inst_com_w_inst_n508,
         round_inst_S_10__sbox_inst_com_w_inst_n507,
         round_inst_S_10__sbox_inst_com_w_inst_n506,
         round_inst_S_10__sbox_inst_com_w_inst_n505,
         round_inst_S_10__sbox_inst_com_w_inst_n504,
         round_inst_S_10__sbox_inst_com_w_inst_n503,
         round_inst_S_10__sbox_inst_com_w_inst_n502,
         round_inst_S_10__sbox_inst_com_w_inst_n501,
         round_inst_S_10__sbox_inst_com_w_inst_n500,
         round_inst_S_10__sbox_inst_com_w_inst_n499,
         round_inst_S_10__sbox_inst_com_w_inst_n498,
         round_inst_S_10__sbox_inst_com_w_inst_n497,
         round_inst_S_10__sbox_inst_com_w_inst_n496,
         round_inst_S_10__sbox_inst_com_w_inst_n495,
         round_inst_S_10__sbox_inst_com_w_inst_n494,
         round_inst_S_10__sbox_inst_com_w_inst_n493,
         round_inst_S_10__sbox_inst_com_w_inst_n492,
         round_inst_S_10__sbox_inst_com_w_inst_n491,
         round_inst_S_10__sbox_inst_com_w_inst_n490,
         round_inst_S_10__sbox_inst_com_w_inst_n489,
         round_inst_S_10__sbox_inst_com_w_inst_n488,
         round_inst_S_10__sbox_inst_com_w_inst_n487,
         round_inst_S_10__sbox_inst_com_w_inst_n486,
         round_inst_S_10__sbox_inst_com_w_inst_n485,
         round_inst_S_10__sbox_inst_com_w_inst_n484,
         round_inst_S_10__sbox_inst_com_w_inst_n483,
         round_inst_S_10__sbox_inst_com_w_inst_n482,
         round_inst_S_10__sbox_inst_com_w_inst_n481,
         round_inst_S_10__sbox_inst_com_w_inst_n480,
         round_inst_S_10__sbox_inst_com_w_inst_n479,
         round_inst_S_10__sbox_inst_com_w_inst_n478,
         round_inst_S_10__sbox_inst_com_w_inst_n477,
         round_inst_S_10__sbox_inst_com_w_inst_n476,
         round_inst_S_10__sbox_inst_com_w_inst_n475,
         round_inst_S_10__sbox_inst_com_w_inst_n474,
         round_inst_S_10__sbox_inst_com_w_inst_n473,
         round_inst_S_10__sbox_inst_com_w_inst_n472,
         round_inst_S_10__sbox_inst_com_w_inst_n471,
         round_inst_S_10__sbox_inst_com_w_inst_n470,
         round_inst_S_10__sbox_inst_com_w_inst_n469,
         round_inst_S_10__sbox_inst_com_w_inst_n468,
         round_inst_S_10__sbox_inst_com_w_inst_n467,
         round_inst_S_10__sbox_inst_com_w_inst_n466,
         round_inst_S_10__sbox_inst_com_w_inst_n465,
         round_inst_S_10__sbox_inst_com_w_inst_n464,
         round_inst_S_10__sbox_inst_com_w_inst_n463,
         round_inst_S_10__sbox_inst_com_w_inst_n462,
         round_inst_S_10__sbox_inst_com_w_inst_n461,
         round_inst_S_10__sbox_inst_com_w_inst_n460,
         round_inst_S_10__sbox_inst_com_w_inst_n459,
         round_inst_S_10__sbox_inst_com_w_inst_n458,
         round_inst_S_10__sbox_inst_com_w_inst_n457,
         round_inst_S_10__sbox_inst_com_w_inst_n456,
         round_inst_S_10__sbox_inst_com_w_inst_n455,
         round_inst_S_10__sbox_inst_com_w_inst_n454,
         round_inst_S_10__sbox_inst_com_w_inst_n453,
         round_inst_S_10__sbox_inst_com_w_inst_n452,
         round_inst_S_10__sbox_inst_com_w_inst_n451,
         round_inst_S_10__sbox_inst_com_w_inst_n450,
         round_inst_S_10__sbox_inst_com_w_inst_n449,
         round_inst_S_10__sbox_inst_com_w_inst_n448,
         round_inst_S_10__sbox_inst_com_w_inst_n447,
         round_inst_S_10__sbox_inst_com_w_inst_n446,
         round_inst_S_10__sbox_inst_com_w_inst_n445,
         round_inst_S_10__sbox_inst_com_w_inst_n444,
         round_inst_S_10__sbox_inst_com_w_inst_n443,
         round_inst_S_10__sbox_inst_com_w_inst_n442,
         round_inst_S_10__sbox_inst_com_w_inst_n441,
         round_inst_S_10__sbox_inst_com_w_inst_n440,
         round_inst_S_10__sbox_inst_com_w_inst_n439,
         round_inst_S_10__sbox_inst_com_w_inst_n438,
         round_inst_S_10__sbox_inst_com_w_inst_n437,
         round_inst_S_10__sbox_inst_com_w_inst_n436,
         round_inst_S_10__sbox_inst_com_w_inst_n435,
         round_inst_S_10__sbox_inst_com_w_inst_n434,
         round_inst_S_10__sbox_inst_com_w_inst_n433,
         round_inst_S_10__sbox_inst_com_w_inst_n432,
         round_inst_S_10__sbox_inst_com_w_inst_n431,
         round_inst_S_10__sbox_inst_com_w_inst_n430,
         round_inst_S_10__sbox_inst_com_w_inst_n429,
         round_inst_S_10__sbox_inst_com_w_inst_n428,
         round_inst_S_10__sbox_inst_com_w_inst_n427,
         round_inst_S_10__sbox_inst_com_w_inst_n426,
         round_inst_S_10__sbox_inst_com_w_inst_n425,
         round_inst_S_10__sbox_inst_com_w_inst_n424,
         round_inst_S_10__sbox_inst_com_w_inst_n423,
         round_inst_S_10__sbox_inst_com_w_inst_n422,
         round_inst_S_10__sbox_inst_com_w_inst_n421,
         round_inst_S_10__sbox_inst_com_w_inst_n420,
         round_inst_S_10__sbox_inst_com_w_inst_n419,
         round_inst_S_10__sbox_inst_com_w_inst_n418,
         round_inst_S_10__sbox_inst_com_w_inst_n417,
         round_inst_S_10__sbox_inst_com_w_inst_n416,
         round_inst_S_10__sbox_inst_com_w_inst_n415,
         round_inst_S_10__sbox_inst_com_w_inst_n414,
         round_inst_S_10__sbox_inst_com_w_inst_n413,
         round_inst_S_10__sbox_inst_com_w_inst_n412,
         round_inst_S_10__sbox_inst_com_w_inst_n411,
         round_inst_S_10__sbox_inst_com_w_inst_n410,
         round_inst_S_10__sbox_inst_com_w_inst_n409,
         round_inst_S_10__sbox_inst_com_w_inst_n408,
         round_inst_S_10__sbox_inst_com_w_inst_n407,
         round_inst_S_10__sbox_inst_com_w_inst_n406,
         round_inst_S_10__sbox_inst_com_w_inst_n405,
         round_inst_S_10__sbox_inst_com_w_inst_n404,
         round_inst_S_10__sbox_inst_com_w_inst_n403,
         round_inst_S_10__sbox_inst_com_w_inst_n402,
         round_inst_S_10__sbox_inst_com_w_inst_n401,
         round_inst_S_10__sbox_inst_com_w_inst_n400,
         round_inst_S_10__sbox_inst_com_w_inst_n399,
         round_inst_S_10__sbox_inst_com_w_inst_n398,
         round_inst_S_10__sbox_inst_com_w_inst_n397,
         round_inst_S_10__sbox_inst_com_w_inst_n396,
         round_inst_S_10__sbox_inst_com_x_inst_n519,
         round_inst_S_10__sbox_inst_com_x_inst_n518,
         round_inst_S_10__sbox_inst_com_x_inst_n517,
         round_inst_S_10__sbox_inst_com_x_inst_n516,
         round_inst_S_10__sbox_inst_com_x_inst_n515,
         round_inst_S_10__sbox_inst_com_x_inst_n514,
         round_inst_S_10__sbox_inst_com_x_inst_n513,
         round_inst_S_10__sbox_inst_com_x_inst_n512,
         round_inst_S_10__sbox_inst_com_x_inst_n511,
         round_inst_S_10__sbox_inst_com_x_inst_n510,
         round_inst_S_10__sbox_inst_com_x_inst_n509,
         round_inst_S_10__sbox_inst_com_x_inst_n508,
         round_inst_S_10__sbox_inst_com_x_inst_n507,
         round_inst_S_10__sbox_inst_com_x_inst_n506,
         round_inst_S_10__sbox_inst_com_x_inst_n505,
         round_inst_S_10__sbox_inst_com_x_inst_n504,
         round_inst_S_10__sbox_inst_com_x_inst_n503,
         round_inst_S_10__sbox_inst_com_x_inst_n502,
         round_inst_S_10__sbox_inst_com_x_inst_n501,
         round_inst_S_10__sbox_inst_com_x_inst_n500,
         round_inst_S_10__sbox_inst_com_x_inst_n499,
         round_inst_S_10__sbox_inst_com_x_inst_n498,
         round_inst_S_10__sbox_inst_com_x_inst_n497,
         round_inst_S_10__sbox_inst_com_x_inst_n496,
         round_inst_S_10__sbox_inst_com_x_inst_n495,
         round_inst_S_10__sbox_inst_com_x_inst_n494,
         round_inst_S_10__sbox_inst_com_x_inst_n493,
         round_inst_S_10__sbox_inst_com_x_inst_n492,
         round_inst_S_10__sbox_inst_com_x_inst_n491,
         round_inst_S_10__sbox_inst_com_x_inst_n490,
         round_inst_S_10__sbox_inst_com_x_inst_n489,
         round_inst_S_10__sbox_inst_com_x_inst_n488,
         round_inst_S_10__sbox_inst_com_x_inst_n487,
         round_inst_S_10__sbox_inst_com_x_inst_n486,
         round_inst_S_10__sbox_inst_com_x_inst_n485,
         round_inst_S_10__sbox_inst_com_x_inst_n484,
         round_inst_S_10__sbox_inst_com_x_inst_n483,
         round_inst_S_10__sbox_inst_com_x_inst_n482,
         round_inst_S_10__sbox_inst_com_x_inst_n481,
         round_inst_S_10__sbox_inst_com_x_inst_n480,
         round_inst_S_10__sbox_inst_com_x_inst_n479,
         round_inst_S_10__sbox_inst_com_x_inst_n478,
         round_inst_S_10__sbox_inst_com_x_inst_n477,
         round_inst_S_10__sbox_inst_com_x_inst_n476,
         round_inst_S_10__sbox_inst_com_x_inst_n475,
         round_inst_S_10__sbox_inst_com_x_inst_n474,
         round_inst_S_10__sbox_inst_com_x_inst_n473,
         round_inst_S_10__sbox_inst_com_x_inst_n472,
         round_inst_S_10__sbox_inst_com_x_inst_n471,
         round_inst_S_10__sbox_inst_com_x_inst_n470,
         round_inst_S_10__sbox_inst_com_x_inst_n469,
         round_inst_S_10__sbox_inst_com_x_inst_n468,
         round_inst_S_10__sbox_inst_com_x_inst_n467,
         round_inst_S_10__sbox_inst_com_x_inst_n466,
         round_inst_S_10__sbox_inst_com_x_inst_n465,
         round_inst_S_10__sbox_inst_com_x_inst_n464,
         round_inst_S_10__sbox_inst_com_x_inst_n463,
         round_inst_S_10__sbox_inst_com_x_inst_n462,
         round_inst_S_10__sbox_inst_com_x_inst_n461,
         round_inst_S_10__sbox_inst_com_x_inst_n460,
         round_inst_S_10__sbox_inst_com_x_inst_n459,
         round_inst_S_10__sbox_inst_com_x_inst_n458,
         round_inst_S_10__sbox_inst_com_x_inst_n457,
         round_inst_S_10__sbox_inst_com_x_inst_n456,
         round_inst_S_10__sbox_inst_com_x_inst_n455,
         round_inst_S_10__sbox_inst_com_x_inst_n454,
         round_inst_S_10__sbox_inst_com_x_inst_n453,
         round_inst_S_10__sbox_inst_com_x_inst_n452,
         round_inst_S_10__sbox_inst_com_x_inst_n451,
         round_inst_S_10__sbox_inst_com_x_inst_n450,
         round_inst_S_10__sbox_inst_com_x_inst_n449,
         round_inst_S_10__sbox_inst_com_x_inst_n448,
         round_inst_S_10__sbox_inst_com_x_inst_n447,
         round_inst_S_10__sbox_inst_com_x_inst_n446,
         round_inst_S_10__sbox_inst_com_x_inst_n445,
         round_inst_S_10__sbox_inst_com_x_inst_n444,
         round_inst_S_10__sbox_inst_com_x_inst_n443,
         round_inst_S_10__sbox_inst_com_x_inst_n442,
         round_inst_S_10__sbox_inst_com_x_inst_n441,
         round_inst_S_10__sbox_inst_com_x_inst_n440,
         round_inst_S_10__sbox_inst_com_x_inst_n439,
         round_inst_S_10__sbox_inst_com_x_inst_n438,
         round_inst_S_10__sbox_inst_com_x_inst_n437,
         round_inst_S_10__sbox_inst_com_x_inst_n436,
         round_inst_S_10__sbox_inst_com_x_inst_n435,
         round_inst_S_10__sbox_inst_com_x_inst_n434,
         round_inst_S_10__sbox_inst_com_x_inst_n433,
         round_inst_S_10__sbox_inst_com_x_inst_n432,
         round_inst_S_10__sbox_inst_com_x_inst_n431,
         round_inst_S_10__sbox_inst_com_x_inst_n430,
         round_inst_S_10__sbox_inst_com_x_inst_n429,
         round_inst_S_10__sbox_inst_com_x_inst_n428,
         round_inst_S_10__sbox_inst_com_x_inst_n427,
         round_inst_S_10__sbox_inst_com_x_inst_n426,
         round_inst_S_10__sbox_inst_com_x_inst_n425,
         round_inst_S_10__sbox_inst_com_x_inst_n424,
         round_inst_S_10__sbox_inst_com_x_inst_n423,
         round_inst_S_10__sbox_inst_com_x_inst_n422,
         round_inst_S_10__sbox_inst_com_x_inst_n421,
         round_inst_S_10__sbox_inst_com_x_inst_n420,
         round_inst_S_10__sbox_inst_com_x_inst_n419,
         round_inst_S_10__sbox_inst_com_x_inst_n418,
         round_inst_S_10__sbox_inst_com_x_inst_n417,
         round_inst_S_10__sbox_inst_com_x_inst_n416,
         round_inst_S_10__sbox_inst_com_x_inst_n415,
         round_inst_S_10__sbox_inst_com_x_inst_n414,
         round_inst_S_10__sbox_inst_com_x_inst_n413,
         round_inst_S_10__sbox_inst_com_x_inst_n412,
         round_inst_S_10__sbox_inst_com_x_inst_n411,
         round_inst_S_10__sbox_inst_com_x_inst_n410,
         round_inst_S_10__sbox_inst_com_x_inst_n409,
         round_inst_S_10__sbox_inst_com_x_inst_n408,
         round_inst_S_10__sbox_inst_com_x_inst_n407,
         round_inst_S_10__sbox_inst_com_x_inst_n406,
         round_inst_S_10__sbox_inst_com_x_inst_n405,
         round_inst_S_10__sbox_inst_com_x_inst_n404,
         round_inst_S_10__sbox_inst_com_x_inst_n403,
         round_inst_S_10__sbox_inst_com_x_inst_n402,
         round_inst_S_10__sbox_inst_com_x_inst_n401,
         round_inst_S_10__sbox_inst_com_x_inst_n400,
         round_inst_S_10__sbox_inst_com_x_inst_n399,
         round_inst_S_10__sbox_inst_com_x_inst_n398,
         round_inst_S_10__sbox_inst_com_x_inst_n397,
         round_inst_S_10__sbox_inst_com_x_inst_n396,
         round_inst_S_10__sbox_inst_com_x_inst_n395,
         round_inst_S_10__sbox_inst_com_x_inst_n394,
         round_inst_S_10__sbox_inst_com_x_inst_n393,
         round_inst_S_10__sbox_inst_com_x_inst_n392,
         round_inst_S_10__sbox_inst_com_x_inst_n391,
         round_inst_S_10__sbox_inst_com_x_inst_n390,
         round_inst_S_10__sbox_inst_com_x_inst_n389,
         round_inst_S_10__sbox_inst_com_x_inst_n388,
         round_inst_S_10__sbox_inst_com_x_inst_n387,
         round_inst_S_10__sbox_inst_com_x_inst_n386,
         round_inst_S_10__sbox_inst_com_x_inst_n385,
         round_inst_S_10__sbox_inst_com_x_inst_n384,
         round_inst_S_10__sbox_inst_com_x_inst_n383,
         round_inst_S_10__sbox_inst_com_x_inst_n382,
         round_inst_S_10__sbox_inst_com_x_inst_n381,
         round_inst_S_10__sbox_inst_com_x_inst_n380,
         round_inst_S_10__sbox_inst_com_y_inst_n517,
         round_inst_S_10__sbox_inst_com_y_inst_n516,
         round_inst_S_10__sbox_inst_com_y_inst_n515,
         round_inst_S_10__sbox_inst_com_y_inst_n514,
         round_inst_S_10__sbox_inst_com_y_inst_n513,
         round_inst_S_10__sbox_inst_com_y_inst_n512,
         round_inst_S_10__sbox_inst_com_y_inst_n511,
         round_inst_S_10__sbox_inst_com_y_inst_n510,
         round_inst_S_10__sbox_inst_com_y_inst_n509,
         round_inst_S_10__sbox_inst_com_y_inst_n508,
         round_inst_S_10__sbox_inst_com_y_inst_n507,
         round_inst_S_10__sbox_inst_com_y_inst_n506,
         round_inst_S_10__sbox_inst_com_y_inst_n505,
         round_inst_S_10__sbox_inst_com_y_inst_n504,
         round_inst_S_10__sbox_inst_com_y_inst_n503,
         round_inst_S_10__sbox_inst_com_y_inst_n502,
         round_inst_S_10__sbox_inst_com_y_inst_n501,
         round_inst_S_10__sbox_inst_com_y_inst_n500,
         round_inst_S_10__sbox_inst_com_y_inst_n499,
         round_inst_S_10__sbox_inst_com_y_inst_n498,
         round_inst_S_10__sbox_inst_com_y_inst_n497,
         round_inst_S_10__sbox_inst_com_y_inst_n496,
         round_inst_S_10__sbox_inst_com_y_inst_n495,
         round_inst_S_10__sbox_inst_com_y_inst_n494,
         round_inst_S_10__sbox_inst_com_y_inst_n493,
         round_inst_S_10__sbox_inst_com_y_inst_n492,
         round_inst_S_10__sbox_inst_com_y_inst_n491,
         round_inst_S_10__sbox_inst_com_y_inst_n490,
         round_inst_S_10__sbox_inst_com_y_inst_n489,
         round_inst_S_10__sbox_inst_com_y_inst_n488,
         round_inst_S_10__sbox_inst_com_y_inst_n487,
         round_inst_S_10__sbox_inst_com_y_inst_n486,
         round_inst_S_10__sbox_inst_com_y_inst_n485,
         round_inst_S_10__sbox_inst_com_y_inst_n484,
         round_inst_S_10__sbox_inst_com_y_inst_n483,
         round_inst_S_10__sbox_inst_com_y_inst_n482,
         round_inst_S_10__sbox_inst_com_y_inst_n481,
         round_inst_S_10__sbox_inst_com_y_inst_n480,
         round_inst_S_10__sbox_inst_com_y_inst_n479,
         round_inst_S_10__sbox_inst_com_y_inst_n478,
         round_inst_S_10__sbox_inst_com_y_inst_n477,
         round_inst_S_10__sbox_inst_com_y_inst_n476,
         round_inst_S_10__sbox_inst_com_y_inst_n475,
         round_inst_S_10__sbox_inst_com_y_inst_n474,
         round_inst_S_10__sbox_inst_com_y_inst_n473,
         round_inst_S_10__sbox_inst_com_y_inst_n472,
         round_inst_S_10__sbox_inst_com_y_inst_n471,
         round_inst_S_10__sbox_inst_com_y_inst_n470,
         round_inst_S_10__sbox_inst_com_y_inst_n469,
         round_inst_S_10__sbox_inst_com_y_inst_n468,
         round_inst_S_10__sbox_inst_com_y_inst_n467,
         round_inst_S_10__sbox_inst_com_y_inst_n466,
         round_inst_S_10__sbox_inst_com_y_inst_n465,
         round_inst_S_10__sbox_inst_com_y_inst_n464,
         round_inst_S_10__sbox_inst_com_y_inst_n463,
         round_inst_S_10__sbox_inst_com_y_inst_n462,
         round_inst_S_10__sbox_inst_com_y_inst_n461,
         round_inst_S_10__sbox_inst_com_y_inst_n460,
         round_inst_S_10__sbox_inst_com_y_inst_n459,
         round_inst_S_10__sbox_inst_com_y_inst_n458,
         round_inst_S_10__sbox_inst_com_y_inst_n457,
         round_inst_S_10__sbox_inst_com_y_inst_n456,
         round_inst_S_10__sbox_inst_com_y_inst_n455,
         round_inst_S_10__sbox_inst_com_y_inst_n454,
         round_inst_S_10__sbox_inst_com_y_inst_n453,
         round_inst_S_10__sbox_inst_com_y_inst_n452,
         round_inst_S_10__sbox_inst_com_y_inst_n451,
         round_inst_S_10__sbox_inst_com_y_inst_n450,
         round_inst_S_10__sbox_inst_com_y_inst_n449,
         round_inst_S_10__sbox_inst_com_y_inst_n448,
         round_inst_S_10__sbox_inst_com_y_inst_n447,
         round_inst_S_10__sbox_inst_com_y_inst_n446,
         round_inst_S_10__sbox_inst_com_y_inst_n445,
         round_inst_S_10__sbox_inst_com_y_inst_n444,
         round_inst_S_10__sbox_inst_com_y_inst_n443,
         round_inst_S_10__sbox_inst_com_y_inst_n442,
         round_inst_S_10__sbox_inst_com_y_inst_n441,
         round_inst_S_10__sbox_inst_com_y_inst_n440,
         round_inst_S_10__sbox_inst_com_y_inst_n439,
         round_inst_S_10__sbox_inst_com_y_inst_n438,
         round_inst_S_10__sbox_inst_com_y_inst_n437,
         round_inst_S_10__sbox_inst_com_y_inst_n436,
         round_inst_S_10__sbox_inst_com_y_inst_n435,
         round_inst_S_10__sbox_inst_com_y_inst_n434,
         round_inst_S_10__sbox_inst_com_y_inst_n433,
         round_inst_S_10__sbox_inst_com_y_inst_n432,
         round_inst_S_10__sbox_inst_com_y_inst_n431,
         round_inst_S_10__sbox_inst_com_y_inst_n430,
         round_inst_S_10__sbox_inst_com_y_inst_n429,
         round_inst_S_10__sbox_inst_com_y_inst_n428,
         round_inst_S_10__sbox_inst_com_y_inst_n427,
         round_inst_S_10__sbox_inst_com_y_inst_n426,
         round_inst_S_10__sbox_inst_com_y_inst_n425,
         round_inst_S_10__sbox_inst_com_y_inst_n424,
         round_inst_S_10__sbox_inst_com_y_inst_n423,
         round_inst_S_10__sbox_inst_com_y_inst_n422,
         round_inst_S_10__sbox_inst_com_y_inst_n421,
         round_inst_S_10__sbox_inst_com_y_inst_n420,
         round_inst_S_10__sbox_inst_com_y_inst_n419,
         round_inst_S_10__sbox_inst_com_y_inst_n418,
         round_inst_S_10__sbox_inst_com_y_inst_n417,
         round_inst_S_10__sbox_inst_com_y_inst_n416,
         round_inst_S_10__sbox_inst_com_y_inst_n415,
         round_inst_S_10__sbox_inst_com_y_inst_n414,
         round_inst_S_10__sbox_inst_com_y_inst_n413,
         round_inst_S_10__sbox_inst_com_y_inst_n412,
         round_inst_S_10__sbox_inst_com_y_inst_n411,
         round_inst_S_10__sbox_inst_com_y_inst_n410,
         round_inst_S_10__sbox_inst_com_y_inst_n409,
         round_inst_S_10__sbox_inst_com_y_inst_n408,
         round_inst_S_10__sbox_inst_com_y_inst_n407,
         round_inst_S_10__sbox_inst_com_y_inst_n406,
         round_inst_S_10__sbox_inst_com_y_inst_n405,
         round_inst_S_10__sbox_inst_com_y_inst_n404,
         round_inst_S_10__sbox_inst_com_y_inst_n403,
         round_inst_S_10__sbox_inst_com_y_inst_n402,
         round_inst_S_10__sbox_inst_com_y_inst_n401,
         round_inst_S_10__sbox_inst_com_y_inst_n400,
         round_inst_S_10__sbox_inst_com_y_inst_n399,
         round_inst_S_10__sbox_inst_com_y_inst_n398,
         round_inst_S_10__sbox_inst_com_y_inst_n397,
         round_inst_S_10__sbox_inst_com_y_inst_n396,
         round_inst_S_10__sbox_inst_com_y_inst_n395,
         round_inst_S_10__sbox_inst_com_y_inst_n394,
         round_inst_S_10__sbox_inst_com_y_inst_n393,
         round_inst_S_10__sbox_inst_com_y_inst_n392,
         round_inst_S_10__sbox_inst_com_y_inst_n391,
         round_inst_S_10__sbox_inst_com_y_inst_n390,
         round_inst_S_10__sbox_inst_com_y_inst_n389,
         round_inst_S_10__sbox_inst_com_y_inst_n388,
         round_inst_S_10__sbox_inst_com_y_inst_n387,
         round_inst_S_10__sbox_inst_com_y_inst_n386,
         round_inst_S_10__sbox_inst_com_z_inst_n523,
         round_inst_S_10__sbox_inst_com_z_inst_n522,
         round_inst_S_10__sbox_inst_com_z_inst_n521,
         round_inst_S_10__sbox_inst_com_z_inst_n520,
         round_inst_S_10__sbox_inst_com_z_inst_n519,
         round_inst_S_10__sbox_inst_com_z_inst_n518,
         round_inst_S_10__sbox_inst_com_z_inst_n517,
         round_inst_S_10__sbox_inst_com_z_inst_n516,
         round_inst_S_10__sbox_inst_com_z_inst_n515,
         round_inst_S_10__sbox_inst_com_z_inst_n514,
         round_inst_S_10__sbox_inst_com_z_inst_n513,
         round_inst_S_10__sbox_inst_com_z_inst_n512,
         round_inst_S_10__sbox_inst_com_z_inst_n511,
         round_inst_S_10__sbox_inst_com_z_inst_n510,
         round_inst_S_10__sbox_inst_com_z_inst_n509,
         round_inst_S_10__sbox_inst_com_z_inst_n508,
         round_inst_S_10__sbox_inst_com_z_inst_n507,
         round_inst_S_10__sbox_inst_com_z_inst_n506,
         round_inst_S_10__sbox_inst_com_z_inst_n505,
         round_inst_S_10__sbox_inst_com_z_inst_n504,
         round_inst_S_10__sbox_inst_com_z_inst_n503,
         round_inst_S_10__sbox_inst_com_z_inst_n502,
         round_inst_S_10__sbox_inst_com_z_inst_n501,
         round_inst_S_10__sbox_inst_com_z_inst_n500,
         round_inst_S_10__sbox_inst_com_z_inst_n499,
         round_inst_S_10__sbox_inst_com_z_inst_n498,
         round_inst_S_10__sbox_inst_com_z_inst_n497,
         round_inst_S_10__sbox_inst_com_z_inst_n496,
         round_inst_S_10__sbox_inst_com_z_inst_n495,
         round_inst_S_10__sbox_inst_com_z_inst_n494,
         round_inst_S_10__sbox_inst_com_z_inst_n493,
         round_inst_S_10__sbox_inst_com_z_inst_n492,
         round_inst_S_10__sbox_inst_com_z_inst_n491,
         round_inst_S_10__sbox_inst_com_z_inst_n490,
         round_inst_S_10__sbox_inst_com_z_inst_n489,
         round_inst_S_10__sbox_inst_com_z_inst_n488,
         round_inst_S_10__sbox_inst_com_z_inst_n487,
         round_inst_S_10__sbox_inst_com_z_inst_n486,
         round_inst_S_10__sbox_inst_com_z_inst_n485,
         round_inst_S_10__sbox_inst_com_z_inst_n484,
         round_inst_S_10__sbox_inst_com_z_inst_n483,
         round_inst_S_10__sbox_inst_com_z_inst_n482,
         round_inst_S_10__sbox_inst_com_z_inst_n481,
         round_inst_S_10__sbox_inst_com_z_inst_n480,
         round_inst_S_10__sbox_inst_com_z_inst_n479,
         round_inst_S_10__sbox_inst_com_z_inst_n478,
         round_inst_S_10__sbox_inst_com_z_inst_n477,
         round_inst_S_10__sbox_inst_com_z_inst_n476,
         round_inst_S_10__sbox_inst_com_z_inst_n475,
         round_inst_S_10__sbox_inst_com_z_inst_n474,
         round_inst_S_10__sbox_inst_com_z_inst_n473,
         round_inst_S_10__sbox_inst_com_z_inst_n472,
         round_inst_S_10__sbox_inst_com_z_inst_n471,
         round_inst_S_10__sbox_inst_com_z_inst_n470,
         round_inst_S_10__sbox_inst_com_z_inst_n469,
         round_inst_S_10__sbox_inst_com_z_inst_n468,
         round_inst_S_10__sbox_inst_com_z_inst_n467,
         round_inst_S_10__sbox_inst_com_z_inst_n466,
         round_inst_S_10__sbox_inst_com_z_inst_n465,
         round_inst_S_10__sbox_inst_com_z_inst_n464,
         round_inst_S_10__sbox_inst_com_z_inst_n463,
         round_inst_S_10__sbox_inst_com_z_inst_n462,
         round_inst_S_10__sbox_inst_com_z_inst_n461,
         round_inst_S_10__sbox_inst_com_z_inst_n460,
         round_inst_S_10__sbox_inst_com_z_inst_n459,
         round_inst_S_10__sbox_inst_com_z_inst_n458,
         round_inst_S_10__sbox_inst_com_z_inst_n457,
         round_inst_S_10__sbox_inst_com_z_inst_n456,
         round_inst_S_10__sbox_inst_com_z_inst_n455,
         round_inst_S_10__sbox_inst_com_z_inst_n454,
         round_inst_S_10__sbox_inst_com_z_inst_n453,
         round_inst_S_10__sbox_inst_com_z_inst_n452,
         round_inst_S_10__sbox_inst_com_z_inst_n451,
         round_inst_S_10__sbox_inst_com_z_inst_n450,
         round_inst_S_10__sbox_inst_com_z_inst_n449,
         round_inst_S_10__sbox_inst_com_z_inst_n448,
         round_inst_S_10__sbox_inst_com_z_inst_n447,
         round_inst_S_10__sbox_inst_com_z_inst_n446,
         round_inst_S_10__sbox_inst_com_z_inst_n445,
         round_inst_S_10__sbox_inst_com_z_inst_n444,
         round_inst_S_10__sbox_inst_com_z_inst_n443,
         round_inst_S_10__sbox_inst_com_z_inst_n442,
         round_inst_S_10__sbox_inst_com_z_inst_n441,
         round_inst_S_10__sbox_inst_com_z_inst_n440,
         round_inst_S_10__sbox_inst_com_z_inst_n439,
         round_inst_S_10__sbox_inst_com_z_inst_n438,
         round_inst_S_10__sbox_inst_com_z_inst_n437,
         round_inst_S_10__sbox_inst_com_z_inst_n436,
         round_inst_S_10__sbox_inst_com_z_inst_n435,
         round_inst_S_10__sbox_inst_com_z_inst_n434,
         round_inst_S_10__sbox_inst_com_z_inst_n433,
         round_inst_S_10__sbox_inst_com_z_inst_n432,
         round_inst_S_10__sbox_inst_com_z_inst_n431,
         round_inst_S_10__sbox_inst_com_z_inst_n430,
         round_inst_S_10__sbox_inst_com_z_inst_n429,
         round_inst_S_10__sbox_inst_com_z_inst_n428,
         round_inst_S_10__sbox_inst_com_z_inst_n427,
         round_inst_S_10__sbox_inst_com_z_inst_n426,
         round_inst_S_10__sbox_inst_com_z_inst_n425,
         round_inst_S_10__sbox_inst_com_z_inst_n424,
         round_inst_S_10__sbox_inst_com_z_inst_n423,
         round_inst_S_10__sbox_inst_com_z_inst_n422,
         round_inst_S_10__sbox_inst_com_z_inst_n421,
         round_inst_S_10__sbox_inst_com_z_inst_n420,
         round_inst_S_10__sbox_inst_com_z_inst_n419,
         round_inst_S_10__sbox_inst_com_z_inst_n418,
         round_inst_S_10__sbox_inst_com_z_inst_n417,
         round_inst_S_10__sbox_inst_com_z_inst_n416,
         round_inst_S_10__sbox_inst_com_z_inst_n415,
         round_inst_S_10__sbox_inst_com_z_inst_n414,
         round_inst_S_10__sbox_inst_com_z_inst_n413,
         round_inst_S_10__sbox_inst_com_z_inst_n412,
         round_inst_S_10__sbox_inst_com_z_inst_n411,
         round_inst_S_10__sbox_inst_com_z_inst_n410,
         round_inst_S_10__sbox_inst_com_z_inst_n409,
         round_inst_S_10__sbox_inst_com_z_inst_n408,
         round_inst_S_10__sbox_inst_com_z_inst_n407,
         round_inst_S_10__sbox_inst_com_z_inst_n406,
         round_inst_S_10__sbox_inst_com_z_inst_n405,
         round_inst_S_10__sbox_inst_com_z_inst_n404,
         round_inst_S_10__sbox_inst_com_z_inst_n403,
         round_inst_S_10__sbox_inst_com_z_inst_n402,
         round_inst_S_10__sbox_inst_com_z_inst_n401,
         round_inst_S_10__sbox_inst_com_z_inst_n400,
         round_inst_S_10__sbox_inst_com_z_inst_n399,
         round_inst_S_10__sbox_inst_com_z_inst_n398,
         round_inst_S_10__sbox_inst_com_z_inst_n397,
         round_inst_S_10__sbox_inst_com_z_inst_n396,
         round_inst_S_10__sbox_inst_com_z_inst_n395,
         round_inst_S_10__sbox_inst_com_z_inst_n394,
         round_inst_S_10__sbox_inst_com_z_inst_n393,
         round_inst_S_10__sbox_inst_com_z_inst_n392,
         round_inst_S_10__sbox_inst_com_z_inst_n391,
         round_inst_S_11__sbox_inst_n6, round_inst_S_11__sbox_inst_n5,
         round_inst_S_11__sbox_inst_n4, round_inst_S_11__sbox_inst_n3,
         round_inst_S_11__sbox_inst_n2, round_inst_S_11__sbox_inst_n1,
         round_inst_S_11__sbox_inst_com_w_inst_n532,
         round_inst_S_11__sbox_inst_com_w_inst_n531,
         round_inst_S_11__sbox_inst_com_w_inst_n530,
         round_inst_S_11__sbox_inst_com_w_inst_n529,
         round_inst_S_11__sbox_inst_com_w_inst_n528,
         round_inst_S_11__sbox_inst_com_w_inst_n527,
         round_inst_S_11__sbox_inst_com_w_inst_n526,
         round_inst_S_11__sbox_inst_com_w_inst_n525,
         round_inst_S_11__sbox_inst_com_w_inst_n524,
         round_inst_S_11__sbox_inst_com_w_inst_n523,
         round_inst_S_11__sbox_inst_com_w_inst_n522,
         round_inst_S_11__sbox_inst_com_w_inst_n521,
         round_inst_S_11__sbox_inst_com_w_inst_n520,
         round_inst_S_11__sbox_inst_com_w_inst_n519,
         round_inst_S_11__sbox_inst_com_w_inst_n518,
         round_inst_S_11__sbox_inst_com_w_inst_n517,
         round_inst_S_11__sbox_inst_com_w_inst_n516,
         round_inst_S_11__sbox_inst_com_w_inst_n515,
         round_inst_S_11__sbox_inst_com_w_inst_n514,
         round_inst_S_11__sbox_inst_com_w_inst_n513,
         round_inst_S_11__sbox_inst_com_w_inst_n512,
         round_inst_S_11__sbox_inst_com_w_inst_n511,
         round_inst_S_11__sbox_inst_com_w_inst_n510,
         round_inst_S_11__sbox_inst_com_w_inst_n509,
         round_inst_S_11__sbox_inst_com_w_inst_n508,
         round_inst_S_11__sbox_inst_com_w_inst_n507,
         round_inst_S_11__sbox_inst_com_w_inst_n506,
         round_inst_S_11__sbox_inst_com_w_inst_n505,
         round_inst_S_11__sbox_inst_com_w_inst_n504,
         round_inst_S_11__sbox_inst_com_w_inst_n503,
         round_inst_S_11__sbox_inst_com_w_inst_n502,
         round_inst_S_11__sbox_inst_com_w_inst_n501,
         round_inst_S_11__sbox_inst_com_w_inst_n500,
         round_inst_S_11__sbox_inst_com_w_inst_n499,
         round_inst_S_11__sbox_inst_com_w_inst_n498,
         round_inst_S_11__sbox_inst_com_w_inst_n497,
         round_inst_S_11__sbox_inst_com_w_inst_n496,
         round_inst_S_11__sbox_inst_com_w_inst_n495,
         round_inst_S_11__sbox_inst_com_w_inst_n494,
         round_inst_S_11__sbox_inst_com_w_inst_n493,
         round_inst_S_11__sbox_inst_com_w_inst_n492,
         round_inst_S_11__sbox_inst_com_w_inst_n491,
         round_inst_S_11__sbox_inst_com_w_inst_n490,
         round_inst_S_11__sbox_inst_com_w_inst_n489,
         round_inst_S_11__sbox_inst_com_w_inst_n488,
         round_inst_S_11__sbox_inst_com_w_inst_n487,
         round_inst_S_11__sbox_inst_com_w_inst_n486,
         round_inst_S_11__sbox_inst_com_w_inst_n485,
         round_inst_S_11__sbox_inst_com_w_inst_n484,
         round_inst_S_11__sbox_inst_com_w_inst_n483,
         round_inst_S_11__sbox_inst_com_w_inst_n482,
         round_inst_S_11__sbox_inst_com_w_inst_n481,
         round_inst_S_11__sbox_inst_com_w_inst_n480,
         round_inst_S_11__sbox_inst_com_w_inst_n479,
         round_inst_S_11__sbox_inst_com_w_inst_n478,
         round_inst_S_11__sbox_inst_com_w_inst_n477,
         round_inst_S_11__sbox_inst_com_w_inst_n476,
         round_inst_S_11__sbox_inst_com_w_inst_n475,
         round_inst_S_11__sbox_inst_com_w_inst_n474,
         round_inst_S_11__sbox_inst_com_w_inst_n473,
         round_inst_S_11__sbox_inst_com_w_inst_n472,
         round_inst_S_11__sbox_inst_com_w_inst_n471,
         round_inst_S_11__sbox_inst_com_w_inst_n470,
         round_inst_S_11__sbox_inst_com_w_inst_n469,
         round_inst_S_11__sbox_inst_com_w_inst_n468,
         round_inst_S_11__sbox_inst_com_w_inst_n467,
         round_inst_S_11__sbox_inst_com_w_inst_n466,
         round_inst_S_11__sbox_inst_com_w_inst_n465,
         round_inst_S_11__sbox_inst_com_w_inst_n464,
         round_inst_S_11__sbox_inst_com_w_inst_n463,
         round_inst_S_11__sbox_inst_com_w_inst_n462,
         round_inst_S_11__sbox_inst_com_w_inst_n461,
         round_inst_S_11__sbox_inst_com_w_inst_n460,
         round_inst_S_11__sbox_inst_com_w_inst_n459,
         round_inst_S_11__sbox_inst_com_w_inst_n458,
         round_inst_S_11__sbox_inst_com_w_inst_n457,
         round_inst_S_11__sbox_inst_com_w_inst_n456,
         round_inst_S_11__sbox_inst_com_w_inst_n455,
         round_inst_S_11__sbox_inst_com_w_inst_n454,
         round_inst_S_11__sbox_inst_com_w_inst_n453,
         round_inst_S_11__sbox_inst_com_w_inst_n452,
         round_inst_S_11__sbox_inst_com_w_inst_n451,
         round_inst_S_11__sbox_inst_com_w_inst_n450,
         round_inst_S_11__sbox_inst_com_w_inst_n449,
         round_inst_S_11__sbox_inst_com_w_inst_n448,
         round_inst_S_11__sbox_inst_com_w_inst_n447,
         round_inst_S_11__sbox_inst_com_w_inst_n446,
         round_inst_S_11__sbox_inst_com_w_inst_n445,
         round_inst_S_11__sbox_inst_com_w_inst_n444,
         round_inst_S_11__sbox_inst_com_w_inst_n443,
         round_inst_S_11__sbox_inst_com_w_inst_n442,
         round_inst_S_11__sbox_inst_com_w_inst_n441,
         round_inst_S_11__sbox_inst_com_w_inst_n440,
         round_inst_S_11__sbox_inst_com_w_inst_n439,
         round_inst_S_11__sbox_inst_com_w_inst_n438,
         round_inst_S_11__sbox_inst_com_w_inst_n437,
         round_inst_S_11__sbox_inst_com_w_inst_n436,
         round_inst_S_11__sbox_inst_com_w_inst_n435,
         round_inst_S_11__sbox_inst_com_w_inst_n434,
         round_inst_S_11__sbox_inst_com_w_inst_n433,
         round_inst_S_11__sbox_inst_com_w_inst_n432,
         round_inst_S_11__sbox_inst_com_w_inst_n431,
         round_inst_S_11__sbox_inst_com_w_inst_n430,
         round_inst_S_11__sbox_inst_com_w_inst_n429,
         round_inst_S_11__sbox_inst_com_w_inst_n428,
         round_inst_S_11__sbox_inst_com_w_inst_n427,
         round_inst_S_11__sbox_inst_com_w_inst_n426,
         round_inst_S_11__sbox_inst_com_w_inst_n425,
         round_inst_S_11__sbox_inst_com_w_inst_n424,
         round_inst_S_11__sbox_inst_com_w_inst_n423,
         round_inst_S_11__sbox_inst_com_w_inst_n422,
         round_inst_S_11__sbox_inst_com_w_inst_n421,
         round_inst_S_11__sbox_inst_com_w_inst_n420,
         round_inst_S_11__sbox_inst_com_w_inst_n419,
         round_inst_S_11__sbox_inst_com_w_inst_n418,
         round_inst_S_11__sbox_inst_com_w_inst_n417,
         round_inst_S_11__sbox_inst_com_w_inst_n416,
         round_inst_S_11__sbox_inst_com_w_inst_n415,
         round_inst_S_11__sbox_inst_com_w_inst_n414,
         round_inst_S_11__sbox_inst_com_w_inst_n413,
         round_inst_S_11__sbox_inst_com_w_inst_n412,
         round_inst_S_11__sbox_inst_com_w_inst_n411,
         round_inst_S_11__sbox_inst_com_w_inst_n410,
         round_inst_S_11__sbox_inst_com_w_inst_n409,
         round_inst_S_11__sbox_inst_com_w_inst_n408,
         round_inst_S_11__sbox_inst_com_w_inst_n407,
         round_inst_S_11__sbox_inst_com_w_inst_n406,
         round_inst_S_11__sbox_inst_com_w_inst_n405,
         round_inst_S_11__sbox_inst_com_w_inst_n404,
         round_inst_S_11__sbox_inst_com_w_inst_n403,
         round_inst_S_11__sbox_inst_com_w_inst_n402,
         round_inst_S_11__sbox_inst_com_w_inst_n401,
         round_inst_S_11__sbox_inst_com_w_inst_n400,
         round_inst_S_11__sbox_inst_com_w_inst_n399,
         round_inst_S_11__sbox_inst_com_w_inst_n398,
         round_inst_S_11__sbox_inst_com_w_inst_n397,
         round_inst_S_11__sbox_inst_com_w_inst_n396,
         round_inst_S_11__sbox_inst_com_x_inst_n519,
         round_inst_S_11__sbox_inst_com_x_inst_n518,
         round_inst_S_11__sbox_inst_com_x_inst_n517,
         round_inst_S_11__sbox_inst_com_x_inst_n516,
         round_inst_S_11__sbox_inst_com_x_inst_n515,
         round_inst_S_11__sbox_inst_com_x_inst_n514,
         round_inst_S_11__sbox_inst_com_x_inst_n513,
         round_inst_S_11__sbox_inst_com_x_inst_n512,
         round_inst_S_11__sbox_inst_com_x_inst_n511,
         round_inst_S_11__sbox_inst_com_x_inst_n510,
         round_inst_S_11__sbox_inst_com_x_inst_n509,
         round_inst_S_11__sbox_inst_com_x_inst_n508,
         round_inst_S_11__sbox_inst_com_x_inst_n507,
         round_inst_S_11__sbox_inst_com_x_inst_n506,
         round_inst_S_11__sbox_inst_com_x_inst_n505,
         round_inst_S_11__sbox_inst_com_x_inst_n504,
         round_inst_S_11__sbox_inst_com_x_inst_n503,
         round_inst_S_11__sbox_inst_com_x_inst_n502,
         round_inst_S_11__sbox_inst_com_x_inst_n501,
         round_inst_S_11__sbox_inst_com_x_inst_n500,
         round_inst_S_11__sbox_inst_com_x_inst_n499,
         round_inst_S_11__sbox_inst_com_x_inst_n498,
         round_inst_S_11__sbox_inst_com_x_inst_n497,
         round_inst_S_11__sbox_inst_com_x_inst_n496,
         round_inst_S_11__sbox_inst_com_x_inst_n495,
         round_inst_S_11__sbox_inst_com_x_inst_n494,
         round_inst_S_11__sbox_inst_com_x_inst_n493,
         round_inst_S_11__sbox_inst_com_x_inst_n492,
         round_inst_S_11__sbox_inst_com_x_inst_n491,
         round_inst_S_11__sbox_inst_com_x_inst_n490,
         round_inst_S_11__sbox_inst_com_x_inst_n489,
         round_inst_S_11__sbox_inst_com_x_inst_n488,
         round_inst_S_11__sbox_inst_com_x_inst_n487,
         round_inst_S_11__sbox_inst_com_x_inst_n486,
         round_inst_S_11__sbox_inst_com_x_inst_n485,
         round_inst_S_11__sbox_inst_com_x_inst_n484,
         round_inst_S_11__sbox_inst_com_x_inst_n483,
         round_inst_S_11__sbox_inst_com_x_inst_n482,
         round_inst_S_11__sbox_inst_com_x_inst_n481,
         round_inst_S_11__sbox_inst_com_x_inst_n480,
         round_inst_S_11__sbox_inst_com_x_inst_n479,
         round_inst_S_11__sbox_inst_com_x_inst_n478,
         round_inst_S_11__sbox_inst_com_x_inst_n477,
         round_inst_S_11__sbox_inst_com_x_inst_n476,
         round_inst_S_11__sbox_inst_com_x_inst_n475,
         round_inst_S_11__sbox_inst_com_x_inst_n474,
         round_inst_S_11__sbox_inst_com_x_inst_n473,
         round_inst_S_11__sbox_inst_com_x_inst_n472,
         round_inst_S_11__sbox_inst_com_x_inst_n471,
         round_inst_S_11__sbox_inst_com_x_inst_n470,
         round_inst_S_11__sbox_inst_com_x_inst_n469,
         round_inst_S_11__sbox_inst_com_x_inst_n468,
         round_inst_S_11__sbox_inst_com_x_inst_n467,
         round_inst_S_11__sbox_inst_com_x_inst_n466,
         round_inst_S_11__sbox_inst_com_x_inst_n465,
         round_inst_S_11__sbox_inst_com_x_inst_n464,
         round_inst_S_11__sbox_inst_com_x_inst_n463,
         round_inst_S_11__sbox_inst_com_x_inst_n462,
         round_inst_S_11__sbox_inst_com_x_inst_n461,
         round_inst_S_11__sbox_inst_com_x_inst_n460,
         round_inst_S_11__sbox_inst_com_x_inst_n459,
         round_inst_S_11__sbox_inst_com_x_inst_n458,
         round_inst_S_11__sbox_inst_com_x_inst_n457,
         round_inst_S_11__sbox_inst_com_x_inst_n456,
         round_inst_S_11__sbox_inst_com_x_inst_n455,
         round_inst_S_11__sbox_inst_com_x_inst_n454,
         round_inst_S_11__sbox_inst_com_x_inst_n453,
         round_inst_S_11__sbox_inst_com_x_inst_n452,
         round_inst_S_11__sbox_inst_com_x_inst_n451,
         round_inst_S_11__sbox_inst_com_x_inst_n450,
         round_inst_S_11__sbox_inst_com_x_inst_n449,
         round_inst_S_11__sbox_inst_com_x_inst_n448,
         round_inst_S_11__sbox_inst_com_x_inst_n447,
         round_inst_S_11__sbox_inst_com_x_inst_n446,
         round_inst_S_11__sbox_inst_com_x_inst_n445,
         round_inst_S_11__sbox_inst_com_x_inst_n444,
         round_inst_S_11__sbox_inst_com_x_inst_n443,
         round_inst_S_11__sbox_inst_com_x_inst_n442,
         round_inst_S_11__sbox_inst_com_x_inst_n441,
         round_inst_S_11__sbox_inst_com_x_inst_n440,
         round_inst_S_11__sbox_inst_com_x_inst_n439,
         round_inst_S_11__sbox_inst_com_x_inst_n438,
         round_inst_S_11__sbox_inst_com_x_inst_n437,
         round_inst_S_11__sbox_inst_com_x_inst_n436,
         round_inst_S_11__sbox_inst_com_x_inst_n435,
         round_inst_S_11__sbox_inst_com_x_inst_n434,
         round_inst_S_11__sbox_inst_com_x_inst_n433,
         round_inst_S_11__sbox_inst_com_x_inst_n432,
         round_inst_S_11__sbox_inst_com_x_inst_n431,
         round_inst_S_11__sbox_inst_com_x_inst_n430,
         round_inst_S_11__sbox_inst_com_x_inst_n429,
         round_inst_S_11__sbox_inst_com_x_inst_n428,
         round_inst_S_11__sbox_inst_com_x_inst_n427,
         round_inst_S_11__sbox_inst_com_x_inst_n426,
         round_inst_S_11__sbox_inst_com_x_inst_n425,
         round_inst_S_11__sbox_inst_com_x_inst_n424,
         round_inst_S_11__sbox_inst_com_x_inst_n423,
         round_inst_S_11__sbox_inst_com_x_inst_n422,
         round_inst_S_11__sbox_inst_com_x_inst_n421,
         round_inst_S_11__sbox_inst_com_x_inst_n420,
         round_inst_S_11__sbox_inst_com_x_inst_n419,
         round_inst_S_11__sbox_inst_com_x_inst_n418,
         round_inst_S_11__sbox_inst_com_x_inst_n417,
         round_inst_S_11__sbox_inst_com_x_inst_n416,
         round_inst_S_11__sbox_inst_com_x_inst_n415,
         round_inst_S_11__sbox_inst_com_x_inst_n414,
         round_inst_S_11__sbox_inst_com_x_inst_n413,
         round_inst_S_11__sbox_inst_com_x_inst_n412,
         round_inst_S_11__sbox_inst_com_x_inst_n411,
         round_inst_S_11__sbox_inst_com_x_inst_n410,
         round_inst_S_11__sbox_inst_com_x_inst_n409,
         round_inst_S_11__sbox_inst_com_x_inst_n408,
         round_inst_S_11__sbox_inst_com_x_inst_n407,
         round_inst_S_11__sbox_inst_com_x_inst_n406,
         round_inst_S_11__sbox_inst_com_x_inst_n405,
         round_inst_S_11__sbox_inst_com_x_inst_n404,
         round_inst_S_11__sbox_inst_com_x_inst_n403,
         round_inst_S_11__sbox_inst_com_x_inst_n402,
         round_inst_S_11__sbox_inst_com_x_inst_n401,
         round_inst_S_11__sbox_inst_com_x_inst_n400,
         round_inst_S_11__sbox_inst_com_x_inst_n399,
         round_inst_S_11__sbox_inst_com_x_inst_n398,
         round_inst_S_11__sbox_inst_com_x_inst_n397,
         round_inst_S_11__sbox_inst_com_x_inst_n396,
         round_inst_S_11__sbox_inst_com_x_inst_n395,
         round_inst_S_11__sbox_inst_com_x_inst_n394,
         round_inst_S_11__sbox_inst_com_x_inst_n393,
         round_inst_S_11__sbox_inst_com_x_inst_n392,
         round_inst_S_11__sbox_inst_com_x_inst_n391,
         round_inst_S_11__sbox_inst_com_x_inst_n390,
         round_inst_S_11__sbox_inst_com_x_inst_n389,
         round_inst_S_11__sbox_inst_com_x_inst_n388,
         round_inst_S_11__sbox_inst_com_x_inst_n387,
         round_inst_S_11__sbox_inst_com_x_inst_n386,
         round_inst_S_11__sbox_inst_com_x_inst_n385,
         round_inst_S_11__sbox_inst_com_x_inst_n384,
         round_inst_S_11__sbox_inst_com_x_inst_n383,
         round_inst_S_11__sbox_inst_com_x_inst_n382,
         round_inst_S_11__sbox_inst_com_x_inst_n381,
         round_inst_S_11__sbox_inst_com_x_inst_n380,
         round_inst_S_11__sbox_inst_com_y_inst_n517,
         round_inst_S_11__sbox_inst_com_y_inst_n516,
         round_inst_S_11__sbox_inst_com_y_inst_n515,
         round_inst_S_11__sbox_inst_com_y_inst_n514,
         round_inst_S_11__sbox_inst_com_y_inst_n513,
         round_inst_S_11__sbox_inst_com_y_inst_n512,
         round_inst_S_11__sbox_inst_com_y_inst_n511,
         round_inst_S_11__sbox_inst_com_y_inst_n510,
         round_inst_S_11__sbox_inst_com_y_inst_n509,
         round_inst_S_11__sbox_inst_com_y_inst_n508,
         round_inst_S_11__sbox_inst_com_y_inst_n507,
         round_inst_S_11__sbox_inst_com_y_inst_n506,
         round_inst_S_11__sbox_inst_com_y_inst_n505,
         round_inst_S_11__sbox_inst_com_y_inst_n504,
         round_inst_S_11__sbox_inst_com_y_inst_n503,
         round_inst_S_11__sbox_inst_com_y_inst_n502,
         round_inst_S_11__sbox_inst_com_y_inst_n501,
         round_inst_S_11__sbox_inst_com_y_inst_n500,
         round_inst_S_11__sbox_inst_com_y_inst_n499,
         round_inst_S_11__sbox_inst_com_y_inst_n498,
         round_inst_S_11__sbox_inst_com_y_inst_n497,
         round_inst_S_11__sbox_inst_com_y_inst_n496,
         round_inst_S_11__sbox_inst_com_y_inst_n495,
         round_inst_S_11__sbox_inst_com_y_inst_n494,
         round_inst_S_11__sbox_inst_com_y_inst_n493,
         round_inst_S_11__sbox_inst_com_y_inst_n492,
         round_inst_S_11__sbox_inst_com_y_inst_n491,
         round_inst_S_11__sbox_inst_com_y_inst_n490,
         round_inst_S_11__sbox_inst_com_y_inst_n489,
         round_inst_S_11__sbox_inst_com_y_inst_n488,
         round_inst_S_11__sbox_inst_com_y_inst_n487,
         round_inst_S_11__sbox_inst_com_y_inst_n486,
         round_inst_S_11__sbox_inst_com_y_inst_n485,
         round_inst_S_11__sbox_inst_com_y_inst_n484,
         round_inst_S_11__sbox_inst_com_y_inst_n483,
         round_inst_S_11__sbox_inst_com_y_inst_n482,
         round_inst_S_11__sbox_inst_com_y_inst_n481,
         round_inst_S_11__sbox_inst_com_y_inst_n480,
         round_inst_S_11__sbox_inst_com_y_inst_n479,
         round_inst_S_11__sbox_inst_com_y_inst_n478,
         round_inst_S_11__sbox_inst_com_y_inst_n477,
         round_inst_S_11__sbox_inst_com_y_inst_n476,
         round_inst_S_11__sbox_inst_com_y_inst_n475,
         round_inst_S_11__sbox_inst_com_y_inst_n474,
         round_inst_S_11__sbox_inst_com_y_inst_n473,
         round_inst_S_11__sbox_inst_com_y_inst_n472,
         round_inst_S_11__sbox_inst_com_y_inst_n471,
         round_inst_S_11__sbox_inst_com_y_inst_n470,
         round_inst_S_11__sbox_inst_com_y_inst_n469,
         round_inst_S_11__sbox_inst_com_y_inst_n468,
         round_inst_S_11__sbox_inst_com_y_inst_n467,
         round_inst_S_11__sbox_inst_com_y_inst_n466,
         round_inst_S_11__sbox_inst_com_y_inst_n465,
         round_inst_S_11__sbox_inst_com_y_inst_n464,
         round_inst_S_11__sbox_inst_com_y_inst_n463,
         round_inst_S_11__sbox_inst_com_y_inst_n462,
         round_inst_S_11__sbox_inst_com_y_inst_n461,
         round_inst_S_11__sbox_inst_com_y_inst_n460,
         round_inst_S_11__sbox_inst_com_y_inst_n459,
         round_inst_S_11__sbox_inst_com_y_inst_n458,
         round_inst_S_11__sbox_inst_com_y_inst_n457,
         round_inst_S_11__sbox_inst_com_y_inst_n456,
         round_inst_S_11__sbox_inst_com_y_inst_n455,
         round_inst_S_11__sbox_inst_com_y_inst_n454,
         round_inst_S_11__sbox_inst_com_y_inst_n453,
         round_inst_S_11__sbox_inst_com_y_inst_n452,
         round_inst_S_11__sbox_inst_com_y_inst_n451,
         round_inst_S_11__sbox_inst_com_y_inst_n450,
         round_inst_S_11__sbox_inst_com_y_inst_n449,
         round_inst_S_11__sbox_inst_com_y_inst_n448,
         round_inst_S_11__sbox_inst_com_y_inst_n447,
         round_inst_S_11__sbox_inst_com_y_inst_n446,
         round_inst_S_11__sbox_inst_com_y_inst_n445,
         round_inst_S_11__sbox_inst_com_y_inst_n444,
         round_inst_S_11__sbox_inst_com_y_inst_n443,
         round_inst_S_11__sbox_inst_com_y_inst_n442,
         round_inst_S_11__sbox_inst_com_y_inst_n441,
         round_inst_S_11__sbox_inst_com_y_inst_n440,
         round_inst_S_11__sbox_inst_com_y_inst_n439,
         round_inst_S_11__sbox_inst_com_y_inst_n438,
         round_inst_S_11__sbox_inst_com_y_inst_n437,
         round_inst_S_11__sbox_inst_com_y_inst_n436,
         round_inst_S_11__sbox_inst_com_y_inst_n435,
         round_inst_S_11__sbox_inst_com_y_inst_n434,
         round_inst_S_11__sbox_inst_com_y_inst_n433,
         round_inst_S_11__sbox_inst_com_y_inst_n432,
         round_inst_S_11__sbox_inst_com_y_inst_n431,
         round_inst_S_11__sbox_inst_com_y_inst_n430,
         round_inst_S_11__sbox_inst_com_y_inst_n429,
         round_inst_S_11__sbox_inst_com_y_inst_n428,
         round_inst_S_11__sbox_inst_com_y_inst_n427,
         round_inst_S_11__sbox_inst_com_y_inst_n426,
         round_inst_S_11__sbox_inst_com_y_inst_n425,
         round_inst_S_11__sbox_inst_com_y_inst_n424,
         round_inst_S_11__sbox_inst_com_y_inst_n423,
         round_inst_S_11__sbox_inst_com_y_inst_n422,
         round_inst_S_11__sbox_inst_com_y_inst_n421,
         round_inst_S_11__sbox_inst_com_y_inst_n420,
         round_inst_S_11__sbox_inst_com_y_inst_n419,
         round_inst_S_11__sbox_inst_com_y_inst_n418,
         round_inst_S_11__sbox_inst_com_y_inst_n417,
         round_inst_S_11__sbox_inst_com_y_inst_n416,
         round_inst_S_11__sbox_inst_com_y_inst_n415,
         round_inst_S_11__sbox_inst_com_y_inst_n414,
         round_inst_S_11__sbox_inst_com_y_inst_n413,
         round_inst_S_11__sbox_inst_com_y_inst_n412,
         round_inst_S_11__sbox_inst_com_y_inst_n411,
         round_inst_S_11__sbox_inst_com_y_inst_n410,
         round_inst_S_11__sbox_inst_com_y_inst_n409,
         round_inst_S_11__sbox_inst_com_y_inst_n408,
         round_inst_S_11__sbox_inst_com_y_inst_n407,
         round_inst_S_11__sbox_inst_com_y_inst_n406,
         round_inst_S_11__sbox_inst_com_y_inst_n405,
         round_inst_S_11__sbox_inst_com_y_inst_n404,
         round_inst_S_11__sbox_inst_com_y_inst_n403,
         round_inst_S_11__sbox_inst_com_y_inst_n402,
         round_inst_S_11__sbox_inst_com_y_inst_n401,
         round_inst_S_11__sbox_inst_com_y_inst_n400,
         round_inst_S_11__sbox_inst_com_y_inst_n399,
         round_inst_S_11__sbox_inst_com_y_inst_n398,
         round_inst_S_11__sbox_inst_com_y_inst_n397,
         round_inst_S_11__sbox_inst_com_y_inst_n396,
         round_inst_S_11__sbox_inst_com_y_inst_n395,
         round_inst_S_11__sbox_inst_com_y_inst_n394,
         round_inst_S_11__sbox_inst_com_y_inst_n393,
         round_inst_S_11__sbox_inst_com_y_inst_n392,
         round_inst_S_11__sbox_inst_com_y_inst_n391,
         round_inst_S_11__sbox_inst_com_y_inst_n390,
         round_inst_S_11__sbox_inst_com_y_inst_n389,
         round_inst_S_11__sbox_inst_com_y_inst_n388,
         round_inst_S_11__sbox_inst_com_y_inst_n387,
         round_inst_S_11__sbox_inst_com_y_inst_n386,
         round_inst_S_11__sbox_inst_com_z_inst_n523,
         round_inst_S_11__sbox_inst_com_z_inst_n522,
         round_inst_S_11__sbox_inst_com_z_inst_n521,
         round_inst_S_11__sbox_inst_com_z_inst_n520,
         round_inst_S_11__sbox_inst_com_z_inst_n519,
         round_inst_S_11__sbox_inst_com_z_inst_n518,
         round_inst_S_11__sbox_inst_com_z_inst_n517,
         round_inst_S_11__sbox_inst_com_z_inst_n516,
         round_inst_S_11__sbox_inst_com_z_inst_n515,
         round_inst_S_11__sbox_inst_com_z_inst_n514,
         round_inst_S_11__sbox_inst_com_z_inst_n513,
         round_inst_S_11__sbox_inst_com_z_inst_n512,
         round_inst_S_11__sbox_inst_com_z_inst_n511,
         round_inst_S_11__sbox_inst_com_z_inst_n510,
         round_inst_S_11__sbox_inst_com_z_inst_n509,
         round_inst_S_11__sbox_inst_com_z_inst_n508,
         round_inst_S_11__sbox_inst_com_z_inst_n507,
         round_inst_S_11__sbox_inst_com_z_inst_n506,
         round_inst_S_11__sbox_inst_com_z_inst_n505,
         round_inst_S_11__sbox_inst_com_z_inst_n504,
         round_inst_S_11__sbox_inst_com_z_inst_n503,
         round_inst_S_11__sbox_inst_com_z_inst_n502,
         round_inst_S_11__sbox_inst_com_z_inst_n501,
         round_inst_S_11__sbox_inst_com_z_inst_n500,
         round_inst_S_11__sbox_inst_com_z_inst_n499,
         round_inst_S_11__sbox_inst_com_z_inst_n498,
         round_inst_S_11__sbox_inst_com_z_inst_n497,
         round_inst_S_11__sbox_inst_com_z_inst_n496,
         round_inst_S_11__sbox_inst_com_z_inst_n495,
         round_inst_S_11__sbox_inst_com_z_inst_n494,
         round_inst_S_11__sbox_inst_com_z_inst_n493,
         round_inst_S_11__sbox_inst_com_z_inst_n492,
         round_inst_S_11__sbox_inst_com_z_inst_n491,
         round_inst_S_11__sbox_inst_com_z_inst_n490,
         round_inst_S_11__sbox_inst_com_z_inst_n489,
         round_inst_S_11__sbox_inst_com_z_inst_n488,
         round_inst_S_11__sbox_inst_com_z_inst_n487,
         round_inst_S_11__sbox_inst_com_z_inst_n486,
         round_inst_S_11__sbox_inst_com_z_inst_n485,
         round_inst_S_11__sbox_inst_com_z_inst_n484,
         round_inst_S_11__sbox_inst_com_z_inst_n483,
         round_inst_S_11__sbox_inst_com_z_inst_n482,
         round_inst_S_11__sbox_inst_com_z_inst_n481,
         round_inst_S_11__sbox_inst_com_z_inst_n480,
         round_inst_S_11__sbox_inst_com_z_inst_n479,
         round_inst_S_11__sbox_inst_com_z_inst_n478,
         round_inst_S_11__sbox_inst_com_z_inst_n477,
         round_inst_S_11__sbox_inst_com_z_inst_n476,
         round_inst_S_11__sbox_inst_com_z_inst_n475,
         round_inst_S_11__sbox_inst_com_z_inst_n474,
         round_inst_S_11__sbox_inst_com_z_inst_n473,
         round_inst_S_11__sbox_inst_com_z_inst_n472,
         round_inst_S_11__sbox_inst_com_z_inst_n471,
         round_inst_S_11__sbox_inst_com_z_inst_n470,
         round_inst_S_11__sbox_inst_com_z_inst_n469,
         round_inst_S_11__sbox_inst_com_z_inst_n468,
         round_inst_S_11__sbox_inst_com_z_inst_n467,
         round_inst_S_11__sbox_inst_com_z_inst_n466,
         round_inst_S_11__sbox_inst_com_z_inst_n465,
         round_inst_S_11__sbox_inst_com_z_inst_n464,
         round_inst_S_11__sbox_inst_com_z_inst_n463,
         round_inst_S_11__sbox_inst_com_z_inst_n462,
         round_inst_S_11__sbox_inst_com_z_inst_n461,
         round_inst_S_11__sbox_inst_com_z_inst_n460,
         round_inst_S_11__sbox_inst_com_z_inst_n459,
         round_inst_S_11__sbox_inst_com_z_inst_n458,
         round_inst_S_11__sbox_inst_com_z_inst_n457,
         round_inst_S_11__sbox_inst_com_z_inst_n456,
         round_inst_S_11__sbox_inst_com_z_inst_n455,
         round_inst_S_11__sbox_inst_com_z_inst_n454,
         round_inst_S_11__sbox_inst_com_z_inst_n453,
         round_inst_S_11__sbox_inst_com_z_inst_n452,
         round_inst_S_11__sbox_inst_com_z_inst_n451,
         round_inst_S_11__sbox_inst_com_z_inst_n450,
         round_inst_S_11__sbox_inst_com_z_inst_n449,
         round_inst_S_11__sbox_inst_com_z_inst_n448,
         round_inst_S_11__sbox_inst_com_z_inst_n447,
         round_inst_S_11__sbox_inst_com_z_inst_n446,
         round_inst_S_11__sbox_inst_com_z_inst_n445,
         round_inst_S_11__sbox_inst_com_z_inst_n444,
         round_inst_S_11__sbox_inst_com_z_inst_n443,
         round_inst_S_11__sbox_inst_com_z_inst_n442,
         round_inst_S_11__sbox_inst_com_z_inst_n441,
         round_inst_S_11__sbox_inst_com_z_inst_n440,
         round_inst_S_11__sbox_inst_com_z_inst_n439,
         round_inst_S_11__sbox_inst_com_z_inst_n438,
         round_inst_S_11__sbox_inst_com_z_inst_n437,
         round_inst_S_11__sbox_inst_com_z_inst_n436,
         round_inst_S_11__sbox_inst_com_z_inst_n435,
         round_inst_S_11__sbox_inst_com_z_inst_n434,
         round_inst_S_11__sbox_inst_com_z_inst_n433,
         round_inst_S_11__sbox_inst_com_z_inst_n432,
         round_inst_S_11__sbox_inst_com_z_inst_n431,
         round_inst_S_11__sbox_inst_com_z_inst_n430,
         round_inst_S_11__sbox_inst_com_z_inst_n429,
         round_inst_S_11__sbox_inst_com_z_inst_n428,
         round_inst_S_11__sbox_inst_com_z_inst_n427,
         round_inst_S_11__sbox_inst_com_z_inst_n426,
         round_inst_S_11__sbox_inst_com_z_inst_n425,
         round_inst_S_11__sbox_inst_com_z_inst_n424,
         round_inst_S_11__sbox_inst_com_z_inst_n423,
         round_inst_S_11__sbox_inst_com_z_inst_n422,
         round_inst_S_11__sbox_inst_com_z_inst_n421,
         round_inst_S_11__sbox_inst_com_z_inst_n420,
         round_inst_S_11__sbox_inst_com_z_inst_n419,
         round_inst_S_11__sbox_inst_com_z_inst_n418,
         round_inst_S_11__sbox_inst_com_z_inst_n417,
         round_inst_S_11__sbox_inst_com_z_inst_n416,
         round_inst_S_11__sbox_inst_com_z_inst_n415,
         round_inst_S_11__sbox_inst_com_z_inst_n414,
         round_inst_S_11__sbox_inst_com_z_inst_n413,
         round_inst_S_11__sbox_inst_com_z_inst_n412,
         round_inst_S_11__sbox_inst_com_z_inst_n411,
         round_inst_S_11__sbox_inst_com_z_inst_n410,
         round_inst_S_11__sbox_inst_com_z_inst_n409,
         round_inst_S_11__sbox_inst_com_z_inst_n408,
         round_inst_S_11__sbox_inst_com_z_inst_n407,
         round_inst_S_11__sbox_inst_com_z_inst_n406,
         round_inst_S_11__sbox_inst_com_z_inst_n405,
         round_inst_S_11__sbox_inst_com_z_inst_n404,
         round_inst_S_11__sbox_inst_com_z_inst_n403,
         round_inst_S_11__sbox_inst_com_z_inst_n402,
         round_inst_S_11__sbox_inst_com_z_inst_n401,
         round_inst_S_11__sbox_inst_com_z_inst_n400,
         round_inst_S_11__sbox_inst_com_z_inst_n399,
         round_inst_S_11__sbox_inst_com_z_inst_n398,
         round_inst_S_11__sbox_inst_com_z_inst_n397,
         round_inst_S_11__sbox_inst_com_z_inst_n396,
         round_inst_S_11__sbox_inst_com_z_inst_n395,
         round_inst_S_11__sbox_inst_com_z_inst_n394,
         round_inst_S_11__sbox_inst_com_z_inst_n393,
         round_inst_S_11__sbox_inst_com_z_inst_n392,
         round_inst_S_11__sbox_inst_com_z_inst_n391,
         round_inst_S_12__sbox_inst_n6, round_inst_S_12__sbox_inst_n5,
         round_inst_S_12__sbox_inst_n4, round_inst_S_12__sbox_inst_n3,
         round_inst_S_12__sbox_inst_n2, round_inst_S_12__sbox_inst_n1,
         round_inst_S_12__sbox_inst_com_w_inst_n529,
         round_inst_S_12__sbox_inst_com_w_inst_n528,
         round_inst_S_12__sbox_inst_com_w_inst_n527,
         round_inst_S_12__sbox_inst_com_w_inst_n526,
         round_inst_S_12__sbox_inst_com_w_inst_n525,
         round_inst_S_12__sbox_inst_com_w_inst_n524,
         round_inst_S_12__sbox_inst_com_w_inst_n523,
         round_inst_S_12__sbox_inst_com_w_inst_n522,
         round_inst_S_12__sbox_inst_com_w_inst_n521,
         round_inst_S_12__sbox_inst_com_w_inst_n520,
         round_inst_S_12__sbox_inst_com_w_inst_n519,
         round_inst_S_12__sbox_inst_com_w_inst_n518,
         round_inst_S_12__sbox_inst_com_w_inst_n517,
         round_inst_S_12__sbox_inst_com_w_inst_n516,
         round_inst_S_12__sbox_inst_com_w_inst_n515,
         round_inst_S_12__sbox_inst_com_w_inst_n514,
         round_inst_S_12__sbox_inst_com_w_inst_n513,
         round_inst_S_12__sbox_inst_com_w_inst_n512,
         round_inst_S_12__sbox_inst_com_w_inst_n511,
         round_inst_S_12__sbox_inst_com_w_inst_n510,
         round_inst_S_12__sbox_inst_com_w_inst_n509,
         round_inst_S_12__sbox_inst_com_w_inst_n508,
         round_inst_S_12__sbox_inst_com_w_inst_n507,
         round_inst_S_12__sbox_inst_com_w_inst_n506,
         round_inst_S_12__sbox_inst_com_w_inst_n505,
         round_inst_S_12__sbox_inst_com_w_inst_n504,
         round_inst_S_12__sbox_inst_com_w_inst_n503,
         round_inst_S_12__sbox_inst_com_w_inst_n502,
         round_inst_S_12__sbox_inst_com_w_inst_n501,
         round_inst_S_12__sbox_inst_com_w_inst_n500,
         round_inst_S_12__sbox_inst_com_w_inst_n499,
         round_inst_S_12__sbox_inst_com_w_inst_n498,
         round_inst_S_12__sbox_inst_com_w_inst_n497,
         round_inst_S_12__sbox_inst_com_w_inst_n496,
         round_inst_S_12__sbox_inst_com_w_inst_n495,
         round_inst_S_12__sbox_inst_com_w_inst_n494,
         round_inst_S_12__sbox_inst_com_w_inst_n493,
         round_inst_S_12__sbox_inst_com_w_inst_n492,
         round_inst_S_12__sbox_inst_com_w_inst_n491,
         round_inst_S_12__sbox_inst_com_w_inst_n490,
         round_inst_S_12__sbox_inst_com_w_inst_n489,
         round_inst_S_12__sbox_inst_com_w_inst_n488,
         round_inst_S_12__sbox_inst_com_w_inst_n487,
         round_inst_S_12__sbox_inst_com_w_inst_n486,
         round_inst_S_12__sbox_inst_com_w_inst_n485,
         round_inst_S_12__sbox_inst_com_w_inst_n484,
         round_inst_S_12__sbox_inst_com_w_inst_n483,
         round_inst_S_12__sbox_inst_com_w_inst_n482,
         round_inst_S_12__sbox_inst_com_w_inst_n481,
         round_inst_S_12__sbox_inst_com_w_inst_n480,
         round_inst_S_12__sbox_inst_com_w_inst_n479,
         round_inst_S_12__sbox_inst_com_w_inst_n478,
         round_inst_S_12__sbox_inst_com_w_inst_n477,
         round_inst_S_12__sbox_inst_com_w_inst_n476,
         round_inst_S_12__sbox_inst_com_w_inst_n475,
         round_inst_S_12__sbox_inst_com_w_inst_n474,
         round_inst_S_12__sbox_inst_com_w_inst_n473,
         round_inst_S_12__sbox_inst_com_w_inst_n472,
         round_inst_S_12__sbox_inst_com_w_inst_n471,
         round_inst_S_12__sbox_inst_com_w_inst_n470,
         round_inst_S_12__sbox_inst_com_w_inst_n469,
         round_inst_S_12__sbox_inst_com_w_inst_n468,
         round_inst_S_12__sbox_inst_com_w_inst_n467,
         round_inst_S_12__sbox_inst_com_w_inst_n466,
         round_inst_S_12__sbox_inst_com_w_inst_n465,
         round_inst_S_12__sbox_inst_com_w_inst_n464,
         round_inst_S_12__sbox_inst_com_w_inst_n463,
         round_inst_S_12__sbox_inst_com_w_inst_n462,
         round_inst_S_12__sbox_inst_com_w_inst_n461,
         round_inst_S_12__sbox_inst_com_w_inst_n460,
         round_inst_S_12__sbox_inst_com_w_inst_n459,
         round_inst_S_12__sbox_inst_com_w_inst_n458,
         round_inst_S_12__sbox_inst_com_w_inst_n457,
         round_inst_S_12__sbox_inst_com_w_inst_n456,
         round_inst_S_12__sbox_inst_com_w_inst_n455,
         round_inst_S_12__sbox_inst_com_w_inst_n454,
         round_inst_S_12__sbox_inst_com_w_inst_n453,
         round_inst_S_12__sbox_inst_com_w_inst_n452,
         round_inst_S_12__sbox_inst_com_w_inst_n451,
         round_inst_S_12__sbox_inst_com_w_inst_n450,
         round_inst_S_12__sbox_inst_com_w_inst_n449,
         round_inst_S_12__sbox_inst_com_w_inst_n448,
         round_inst_S_12__sbox_inst_com_w_inst_n447,
         round_inst_S_12__sbox_inst_com_w_inst_n446,
         round_inst_S_12__sbox_inst_com_w_inst_n445,
         round_inst_S_12__sbox_inst_com_w_inst_n444,
         round_inst_S_12__sbox_inst_com_w_inst_n443,
         round_inst_S_12__sbox_inst_com_w_inst_n442,
         round_inst_S_12__sbox_inst_com_w_inst_n441,
         round_inst_S_12__sbox_inst_com_w_inst_n440,
         round_inst_S_12__sbox_inst_com_w_inst_n439,
         round_inst_S_12__sbox_inst_com_w_inst_n438,
         round_inst_S_12__sbox_inst_com_w_inst_n437,
         round_inst_S_12__sbox_inst_com_w_inst_n436,
         round_inst_S_12__sbox_inst_com_w_inst_n435,
         round_inst_S_12__sbox_inst_com_w_inst_n434,
         round_inst_S_12__sbox_inst_com_w_inst_n433,
         round_inst_S_12__sbox_inst_com_w_inst_n432,
         round_inst_S_12__sbox_inst_com_w_inst_n431,
         round_inst_S_12__sbox_inst_com_w_inst_n430,
         round_inst_S_12__sbox_inst_com_w_inst_n429,
         round_inst_S_12__sbox_inst_com_w_inst_n428,
         round_inst_S_12__sbox_inst_com_w_inst_n427,
         round_inst_S_12__sbox_inst_com_w_inst_n426,
         round_inst_S_12__sbox_inst_com_w_inst_n425,
         round_inst_S_12__sbox_inst_com_w_inst_n424,
         round_inst_S_12__sbox_inst_com_w_inst_n423,
         round_inst_S_12__sbox_inst_com_w_inst_n422,
         round_inst_S_12__sbox_inst_com_w_inst_n421,
         round_inst_S_12__sbox_inst_com_w_inst_n420,
         round_inst_S_12__sbox_inst_com_w_inst_n419,
         round_inst_S_12__sbox_inst_com_w_inst_n418,
         round_inst_S_12__sbox_inst_com_w_inst_n417,
         round_inst_S_12__sbox_inst_com_w_inst_n416,
         round_inst_S_12__sbox_inst_com_w_inst_n415,
         round_inst_S_12__sbox_inst_com_w_inst_n414,
         round_inst_S_12__sbox_inst_com_w_inst_n413,
         round_inst_S_12__sbox_inst_com_w_inst_n412,
         round_inst_S_12__sbox_inst_com_w_inst_n411,
         round_inst_S_12__sbox_inst_com_w_inst_n410,
         round_inst_S_12__sbox_inst_com_w_inst_n409,
         round_inst_S_12__sbox_inst_com_w_inst_n408,
         round_inst_S_12__sbox_inst_com_w_inst_n407,
         round_inst_S_12__sbox_inst_com_w_inst_n406,
         round_inst_S_12__sbox_inst_com_w_inst_n405,
         round_inst_S_12__sbox_inst_com_w_inst_n404,
         round_inst_S_12__sbox_inst_com_w_inst_n403,
         round_inst_S_12__sbox_inst_com_w_inst_n402,
         round_inst_S_12__sbox_inst_com_w_inst_n401,
         round_inst_S_12__sbox_inst_com_w_inst_n400,
         round_inst_S_12__sbox_inst_com_w_inst_n399,
         round_inst_S_12__sbox_inst_com_w_inst_n398,
         round_inst_S_12__sbox_inst_com_w_inst_n397,
         round_inst_S_12__sbox_inst_com_w_inst_n396,
         round_inst_S_12__sbox_inst_com_x_inst_n512,
         round_inst_S_12__sbox_inst_com_x_inst_n511,
         round_inst_S_12__sbox_inst_com_x_inst_n510,
         round_inst_S_12__sbox_inst_com_x_inst_n509,
         round_inst_S_12__sbox_inst_com_x_inst_n508,
         round_inst_S_12__sbox_inst_com_x_inst_n507,
         round_inst_S_12__sbox_inst_com_x_inst_n506,
         round_inst_S_12__sbox_inst_com_x_inst_n505,
         round_inst_S_12__sbox_inst_com_x_inst_n504,
         round_inst_S_12__sbox_inst_com_x_inst_n503,
         round_inst_S_12__sbox_inst_com_x_inst_n502,
         round_inst_S_12__sbox_inst_com_x_inst_n501,
         round_inst_S_12__sbox_inst_com_x_inst_n500,
         round_inst_S_12__sbox_inst_com_x_inst_n499,
         round_inst_S_12__sbox_inst_com_x_inst_n498,
         round_inst_S_12__sbox_inst_com_x_inst_n497,
         round_inst_S_12__sbox_inst_com_x_inst_n496,
         round_inst_S_12__sbox_inst_com_x_inst_n495,
         round_inst_S_12__sbox_inst_com_x_inst_n494,
         round_inst_S_12__sbox_inst_com_x_inst_n493,
         round_inst_S_12__sbox_inst_com_x_inst_n492,
         round_inst_S_12__sbox_inst_com_x_inst_n491,
         round_inst_S_12__sbox_inst_com_x_inst_n490,
         round_inst_S_12__sbox_inst_com_x_inst_n489,
         round_inst_S_12__sbox_inst_com_x_inst_n488,
         round_inst_S_12__sbox_inst_com_x_inst_n487,
         round_inst_S_12__sbox_inst_com_x_inst_n486,
         round_inst_S_12__sbox_inst_com_x_inst_n485,
         round_inst_S_12__sbox_inst_com_x_inst_n484,
         round_inst_S_12__sbox_inst_com_x_inst_n483,
         round_inst_S_12__sbox_inst_com_x_inst_n482,
         round_inst_S_12__sbox_inst_com_x_inst_n481,
         round_inst_S_12__sbox_inst_com_x_inst_n480,
         round_inst_S_12__sbox_inst_com_x_inst_n479,
         round_inst_S_12__sbox_inst_com_x_inst_n478,
         round_inst_S_12__sbox_inst_com_x_inst_n477,
         round_inst_S_12__sbox_inst_com_x_inst_n476,
         round_inst_S_12__sbox_inst_com_x_inst_n475,
         round_inst_S_12__sbox_inst_com_x_inst_n474,
         round_inst_S_12__sbox_inst_com_x_inst_n473,
         round_inst_S_12__sbox_inst_com_x_inst_n472,
         round_inst_S_12__sbox_inst_com_x_inst_n471,
         round_inst_S_12__sbox_inst_com_x_inst_n470,
         round_inst_S_12__sbox_inst_com_x_inst_n469,
         round_inst_S_12__sbox_inst_com_x_inst_n468,
         round_inst_S_12__sbox_inst_com_x_inst_n467,
         round_inst_S_12__sbox_inst_com_x_inst_n466,
         round_inst_S_12__sbox_inst_com_x_inst_n465,
         round_inst_S_12__sbox_inst_com_x_inst_n464,
         round_inst_S_12__sbox_inst_com_x_inst_n463,
         round_inst_S_12__sbox_inst_com_x_inst_n462,
         round_inst_S_12__sbox_inst_com_x_inst_n461,
         round_inst_S_12__sbox_inst_com_x_inst_n460,
         round_inst_S_12__sbox_inst_com_x_inst_n459,
         round_inst_S_12__sbox_inst_com_x_inst_n458,
         round_inst_S_12__sbox_inst_com_x_inst_n457,
         round_inst_S_12__sbox_inst_com_x_inst_n456,
         round_inst_S_12__sbox_inst_com_x_inst_n455,
         round_inst_S_12__sbox_inst_com_x_inst_n454,
         round_inst_S_12__sbox_inst_com_x_inst_n453,
         round_inst_S_12__sbox_inst_com_x_inst_n452,
         round_inst_S_12__sbox_inst_com_x_inst_n451,
         round_inst_S_12__sbox_inst_com_x_inst_n450,
         round_inst_S_12__sbox_inst_com_x_inst_n449,
         round_inst_S_12__sbox_inst_com_x_inst_n448,
         round_inst_S_12__sbox_inst_com_x_inst_n447,
         round_inst_S_12__sbox_inst_com_x_inst_n446,
         round_inst_S_12__sbox_inst_com_x_inst_n445,
         round_inst_S_12__sbox_inst_com_x_inst_n444,
         round_inst_S_12__sbox_inst_com_x_inst_n443,
         round_inst_S_12__sbox_inst_com_x_inst_n442,
         round_inst_S_12__sbox_inst_com_x_inst_n441,
         round_inst_S_12__sbox_inst_com_x_inst_n440,
         round_inst_S_12__sbox_inst_com_x_inst_n439,
         round_inst_S_12__sbox_inst_com_x_inst_n438,
         round_inst_S_12__sbox_inst_com_x_inst_n437,
         round_inst_S_12__sbox_inst_com_x_inst_n436,
         round_inst_S_12__sbox_inst_com_x_inst_n435,
         round_inst_S_12__sbox_inst_com_x_inst_n434,
         round_inst_S_12__sbox_inst_com_x_inst_n433,
         round_inst_S_12__sbox_inst_com_x_inst_n432,
         round_inst_S_12__sbox_inst_com_x_inst_n431,
         round_inst_S_12__sbox_inst_com_x_inst_n430,
         round_inst_S_12__sbox_inst_com_x_inst_n429,
         round_inst_S_12__sbox_inst_com_x_inst_n428,
         round_inst_S_12__sbox_inst_com_x_inst_n427,
         round_inst_S_12__sbox_inst_com_x_inst_n426,
         round_inst_S_12__sbox_inst_com_x_inst_n425,
         round_inst_S_12__sbox_inst_com_x_inst_n424,
         round_inst_S_12__sbox_inst_com_x_inst_n423,
         round_inst_S_12__sbox_inst_com_x_inst_n422,
         round_inst_S_12__sbox_inst_com_x_inst_n421,
         round_inst_S_12__sbox_inst_com_x_inst_n420,
         round_inst_S_12__sbox_inst_com_x_inst_n419,
         round_inst_S_12__sbox_inst_com_x_inst_n418,
         round_inst_S_12__sbox_inst_com_x_inst_n417,
         round_inst_S_12__sbox_inst_com_x_inst_n416,
         round_inst_S_12__sbox_inst_com_x_inst_n415,
         round_inst_S_12__sbox_inst_com_x_inst_n414,
         round_inst_S_12__sbox_inst_com_x_inst_n413,
         round_inst_S_12__sbox_inst_com_x_inst_n412,
         round_inst_S_12__sbox_inst_com_x_inst_n411,
         round_inst_S_12__sbox_inst_com_x_inst_n410,
         round_inst_S_12__sbox_inst_com_x_inst_n409,
         round_inst_S_12__sbox_inst_com_x_inst_n408,
         round_inst_S_12__sbox_inst_com_x_inst_n407,
         round_inst_S_12__sbox_inst_com_x_inst_n406,
         round_inst_S_12__sbox_inst_com_x_inst_n405,
         round_inst_S_12__sbox_inst_com_x_inst_n404,
         round_inst_S_12__sbox_inst_com_x_inst_n403,
         round_inst_S_12__sbox_inst_com_x_inst_n402,
         round_inst_S_12__sbox_inst_com_x_inst_n401,
         round_inst_S_12__sbox_inst_com_x_inst_n400,
         round_inst_S_12__sbox_inst_com_x_inst_n399,
         round_inst_S_12__sbox_inst_com_x_inst_n398,
         round_inst_S_12__sbox_inst_com_x_inst_n397,
         round_inst_S_12__sbox_inst_com_x_inst_n396,
         round_inst_S_12__sbox_inst_com_x_inst_n395,
         round_inst_S_12__sbox_inst_com_x_inst_n394,
         round_inst_S_12__sbox_inst_com_x_inst_n393,
         round_inst_S_12__sbox_inst_com_x_inst_n392,
         round_inst_S_12__sbox_inst_com_x_inst_n391,
         round_inst_S_12__sbox_inst_com_x_inst_n390,
         round_inst_S_12__sbox_inst_com_x_inst_n389,
         round_inst_S_12__sbox_inst_com_x_inst_n388,
         round_inst_S_12__sbox_inst_com_x_inst_n387,
         round_inst_S_12__sbox_inst_com_x_inst_n386,
         round_inst_S_12__sbox_inst_com_x_inst_n385,
         round_inst_S_12__sbox_inst_com_x_inst_n384,
         round_inst_S_12__sbox_inst_com_x_inst_n383,
         round_inst_S_12__sbox_inst_com_x_inst_n382,
         round_inst_S_12__sbox_inst_com_x_inst_n381,
         round_inst_S_12__sbox_inst_com_y_inst_n519,
         round_inst_S_12__sbox_inst_com_y_inst_n518,
         round_inst_S_12__sbox_inst_com_y_inst_n517,
         round_inst_S_12__sbox_inst_com_y_inst_n516,
         round_inst_S_12__sbox_inst_com_y_inst_n515,
         round_inst_S_12__sbox_inst_com_y_inst_n514,
         round_inst_S_12__sbox_inst_com_y_inst_n513,
         round_inst_S_12__sbox_inst_com_y_inst_n512,
         round_inst_S_12__sbox_inst_com_y_inst_n511,
         round_inst_S_12__sbox_inst_com_y_inst_n510,
         round_inst_S_12__sbox_inst_com_y_inst_n509,
         round_inst_S_12__sbox_inst_com_y_inst_n508,
         round_inst_S_12__sbox_inst_com_y_inst_n507,
         round_inst_S_12__sbox_inst_com_y_inst_n506,
         round_inst_S_12__sbox_inst_com_y_inst_n505,
         round_inst_S_12__sbox_inst_com_y_inst_n504,
         round_inst_S_12__sbox_inst_com_y_inst_n503,
         round_inst_S_12__sbox_inst_com_y_inst_n502,
         round_inst_S_12__sbox_inst_com_y_inst_n501,
         round_inst_S_12__sbox_inst_com_y_inst_n500,
         round_inst_S_12__sbox_inst_com_y_inst_n499,
         round_inst_S_12__sbox_inst_com_y_inst_n498,
         round_inst_S_12__sbox_inst_com_y_inst_n497,
         round_inst_S_12__sbox_inst_com_y_inst_n496,
         round_inst_S_12__sbox_inst_com_y_inst_n495,
         round_inst_S_12__sbox_inst_com_y_inst_n494,
         round_inst_S_12__sbox_inst_com_y_inst_n493,
         round_inst_S_12__sbox_inst_com_y_inst_n492,
         round_inst_S_12__sbox_inst_com_y_inst_n491,
         round_inst_S_12__sbox_inst_com_y_inst_n490,
         round_inst_S_12__sbox_inst_com_y_inst_n489,
         round_inst_S_12__sbox_inst_com_y_inst_n488,
         round_inst_S_12__sbox_inst_com_y_inst_n487,
         round_inst_S_12__sbox_inst_com_y_inst_n486,
         round_inst_S_12__sbox_inst_com_y_inst_n485,
         round_inst_S_12__sbox_inst_com_y_inst_n484,
         round_inst_S_12__sbox_inst_com_y_inst_n483,
         round_inst_S_12__sbox_inst_com_y_inst_n482,
         round_inst_S_12__sbox_inst_com_y_inst_n481,
         round_inst_S_12__sbox_inst_com_y_inst_n480,
         round_inst_S_12__sbox_inst_com_y_inst_n479,
         round_inst_S_12__sbox_inst_com_y_inst_n478,
         round_inst_S_12__sbox_inst_com_y_inst_n477,
         round_inst_S_12__sbox_inst_com_y_inst_n476,
         round_inst_S_12__sbox_inst_com_y_inst_n475,
         round_inst_S_12__sbox_inst_com_y_inst_n474,
         round_inst_S_12__sbox_inst_com_y_inst_n473,
         round_inst_S_12__sbox_inst_com_y_inst_n472,
         round_inst_S_12__sbox_inst_com_y_inst_n471,
         round_inst_S_12__sbox_inst_com_y_inst_n470,
         round_inst_S_12__sbox_inst_com_y_inst_n469,
         round_inst_S_12__sbox_inst_com_y_inst_n468,
         round_inst_S_12__sbox_inst_com_y_inst_n467,
         round_inst_S_12__sbox_inst_com_y_inst_n466,
         round_inst_S_12__sbox_inst_com_y_inst_n465,
         round_inst_S_12__sbox_inst_com_y_inst_n464,
         round_inst_S_12__sbox_inst_com_y_inst_n463,
         round_inst_S_12__sbox_inst_com_y_inst_n462,
         round_inst_S_12__sbox_inst_com_y_inst_n461,
         round_inst_S_12__sbox_inst_com_y_inst_n460,
         round_inst_S_12__sbox_inst_com_y_inst_n459,
         round_inst_S_12__sbox_inst_com_y_inst_n458,
         round_inst_S_12__sbox_inst_com_y_inst_n457,
         round_inst_S_12__sbox_inst_com_y_inst_n456,
         round_inst_S_12__sbox_inst_com_y_inst_n455,
         round_inst_S_12__sbox_inst_com_y_inst_n454,
         round_inst_S_12__sbox_inst_com_y_inst_n453,
         round_inst_S_12__sbox_inst_com_y_inst_n452,
         round_inst_S_12__sbox_inst_com_y_inst_n451,
         round_inst_S_12__sbox_inst_com_y_inst_n450,
         round_inst_S_12__sbox_inst_com_y_inst_n449,
         round_inst_S_12__sbox_inst_com_y_inst_n448,
         round_inst_S_12__sbox_inst_com_y_inst_n447,
         round_inst_S_12__sbox_inst_com_y_inst_n446,
         round_inst_S_12__sbox_inst_com_y_inst_n445,
         round_inst_S_12__sbox_inst_com_y_inst_n444,
         round_inst_S_12__sbox_inst_com_y_inst_n443,
         round_inst_S_12__sbox_inst_com_y_inst_n442,
         round_inst_S_12__sbox_inst_com_y_inst_n441,
         round_inst_S_12__sbox_inst_com_y_inst_n440,
         round_inst_S_12__sbox_inst_com_y_inst_n439,
         round_inst_S_12__sbox_inst_com_y_inst_n438,
         round_inst_S_12__sbox_inst_com_y_inst_n437,
         round_inst_S_12__sbox_inst_com_y_inst_n436,
         round_inst_S_12__sbox_inst_com_y_inst_n435,
         round_inst_S_12__sbox_inst_com_y_inst_n434,
         round_inst_S_12__sbox_inst_com_y_inst_n433,
         round_inst_S_12__sbox_inst_com_y_inst_n432,
         round_inst_S_12__sbox_inst_com_y_inst_n431,
         round_inst_S_12__sbox_inst_com_y_inst_n430,
         round_inst_S_12__sbox_inst_com_y_inst_n429,
         round_inst_S_12__sbox_inst_com_y_inst_n428,
         round_inst_S_12__sbox_inst_com_y_inst_n427,
         round_inst_S_12__sbox_inst_com_y_inst_n426,
         round_inst_S_12__sbox_inst_com_y_inst_n425,
         round_inst_S_12__sbox_inst_com_y_inst_n424,
         round_inst_S_12__sbox_inst_com_y_inst_n423,
         round_inst_S_12__sbox_inst_com_y_inst_n422,
         round_inst_S_12__sbox_inst_com_y_inst_n421,
         round_inst_S_12__sbox_inst_com_y_inst_n420,
         round_inst_S_12__sbox_inst_com_y_inst_n419,
         round_inst_S_12__sbox_inst_com_y_inst_n418,
         round_inst_S_12__sbox_inst_com_y_inst_n417,
         round_inst_S_12__sbox_inst_com_y_inst_n416,
         round_inst_S_12__sbox_inst_com_y_inst_n415,
         round_inst_S_12__sbox_inst_com_y_inst_n414,
         round_inst_S_12__sbox_inst_com_y_inst_n413,
         round_inst_S_12__sbox_inst_com_y_inst_n412,
         round_inst_S_12__sbox_inst_com_y_inst_n411,
         round_inst_S_12__sbox_inst_com_y_inst_n410,
         round_inst_S_12__sbox_inst_com_y_inst_n409,
         round_inst_S_12__sbox_inst_com_y_inst_n408,
         round_inst_S_12__sbox_inst_com_y_inst_n407,
         round_inst_S_12__sbox_inst_com_y_inst_n406,
         round_inst_S_12__sbox_inst_com_y_inst_n405,
         round_inst_S_12__sbox_inst_com_y_inst_n404,
         round_inst_S_12__sbox_inst_com_y_inst_n403,
         round_inst_S_12__sbox_inst_com_y_inst_n402,
         round_inst_S_12__sbox_inst_com_y_inst_n401,
         round_inst_S_12__sbox_inst_com_y_inst_n400,
         round_inst_S_12__sbox_inst_com_y_inst_n399,
         round_inst_S_12__sbox_inst_com_y_inst_n398,
         round_inst_S_12__sbox_inst_com_y_inst_n397,
         round_inst_S_12__sbox_inst_com_y_inst_n396,
         round_inst_S_12__sbox_inst_com_y_inst_n395,
         round_inst_S_12__sbox_inst_com_y_inst_n394,
         round_inst_S_12__sbox_inst_com_y_inst_n393,
         round_inst_S_12__sbox_inst_com_y_inst_n392,
         round_inst_S_12__sbox_inst_com_y_inst_n391,
         round_inst_S_12__sbox_inst_com_y_inst_n390,
         round_inst_S_12__sbox_inst_com_y_inst_n389,
         round_inst_S_12__sbox_inst_com_y_inst_n388,
         round_inst_S_12__sbox_inst_com_y_inst_n387,
         round_inst_S_12__sbox_inst_com_y_inst_n386,
         round_inst_S_12__sbox_inst_com_z_inst_n517,
         round_inst_S_12__sbox_inst_com_z_inst_n516,
         round_inst_S_12__sbox_inst_com_z_inst_n515,
         round_inst_S_12__sbox_inst_com_z_inst_n514,
         round_inst_S_12__sbox_inst_com_z_inst_n513,
         round_inst_S_12__sbox_inst_com_z_inst_n512,
         round_inst_S_12__sbox_inst_com_z_inst_n511,
         round_inst_S_12__sbox_inst_com_z_inst_n510,
         round_inst_S_12__sbox_inst_com_z_inst_n509,
         round_inst_S_12__sbox_inst_com_z_inst_n508,
         round_inst_S_12__sbox_inst_com_z_inst_n507,
         round_inst_S_12__sbox_inst_com_z_inst_n506,
         round_inst_S_12__sbox_inst_com_z_inst_n505,
         round_inst_S_12__sbox_inst_com_z_inst_n504,
         round_inst_S_12__sbox_inst_com_z_inst_n503,
         round_inst_S_12__sbox_inst_com_z_inst_n502,
         round_inst_S_12__sbox_inst_com_z_inst_n501,
         round_inst_S_12__sbox_inst_com_z_inst_n500,
         round_inst_S_12__sbox_inst_com_z_inst_n499,
         round_inst_S_12__sbox_inst_com_z_inst_n498,
         round_inst_S_12__sbox_inst_com_z_inst_n497,
         round_inst_S_12__sbox_inst_com_z_inst_n496,
         round_inst_S_12__sbox_inst_com_z_inst_n495,
         round_inst_S_12__sbox_inst_com_z_inst_n494,
         round_inst_S_12__sbox_inst_com_z_inst_n493,
         round_inst_S_12__sbox_inst_com_z_inst_n492,
         round_inst_S_12__sbox_inst_com_z_inst_n491,
         round_inst_S_12__sbox_inst_com_z_inst_n490,
         round_inst_S_12__sbox_inst_com_z_inst_n489,
         round_inst_S_12__sbox_inst_com_z_inst_n488,
         round_inst_S_12__sbox_inst_com_z_inst_n487,
         round_inst_S_12__sbox_inst_com_z_inst_n486,
         round_inst_S_12__sbox_inst_com_z_inst_n485,
         round_inst_S_12__sbox_inst_com_z_inst_n484,
         round_inst_S_12__sbox_inst_com_z_inst_n483,
         round_inst_S_12__sbox_inst_com_z_inst_n482,
         round_inst_S_12__sbox_inst_com_z_inst_n481,
         round_inst_S_12__sbox_inst_com_z_inst_n480,
         round_inst_S_12__sbox_inst_com_z_inst_n479,
         round_inst_S_12__sbox_inst_com_z_inst_n478,
         round_inst_S_12__sbox_inst_com_z_inst_n477,
         round_inst_S_12__sbox_inst_com_z_inst_n476,
         round_inst_S_12__sbox_inst_com_z_inst_n475,
         round_inst_S_12__sbox_inst_com_z_inst_n474,
         round_inst_S_12__sbox_inst_com_z_inst_n473,
         round_inst_S_12__sbox_inst_com_z_inst_n472,
         round_inst_S_12__sbox_inst_com_z_inst_n471,
         round_inst_S_12__sbox_inst_com_z_inst_n470,
         round_inst_S_12__sbox_inst_com_z_inst_n469,
         round_inst_S_12__sbox_inst_com_z_inst_n468,
         round_inst_S_12__sbox_inst_com_z_inst_n467,
         round_inst_S_12__sbox_inst_com_z_inst_n466,
         round_inst_S_12__sbox_inst_com_z_inst_n465,
         round_inst_S_12__sbox_inst_com_z_inst_n464,
         round_inst_S_12__sbox_inst_com_z_inst_n463,
         round_inst_S_12__sbox_inst_com_z_inst_n462,
         round_inst_S_12__sbox_inst_com_z_inst_n461,
         round_inst_S_12__sbox_inst_com_z_inst_n460,
         round_inst_S_12__sbox_inst_com_z_inst_n459,
         round_inst_S_12__sbox_inst_com_z_inst_n458,
         round_inst_S_12__sbox_inst_com_z_inst_n457,
         round_inst_S_12__sbox_inst_com_z_inst_n456,
         round_inst_S_12__sbox_inst_com_z_inst_n455,
         round_inst_S_12__sbox_inst_com_z_inst_n454,
         round_inst_S_12__sbox_inst_com_z_inst_n453,
         round_inst_S_12__sbox_inst_com_z_inst_n452,
         round_inst_S_12__sbox_inst_com_z_inst_n451,
         round_inst_S_12__sbox_inst_com_z_inst_n450,
         round_inst_S_12__sbox_inst_com_z_inst_n449,
         round_inst_S_12__sbox_inst_com_z_inst_n448,
         round_inst_S_12__sbox_inst_com_z_inst_n447,
         round_inst_S_12__sbox_inst_com_z_inst_n446,
         round_inst_S_12__sbox_inst_com_z_inst_n445,
         round_inst_S_12__sbox_inst_com_z_inst_n444,
         round_inst_S_12__sbox_inst_com_z_inst_n443,
         round_inst_S_12__sbox_inst_com_z_inst_n442,
         round_inst_S_12__sbox_inst_com_z_inst_n441,
         round_inst_S_12__sbox_inst_com_z_inst_n440,
         round_inst_S_12__sbox_inst_com_z_inst_n439,
         round_inst_S_12__sbox_inst_com_z_inst_n438,
         round_inst_S_12__sbox_inst_com_z_inst_n437,
         round_inst_S_12__sbox_inst_com_z_inst_n436,
         round_inst_S_12__sbox_inst_com_z_inst_n435,
         round_inst_S_12__sbox_inst_com_z_inst_n434,
         round_inst_S_12__sbox_inst_com_z_inst_n433,
         round_inst_S_12__sbox_inst_com_z_inst_n432,
         round_inst_S_12__sbox_inst_com_z_inst_n431,
         round_inst_S_12__sbox_inst_com_z_inst_n430,
         round_inst_S_12__sbox_inst_com_z_inst_n429,
         round_inst_S_12__sbox_inst_com_z_inst_n428,
         round_inst_S_12__sbox_inst_com_z_inst_n427,
         round_inst_S_12__sbox_inst_com_z_inst_n426,
         round_inst_S_12__sbox_inst_com_z_inst_n425,
         round_inst_S_12__sbox_inst_com_z_inst_n424,
         round_inst_S_12__sbox_inst_com_z_inst_n423,
         round_inst_S_12__sbox_inst_com_z_inst_n422,
         round_inst_S_12__sbox_inst_com_z_inst_n421,
         round_inst_S_12__sbox_inst_com_z_inst_n420,
         round_inst_S_12__sbox_inst_com_z_inst_n419,
         round_inst_S_12__sbox_inst_com_z_inst_n418,
         round_inst_S_12__sbox_inst_com_z_inst_n417,
         round_inst_S_12__sbox_inst_com_z_inst_n416,
         round_inst_S_12__sbox_inst_com_z_inst_n415,
         round_inst_S_12__sbox_inst_com_z_inst_n414,
         round_inst_S_12__sbox_inst_com_z_inst_n413,
         round_inst_S_12__sbox_inst_com_z_inst_n412,
         round_inst_S_12__sbox_inst_com_z_inst_n411,
         round_inst_S_12__sbox_inst_com_z_inst_n410,
         round_inst_S_12__sbox_inst_com_z_inst_n409,
         round_inst_S_12__sbox_inst_com_z_inst_n408,
         round_inst_S_12__sbox_inst_com_z_inst_n407,
         round_inst_S_12__sbox_inst_com_z_inst_n406,
         round_inst_S_12__sbox_inst_com_z_inst_n405,
         round_inst_S_12__sbox_inst_com_z_inst_n404,
         round_inst_S_12__sbox_inst_com_z_inst_n403,
         round_inst_S_12__sbox_inst_com_z_inst_n402,
         round_inst_S_12__sbox_inst_com_z_inst_n401,
         round_inst_S_12__sbox_inst_com_z_inst_n400,
         round_inst_S_12__sbox_inst_com_z_inst_n399,
         round_inst_S_12__sbox_inst_com_z_inst_n398,
         round_inst_S_12__sbox_inst_com_z_inst_n397,
         round_inst_S_12__sbox_inst_com_z_inst_n396,
         round_inst_S_12__sbox_inst_com_z_inst_n395,
         round_inst_S_12__sbox_inst_com_z_inst_n394,
         round_inst_S_12__sbox_inst_com_z_inst_n393,
         round_inst_S_12__sbox_inst_com_z_inst_n392,
         round_inst_S_12__sbox_inst_com_z_inst_n391,
         round_inst_S_12__sbox_inst_com_z_inst_n390,
         round_inst_S_13__sbox_inst_n4, round_inst_S_13__sbox_inst_n3,
         round_inst_S_13__sbox_inst_n2, round_inst_S_13__sbox_inst_n1,
         round_inst_S_13__sbox_inst_com_w_inst_n531,
         round_inst_S_13__sbox_inst_com_w_inst_n530,
         round_inst_S_13__sbox_inst_com_w_inst_n529,
         round_inst_S_13__sbox_inst_com_w_inst_n528,
         round_inst_S_13__sbox_inst_com_w_inst_n527,
         round_inst_S_13__sbox_inst_com_w_inst_n526,
         round_inst_S_13__sbox_inst_com_w_inst_n525,
         round_inst_S_13__sbox_inst_com_w_inst_n524,
         round_inst_S_13__sbox_inst_com_w_inst_n523,
         round_inst_S_13__sbox_inst_com_w_inst_n522,
         round_inst_S_13__sbox_inst_com_w_inst_n521,
         round_inst_S_13__sbox_inst_com_w_inst_n520,
         round_inst_S_13__sbox_inst_com_w_inst_n519,
         round_inst_S_13__sbox_inst_com_w_inst_n518,
         round_inst_S_13__sbox_inst_com_w_inst_n517,
         round_inst_S_13__sbox_inst_com_w_inst_n516,
         round_inst_S_13__sbox_inst_com_w_inst_n515,
         round_inst_S_13__sbox_inst_com_w_inst_n514,
         round_inst_S_13__sbox_inst_com_w_inst_n513,
         round_inst_S_13__sbox_inst_com_w_inst_n512,
         round_inst_S_13__sbox_inst_com_w_inst_n511,
         round_inst_S_13__sbox_inst_com_w_inst_n510,
         round_inst_S_13__sbox_inst_com_w_inst_n509,
         round_inst_S_13__sbox_inst_com_w_inst_n508,
         round_inst_S_13__sbox_inst_com_w_inst_n507,
         round_inst_S_13__sbox_inst_com_w_inst_n506,
         round_inst_S_13__sbox_inst_com_w_inst_n505,
         round_inst_S_13__sbox_inst_com_w_inst_n504,
         round_inst_S_13__sbox_inst_com_w_inst_n503,
         round_inst_S_13__sbox_inst_com_w_inst_n502,
         round_inst_S_13__sbox_inst_com_w_inst_n501,
         round_inst_S_13__sbox_inst_com_w_inst_n500,
         round_inst_S_13__sbox_inst_com_w_inst_n499,
         round_inst_S_13__sbox_inst_com_w_inst_n498,
         round_inst_S_13__sbox_inst_com_w_inst_n497,
         round_inst_S_13__sbox_inst_com_w_inst_n496,
         round_inst_S_13__sbox_inst_com_w_inst_n495,
         round_inst_S_13__sbox_inst_com_w_inst_n494,
         round_inst_S_13__sbox_inst_com_w_inst_n493,
         round_inst_S_13__sbox_inst_com_w_inst_n492,
         round_inst_S_13__sbox_inst_com_w_inst_n491,
         round_inst_S_13__sbox_inst_com_w_inst_n490,
         round_inst_S_13__sbox_inst_com_w_inst_n489,
         round_inst_S_13__sbox_inst_com_w_inst_n488,
         round_inst_S_13__sbox_inst_com_w_inst_n487,
         round_inst_S_13__sbox_inst_com_w_inst_n486,
         round_inst_S_13__sbox_inst_com_w_inst_n485,
         round_inst_S_13__sbox_inst_com_w_inst_n484,
         round_inst_S_13__sbox_inst_com_w_inst_n483,
         round_inst_S_13__sbox_inst_com_w_inst_n482,
         round_inst_S_13__sbox_inst_com_w_inst_n481,
         round_inst_S_13__sbox_inst_com_w_inst_n480,
         round_inst_S_13__sbox_inst_com_w_inst_n479,
         round_inst_S_13__sbox_inst_com_w_inst_n478,
         round_inst_S_13__sbox_inst_com_w_inst_n477,
         round_inst_S_13__sbox_inst_com_w_inst_n476,
         round_inst_S_13__sbox_inst_com_w_inst_n475,
         round_inst_S_13__sbox_inst_com_w_inst_n474,
         round_inst_S_13__sbox_inst_com_w_inst_n473,
         round_inst_S_13__sbox_inst_com_w_inst_n472,
         round_inst_S_13__sbox_inst_com_w_inst_n471,
         round_inst_S_13__sbox_inst_com_w_inst_n470,
         round_inst_S_13__sbox_inst_com_w_inst_n469,
         round_inst_S_13__sbox_inst_com_w_inst_n468,
         round_inst_S_13__sbox_inst_com_w_inst_n467,
         round_inst_S_13__sbox_inst_com_w_inst_n466,
         round_inst_S_13__sbox_inst_com_w_inst_n465,
         round_inst_S_13__sbox_inst_com_w_inst_n464,
         round_inst_S_13__sbox_inst_com_w_inst_n463,
         round_inst_S_13__sbox_inst_com_w_inst_n462,
         round_inst_S_13__sbox_inst_com_w_inst_n461,
         round_inst_S_13__sbox_inst_com_w_inst_n460,
         round_inst_S_13__sbox_inst_com_w_inst_n459,
         round_inst_S_13__sbox_inst_com_w_inst_n458,
         round_inst_S_13__sbox_inst_com_w_inst_n457,
         round_inst_S_13__sbox_inst_com_w_inst_n456,
         round_inst_S_13__sbox_inst_com_w_inst_n455,
         round_inst_S_13__sbox_inst_com_w_inst_n454,
         round_inst_S_13__sbox_inst_com_w_inst_n453,
         round_inst_S_13__sbox_inst_com_w_inst_n452,
         round_inst_S_13__sbox_inst_com_w_inst_n451,
         round_inst_S_13__sbox_inst_com_w_inst_n450,
         round_inst_S_13__sbox_inst_com_w_inst_n449,
         round_inst_S_13__sbox_inst_com_w_inst_n448,
         round_inst_S_13__sbox_inst_com_w_inst_n447,
         round_inst_S_13__sbox_inst_com_w_inst_n446,
         round_inst_S_13__sbox_inst_com_w_inst_n445,
         round_inst_S_13__sbox_inst_com_w_inst_n444,
         round_inst_S_13__sbox_inst_com_w_inst_n443,
         round_inst_S_13__sbox_inst_com_w_inst_n442,
         round_inst_S_13__sbox_inst_com_w_inst_n441,
         round_inst_S_13__sbox_inst_com_w_inst_n440,
         round_inst_S_13__sbox_inst_com_w_inst_n439,
         round_inst_S_13__sbox_inst_com_w_inst_n438,
         round_inst_S_13__sbox_inst_com_w_inst_n437,
         round_inst_S_13__sbox_inst_com_w_inst_n436,
         round_inst_S_13__sbox_inst_com_w_inst_n435,
         round_inst_S_13__sbox_inst_com_w_inst_n434,
         round_inst_S_13__sbox_inst_com_w_inst_n433,
         round_inst_S_13__sbox_inst_com_w_inst_n432,
         round_inst_S_13__sbox_inst_com_w_inst_n431,
         round_inst_S_13__sbox_inst_com_w_inst_n430,
         round_inst_S_13__sbox_inst_com_w_inst_n429,
         round_inst_S_13__sbox_inst_com_w_inst_n428,
         round_inst_S_13__sbox_inst_com_w_inst_n427,
         round_inst_S_13__sbox_inst_com_w_inst_n426,
         round_inst_S_13__sbox_inst_com_w_inst_n425,
         round_inst_S_13__sbox_inst_com_w_inst_n424,
         round_inst_S_13__sbox_inst_com_w_inst_n423,
         round_inst_S_13__sbox_inst_com_w_inst_n422,
         round_inst_S_13__sbox_inst_com_w_inst_n421,
         round_inst_S_13__sbox_inst_com_w_inst_n420,
         round_inst_S_13__sbox_inst_com_w_inst_n419,
         round_inst_S_13__sbox_inst_com_w_inst_n418,
         round_inst_S_13__sbox_inst_com_w_inst_n417,
         round_inst_S_13__sbox_inst_com_w_inst_n416,
         round_inst_S_13__sbox_inst_com_w_inst_n415,
         round_inst_S_13__sbox_inst_com_w_inst_n414,
         round_inst_S_13__sbox_inst_com_w_inst_n413,
         round_inst_S_13__sbox_inst_com_w_inst_n412,
         round_inst_S_13__sbox_inst_com_w_inst_n411,
         round_inst_S_13__sbox_inst_com_w_inst_n410,
         round_inst_S_13__sbox_inst_com_w_inst_n409,
         round_inst_S_13__sbox_inst_com_w_inst_n408,
         round_inst_S_13__sbox_inst_com_w_inst_n407,
         round_inst_S_13__sbox_inst_com_w_inst_n406,
         round_inst_S_13__sbox_inst_com_w_inst_n405,
         round_inst_S_13__sbox_inst_com_w_inst_n404,
         round_inst_S_13__sbox_inst_com_w_inst_n403,
         round_inst_S_13__sbox_inst_com_w_inst_n402,
         round_inst_S_13__sbox_inst_com_w_inst_n401,
         round_inst_S_13__sbox_inst_com_w_inst_n400,
         round_inst_S_13__sbox_inst_com_w_inst_n399,
         round_inst_S_13__sbox_inst_com_w_inst_n398,
         round_inst_S_13__sbox_inst_com_w_inst_n397,
         round_inst_S_13__sbox_inst_com_w_inst_n396,
         round_inst_S_13__sbox_inst_com_x_inst_n518,
         round_inst_S_13__sbox_inst_com_x_inst_n517,
         round_inst_S_13__sbox_inst_com_x_inst_n516,
         round_inst_S_13__sbox_inst_com_x_inst_n515,
         round_inst_S_13__sbox_inst_com_x_inst_n514,
         round_inst_S_13__sbox_inst_com_x_inst_n513,
         round_inst_S_13__sbox_inst_com_x_inst_n512,
         round_inst_S_13__sbox_inst_com_x_inst_n511,
         round_inst_S_13__sbox_inst_com_x_inst_n510,
         round_inst_S_13__sbox_inst_com_x_inst_n509,
         round_inst_S_13__sbox_inst_com_x_inst_n508,
         round_inst_S_13__sbox_inst_com_x_inst_n507,
         round_inst_S_13__sbox_inst_com_x_inst_n506,
         round_inst_S_13__sbox_inst_com_x_inst_n505,
         round_inst_S_13__sbox_inst_com_x_inst_n504,
         round_inst_S_13__sbox_inst_com_x_inst_n503,
         round_inst_S_13__sbox_inst_com_x_inst_n502,
         round_inst_S_13__sbox_inst_com_x_inst_n501,
         round_inst_S_13__sbox_inst_com_x_inst_n500,
         round_inst_S_13__sbox_inst_com_x_inst_n499,
         round_inst_S_13__sbox_inst_com_x_inst_n498,
         round_inst_S_13__sbox_inst_com_x_inst_n497,
         round_inst_S_13__sbox_inst_com_x_inst_n496,
         round_inst_S_13__sbox_inst_com_x_inst_n495,
         round_inst_S_13__sbox_inst_com_x_inst_n494,
         round_inst_S_13__sbox_inst_com_x_inst_n493,
         round_inst_S_13__sbox_inst_com_x_inst_n492,
         round_inst_S_13__sbox_inst_com_x_inst_n491,
         round_inst_S_13__sbox_inst_com_x_inst_n490,
         round_inst_S_13__sbox_inst_com_x_inst_n489,
         round_inst_S_13__sbox_inst_com_x_inst_n488,
         round_inst_S_13__sbox_inst_com_x_inst_n487,
         round_inst_S_13__sbox_inst_com_x_inst_n486,
         round_inst_S_13__sbox_inst_com_x_inst_n485,
         round_inst_S_13__sbox_inst_com_x_inst_n484,
         round_inst_S_13__sbox_inst_com_x_inst_n483,
         round_inst_S_13__sbox_inst_com_x_inst_n482,
         round_inst_S_13__sbox_inst_com_x_inst_n481,
         round_inst_S_13__sbox_inst_com_x_inst_n480,
         round_inst_S_13__sbox_inst_com_x_inst_n479,
         round_inst_S_13__sbox_inst_com_x_inst_n478,
         round_inst_S_13__sbox_inst_com_x_inst_n477,
         round_inst_S_13__sbox_inst_com_x_inst_n476,
         round_inst_S_13__sbox_inst_com_x_inst_n475,
         round_inst_S_13__sbox_inst_com_x_inst_n474,
         round_inst_S_13__sbox_inst_com_x_inst_n473,
         round_inst_S_13__sbox_inst_com_x_inst_n472,
         round_inst_S_13__sbox_inst_com_x_inst_n471,
         round_inst_S_13__sbox_inst_com_x_inst_n470,
         round_inst_S_13__sbox_inst_com_x_inst_n469,
         round_inst_S_13__sbox_inst_com_x_inst_n468,
         round_inst_S_13__sbox_inst_com_x_inst_n467,
         round_inst_S_13__sbox_inst_com_x_inst_n466,
         round_inst_S_13__sbox_inst_com_x_inst_n465,
         round_inst_S_13__sbox_inst_com_x_inst_n464,
         round_inst_S_13__sbox_inst_com_x_inst_n463,
         round_inst_S_13__sbox_inst_com_x_inst_n462,
         round_inst_S_13__sbox_inst_com_x_inst_n461,
         round_inst_S_13__sbox_inst_com_x_inst_n460,
         round_inst_S_13__sbox_inst_com_x_inst_n459,
         round_inst_S_13__sbox_inst_com_x_inst_n458,
         round_inst_S_13__sbox_inst_com_x_inst_n457,
         round_inst_S_13__sbox_inst_com_x_inst_n456,
         round_inst_S_13__sbox_inst_com_x_inst_n455,
         round_inst_S_13__sbox_inst_com_x_inst_n454,
         round_inst_S_13__sbox_inst_com_x_inst_n453,
         round_inst_S_13__sbox_inst_com_x_inst_n452,
         round_inst_S_13__sbox_inst_com_x_inst_n451,
         round_inst_S_13__sbox_inst_com_x_inst_n450,
         round_inst_S_13__sbox_inst_com_x_inst_n449,
         round_inst_S_13__sbox_inst_com_x_inst_n448,
         round_inst_S_13__sbox_inst_com_x_inst_n447,
         round_inst_S_13__sbox_inst_com_x_inst_n446,
         round_inst_S_13__sbox_inst_com_x_inst_n445,
         round_inst_S_13__sbox_inst_com_x_inst_n444,
         round_inst_S_13__sbox_inst_com_x_inst_n443,
         round_inst_S_13__sbox_inst_com_x_inst_n442,
         round_inst_S_13__sbox_inst_com_x_inst_n441,
         round_inst_S_13__sbox_inst_com_x_inst_n440,
         round_inst_S_13__sbox_inst_com_x_inst_n439,
         round_inst_S_13__sbox_inst_com_x_inst_n438,
         round_inst_S_13__sbox_inst_com_x_inst_n437,
         round_inst_S_13__sbox_inst_com_x_inst_n436,
         round_inst_S_13__sbox_inst_com_x_inst_n435,
         round_inst_S_13__sbox_inst_com_x_inst_n434,
         round_inst_S_13__sbox_inst_com_x_inst_n433,
         round_inst_S_13__sbox_inst_com_x_inst_n432,
         round_inst_S_13__sbox_inst_com_x_inst_n431,
         round_inst_S_13__sbox_inst_com_x_inst_n430,
         round_inst_S_13__sbox_inst_com_x_inst_n429,
         round_inst_S_13__sbox_inst_com_x_inst_n428,
         round_inst_S_13__sbox_inst_com_x_inst_n427,
         round_inst_S_13__sbox_inst_com_x_inst_n426,
         round_inst_S_13__sbox_inst_com_x_inst_n425,
         round_inst_S_13__sbox_inst_com_x_inst_n424,
         round_inst_S_13__sbox_inst_com_x_inst_n423,
         round_inst_S_13__sbox_inst_com_x_inst_n422,
         round_inst_S_13__sbox_inst_com_x_inst_n421,
         round_inst_S_13__sbox_inst_com_x_inst_n420,
         round_inst_S_13__sbox_inst_com_x_inst_n419,
         round_inst_S_13__sbox_inst_com_x_inst_n418,
         round_inst_S_13__sbox_inst_com_x_inst_n417,
         round_inst_S_13__sbox_inst_com_x_inst_n416,
         round_inst_S_13__sbox_inst_com_x_inst_n415,
         round_inst_S_13__sbox_inst_com_x_inst_n414,
         round_inst_S_13__sbox_inst_com_x_inst_n413,
         round_inst_S_13__sbox_inst_com_x_inst_n412,
         round_inst_S_13__sbox_inst_com_x_inst_n411,
         round_inst_S_13__sbox_inst_com_x_inst_n410,
         round_inst_S_13__sbox_inst_com_x_inst_n409,
         round_inst_S_13__sbox_inst_com_x_inst_n408,
         round_inst_S_13__sbox_inst_com_x_inst_n407,
         round_inst_S_13__sbox_inst_com_x_inst_n406,
         round_inst_S_13__sbox_inst_com_x_inst_n405,
         round_inst_S_13__sbox_inst_com_x_inst_n404,
         round_inst_S_13__sbox_inst_com_x_inst_n403,
         round_inst_S_13__sbox_inst_com_x_inst_n402,
         round_inst_S_13__sbox_inst_com_x_inst_n401,
         round_inst_S_13__sbox_inst_com_x_inst_n400,
         round_inst_S_13__sbox_inst_com_x_inst_n399,
         round_inst_S_13__sbox_inst_com_x_inst_n398,
         round_inst_S_13__sbox_inst_com_x_inst_n397,
         round_inst_S_13__sbox_inst_com_x_inst_n396,
         round_inst_S_13__sbox_inst_com_x_inst_n395,
         round_inst_S_13__sbox_inst_com_x_inst_n394,
         round_inst_S_13__sbox_inst_com_x_inst_n393,
         round_inst_S_13__sbox_inst_com_x_inst_n392,
         round_inst_S_13__sbox_inst_com_x_inst_n391,
         round_inst_S_13__sbox_inst_com_x_inst_n390,
         round_inst_S_13__sbox_inst_com_x_inst_n389,
         round_inst_S_13__sbox_inst_com_x_inst_n388,
         round_inst_S_13__sbox_inst_com_x_inst_n387,
         round_inst_S_13__sbox_inst_com_x_inst_n386,
         round_inst_S_13__sbox_inst_com_x_inst_n385,
         round_inst_S_13__sbox_inst_com_x_inst_n384,
         round_inst_S_13__sbox_inst_com_x_inst_n383,
         round_inst_S_13__sbox_inst_com_x_inst_n382,
         round_inst_S_13__sbox_inst_com_x_inst_n381,
         round_inst_S_13__sbox_inst_com_x_inst_n380,
         round_inst_S_13__sbox_inst_com_y_inst_n517,
         round_inst_S_13__sbox_inst_com_y_inst_n516,
         round_inst_S_13__sbox_inst_com_y_inst_n515,
         round_inst_S_13__sbox_inst_com_y_inst_n514,
         round_inst_S_13__sbox_inst_com_y_inst_n513,
         round_inst_S_13__sbox_inst_com_y_inst_n512,
         round_inst_S_13__sbox_inst_com_y_inst_n511,
         round_inst_S_13__sbox_inst_com_y_inst_n510,
         round_inst_S_13__sbox_inst_com_y_inst_n509,
         round_inst_S_13__sbox_inst_com_y_inst_n508,
         round_inst_S_13__sbox_inst_com_y_inst_n507,
         round_inst_S_13__sbox_inst_com_y_inst_n506,
         round_inst_S_13__sbox_inst_com_y_inst_n505,
         round_inst_S_13__sbox_inst_com_y_inst_n504,
         round_inst_S_13__sbox_inst_com_y_inst_n503,
         round_inst_S_13__sbox_inst_com_y_inst_n502,
         round_inst_S_13__sbox_inst_com_y_inst_n501,
         round_inst_S_13__sbox_inst_com_y_inst_n500,
         round_inst_S_13__sbox_inst_com_y_inst_n499,
         round_inst_S_13__sbox_inst_com_y_inst_n498,
         round_inst_S_13__sbox_inst_com_y_inst_n497,
         round_inst_S_13__sbox_inst_com_y_inst_n496,
         round_inst_S_13__sbox_inst_com_y_inst_n495,
         round_inst_S_13__sbox_inst_com_y_inst_n494,
         round_inst_S_13__sbox_inst_com_y_inst_n493,
         round_inst_S_13__sbox_inst_com_y_inst_n492,
         round_inst_S_13__sbox_inst_com_y_inst_n491,
         round_inst_S_13__sbox_inst_com_y_inst_n490,
         round_inst_S_13__sbox_inst_com_y_inst_n489,
         round_inst_S_13__sbox_inst_com_y_inst_n488,
         round_inst_S_13__sbox_inst_com_y_inst_n487,
         round_inst_S_13__sbox_inst_com_y_inst_n486,
         round_inst_S_13__sbox_inst_com_y_inst_n485,
         round_inst_S_13__sbox_inst_com_y_inst_n484,
         round_inst_S_13__sbox_inst_com_y_inst_n483,
         round_inst_S_13__sbox_inst_com_y_inst_n482,
         round_inst_S_13__sbox_inst_com_y_inst_n481,
         round_inst_S_13__sbox_inst_com_y_inst_n480,
         round_inst_S_13__sbox_inst_com_y_inst_n479,
         round_inst_S_13__sbox_inst_com_y_inst_n478,
         round_inst_S_13__sbox_inst_com_y_inst_n477,
         round_inst_S_13__sbox_inst_com_y_inst_n476,
         round_inst_S_13__sbox_inst_com_y_inst_n475,
         round_inst_S_13__sbox_inst_com_y_inst_n474,
         round_inst_S_13__sbox_inst_com_y_inst_n473,
         round_inst_S_13__sbox_inst_com_y_inst_n472,
         round_inst_S_13__sbox_inst_com_y_inst_n471,
         round_inst_S_13__sbox_inst_com_y_inst_n470,
         round_inst_S_13__sbox_inst_com_y_inst_n469,
         round_inst_S_13__sbox_inst_com_y_inst_n468,
         round_inst_S_13__sbox_inst_com_y_inst_n467,
         round_inst_S_13__sbox_inst_com_y_inst_n466,
         round_inst_S_13__sbox_inst_com_y_inst_n465,
         round_inst_S_13__sbox_inst_com_y_inst_n464,
         round_inst_S_13__sbox_inst_com_y_inst_n463,
         round_inst_S_13__sbox_inst_com_y_inst_n462,
         round_inst_S_13__sbox_inst_com_y_inst_n461,
         round_inst_S_13__sbox_inst_com_y_inst_n460,
         round_inst_S_13__sbox_inst_com_y_inst_n459,
         round_inst_S_13__sbox_inst_com_y_inst_n458,
         round_inst_S_13__sbox_inst_com_y_inst_n457,
         round_inst_S_13__sbox_inst_com_y_inst_n456,
         round_inst_S_13__sbox_inst_com_y_inst_n455,
         round_inst_S_13__sbox_inst_com_y_inst_n454,
         round_inst_S_13__sbox_inst_com_y_inst_n453,
         round_inst_S_13__sbox_inst_com_y_inst_n452,
         round_inst_S_13__sbox_inst_com_y_inst_n451,
         round_inst_S_13__sbox_inst_com_y_inst_n450,
         round_inst_S_13__sbox_inst_com_y_inst_n449,
         round_inst_S_13__sbox_inst_com_y_inst_n448,
         round_inst_S_13__sbox_inst_com_y_inst_n447,
         round_inst_S_13__sbox_inst_com_y_inst_n446,
         round_inst_S_13__sbox_inst_com_y_inst_n445,
         round_inst_S_13__sbox_inst_com_y_inst_n444,
         round_inst_S_13__sbox_inst_com_y_inst_n443,
         round_inst_S_13__sbox_inst_com_y_inst_n442,
         round_inst_S_13__sbox_inst_com_y_inst_n441,
         round_inst_S_13__sbox_inst_com_y_inst_n440,
         round_inst_S_13__sbox_inst_com_y_inst_n439,
         round_inst_S_13__sbox_inst_com_y_inst_n438,
         round_inst_S_13__sbox_inst_com_y_inst_n437,
         round_inst_S_13__sbox_inst_com_y_inst_n436,
         round_inst_S_13__sbox_inst_com_y_inst_n435,
         round_inst_S_13__sbox_inst_com_y_inst_n434,
         round_inst_S_13__sbox_inst_com_y_inst_n433,
         round_inst_S_13__sbox_inst_com_y_inst_n432,
         round_inst_S_13__sbox_inst_com_y_inst_n431,
         round_inst_S_13__sbox_inst_com_y_inst_n430,
         round_inst_S_13__sbox_inst_com_y_inst_n429,
         round_inst_S_13__sbox_inst_com_y_inst_n428,
         round_inst_S_13__sbox_inst_com_y_inst_n427,
         round_inst_S_13__sbox_inst_com_y_inst_n426,
         round_inst_S_13__sbox_inst_com_y_inst_n425,
         round_inst_S_13__sbox_inst_com_y_inst_n424,
         round_inst_S_13__sbox_inst_com_y_inst_n423,
         round_inst_S_13__sbox_inst_com_y_inst_n422,
         round_inst_S_13__sbox_inst_com_y_inst_n421,
         round_inst_S_13__sbox_inst_com_y_inst_n420,
         round_inst_S_13__sbox_inst_com_y_inst_n419,
         round_inst_S_13__sbox_inst_com_y_inst_n418,
         round_inst_S_13__sbox_inst_com_y_inst_n417,
         round_inst_S_13__sbox_inst_com_y_inst_n416,
         round_inst_S_13__sbox_inst_com_y_inst_n415,
         round_inst_S_13__sbox_inst_com_y_inst_n414,
         round_inst_S_13__sbox_inst_com_y_inst_n413,
         round_inst_S_13__sbox_inst_com_y_inst_n412,
         round_inst_S_13__sbox_inst_com_y_inst_n411,
         round_inst_S_13__sbox_inst_com_y_inst_n410,
         round_inst_S_13__sbox_inst_com_y_inst_n409,
         round_inst_S_13__sbox_inst_com_y_inst_n408,
         round_inst_S_13__sbox_inst_com_y_inst_n407,
         round_inst_S_13__sbox_inst_com_y_inst_n406,
         round_inst_S_13__sbox_inst_com_y_inst_n405,
         round_inst_S_13__sbox_inst_com_y_inst_n404,
         round_inst_S_13__sbox_inst_com_y_inst_n403,
         round_inst_S_13__sbox_inst_com_y_inst_n402,
         round_inst_S_13__sbox_inst_com_y_inst_n401,
         round_inst_S_13__sbox_inst_com_y_inst_n400,
         round_inst_S_13__sbox_inst_com_y_inst_n399,
         round_inst_S_13__sbox_inst_com_y_inst_n398,
         round_inst_S_13__sbox_inst_com_y_inst_n397,
         round_inst_S_13__sbox_inst_com_y_inst_n396,
         round_inst_S_13__sbox_inst_com_y_inst_n395,
         round_inst_S_13__sbox_inst_com_y_inst_n394,
         round_inst_S_13__sbox_inst_com_y_inst_n393,
         round_inst_S_13__sbox_inst_com_y_inst_n392,
         round_inst_S_13__sbox_inst_com_y_inst_n391,
         round_inst_S_13__sbox_inst_com_y_inst_n390,
         round_inst_S_13__sbox_inst_com_y_inst_n389,
         round_inst_S_13__sbox_inst_com_y_inst_n388,
         round_inst_S_13__sbox_inst_com_y_inst_n387,
         round_inst_S_13__sbox_inst_com_y_inst_n386,
         round_inst_S_13__sbox_inst_com_z_inst_n513,
         round_inst_S_13__sbox_inst_com_z_inst_n512,
         round_inst_S_13__sbox_inst_com_z_inst_n511,
         round_inst_S_13__sbox_inst_com_z_inst_n510,
         round_inst_S_13__sbox_inst_com_z_inst_n509,
         round_inst_S_13__sbox_inst_com_z_inst_n508,
         round_inst_S_13__sbox_inst_com_z_inst_n507,
         round_inst_S_13__sbox_inst_com_z_inst_n506,
         round_inst_S_13__sbox_inst_com_z_inst_n505,
         round_inst_S_13__sbox_inst_com_z_inst_n504,
         round_inst_S_13__sbox_inst_com_z_inst_n503,
         round_inst_S_13__sbox_inst_com_z_inst_n502,
         round_inst_S_13__sbox_inst_com_z_inst_n501,
         round_inst_S_13__sbox_inst_com_z_inst_n500,
         round_inst_S_13__sbox_inst_com_z_inst_n499,
         round_inst_S_13__sbox_inst_com_z_inst_n498,
         round_inst_S_13__sbox_inst_com_z_inst_n497,
         round_inst_S_13__sbox_inst_com_z_inst_n496,
         round_inst_S_13__sbox_inst_com_z_inst_n495,
         round_inst_S_13__sbox_inst_com_z_inst_n494,
         round_inst_S_13__sbox_inst_com_z_inst_n493,
         round_inst_S_13__sbox_inst_com_z_inst_n492,
         round_inst_S_13__sbox_inst_com_z_inst_n491,
         round_inst_S_13__sbox_inst_com_z_inst_n490,
         round_inst_S_13__sbox_inst_com_z_inst_n489,
         round_inst_S_13__sbox_inst_com_z_inst_n488,
         round_inst_S_13__sbox_inst_com_z_inst_n487,
         round_inst_S_13__sbox_inst_com_z_inst_n486,
         round_inst_S_13__sbox_inst_com_z_inst_n485,
         round_inst_S_13__sbox_inst_com_z_inst_n484,
         round_inst_S_13__sbox_inst_com_z_inst_n483,
         round_inst_S_13__sbox_inst_com_z_inst_n482,
         round_inst_S_13__sbox_inst_com_z_inst_n481,
         round_inst_S_13__sbox_inst_com_z_inst_n480,
         round_inst_S_13__sbox_inst_com_z_inst_n479,
         round_inst_S_13__sbox_inst_com_z_inst_n478,
         round_inst_S_13__sbox_inst_com_z_inst_n477,
         round_inst_S_13__sbox_inst_com_z_inst_n476,
         round_inst_S_13__sbox_inst_com_z_inst_n475,
         round_inst_S_13__sbox_inst_com_z_inst_n474,
         round_inst_S_13__sbox_inst_com_z_inst_n473,
         round_inst_S_13__sbox_inst_com_z_inst_n472,
         round_inst_S_13__sbox_inst_com_z_inst_n471,
         round_inst_S_13__sbox_inst_com_z_inst_n470,
         round_inst_S_13__sbox_inst_com_z_inst_n469,
         round_inst_S_13__sbox_inst_com_z_inst_n468,
         round_inst_S_13__sbox_inst_com_z_inst_n467,
         round_inst_S_13__sbox_inst_com_z_inst_n466,
         round_inst_S_13__sbox_inst_com_z_inst_n465,
         round_inst_S_13__sbox_inst_com_z_inst_n464,
         round_inst_S_13__sbox_inst_com_z_inst_n463,
         round_inst_S_13__sbox_inst_com_z_inst_n462,
         round_inst_S_13__sbox_inst_com_z_inst_n461,
         round_inst_S_13__sbox_inst_com_z_inst_n460,
         round_inst_S_13__sbox_inst_com_z_inst_n459,
         round_inst_S_13__sbox_inst_com_z_inst_n458,
         round_inst_S_13__sbox_inst_com_z_inst_n457,
         round_inst_S_13__sbox_inst_com_z_inst_n456,
         round_inst_S_13__sbox_inst_com_z_inst_n455,
         round_inst_S_13__sbox_inst_com_z_inst_n454,
         round_inst_S_13__sbox_inst_com_z_inst_n453,
         round_inst_S_13__sbox_inst_com_z_inst_n452,
         round_inst_S_13__sbox_inst_com_z_inst_n451,
         round_inst_S_13__sbox_inst_com_z_inst_n450,
         round_inst_S_13__sbox_inst_com_z_inst_n449,
         round_inst_S_13__sbox_inst_com_z_inst_n448,
         round_inst_S_13__sbox_inst_com_z_inst_n447,
         round_inst_S_13__sbox_inst_com_z_inst_n446,
         round_inst_S_13__sbox_inst_com_z_inst_n445,
         round_inst_S_13__sbox_inst_com_z_inst_n444,
         round_inst_S_13__sbox_inst_com_z_inst_n443,
         round_inst_S_13__sbox_inst_com_z_inst_n442,
         round_inst_S_13__sbox_inst_com_z_inst_n441,
         round_inst_S_13__sbox_inst_com_z_inst_n440,
         round_inst_S_13__sbox_inst_com_z_inst_n439,
         round_inst_S_13__sbox_inst_com_z_inst_n438,
         round_inst_S_13__sbox_inst_com_z_inst_n437,
         round_inst_S_13__sbox_inst_com_z_inst_n436,
         round_inst_S_13__sbox_inst_com_z_inst_n435,
         round_inst_S_13__sbox_inst_com_z_inst_n434,
         round_inst_S_13__sbox_inst_com_z_inst_n433,
         round_inst_S_13__sbox_inst_com_z_inst_n432,
         round_inst_S_13__sbox_inst_com_z_inst_n431,
         round_inst_S_13__sbox_inst_com_z_inst_n430,
         round_inst_S_13__sbox_inst_com_z_inst_n429,
         round_inst_S_13__sbox_inst_com_z_inst_n428,
         round_inst_S_13__sbox_inst_com_z_inst_n427,
         round_inst_S_13__sbox_inst_com_z_inst_n426,
         round_inst_S_13__sbox_inst_com_z_inst_n425,
         round_inst_S_13__sbox_inst_com_z_inst_n424,
         round_inst_S_13__sbox_inst_com_z_inst_n423,
         round_inst_S_13__sbox_inst_com_z_inst_n422,
         round_inst_S_13__sbox_inst_com_z_inst_n421,
         round_inst_S_13__sbox_inst_com_z_inst_n420,
         round_inst_S_13__sbox_inst_com_z_inst_n419,
         round_inst_S_13__sbox_inst_com_z_inst_n418,
         round_inst_S_13__sbox_inst_com_z_inst_n417,
         round_inst_S_13__sbox_inst_com_z_inst_n416,
         round_inst_S_13__sbox_inst_com_z_inst_n415,
         round_inst_S_13__sbox_inst_com_z_inst_n414,
         round_inst_S_13__sbox_inst_com_z_inst_n413,
         round_inst_S_13__sbox_inst_com_z_inst_n412,
         round_inst_S_13__sbox_inst_com_z_inst_n411,
         round_inst_S_13__sbox_inst_com_z_inst_n410,
         round_inst_S_13__sbox_inst_com_z_inst_n409,
         round_inst_S_13__sbox_inst_com_z_inst_n408,
         round_inst_S_13__sbox_inst_com_z_inst_n407,
         round_inst_S_13__sbox_inst_com_z_inst_n406,
         round_inst_S_13__sbox_inst_com_z_inst_n405,
         round_inst_S_13__sbox_inst_com_z_inst_n404,
         round_inst_S_13__sbox_inst_com_z_inst_n403,
         round_inst_S_13__sbox_inst_com_z_inst_n402,
         round_inst_S_13__sbox_inst_com_z_inst_n401,
         round_inst_S_13__sbox_inst_com_z_inst_n400,
         round_inst_S_13__sbox_inst_com_z_inst_n399,
         round_inst_S_13__sbox_inst_com_z_inst_n398,
         round_inst_S_13__sbox_inst_com_z_inst_n397,
         round_inst_S_13__sbox_inst_com_z_inst_n396,
         round_inst_S_13__sbox_inst_com_z_inst_n395,
         round_inst_S_13__sbox_inst_com_z_inst_n394,
         round_inst_S_13__sbox_inst_com_z_inst_n393,
         round_inst_S_13__sbox_inst_com_z_inst_n392,
         round_inst_S_13__sbox_inst_com_z_inst_n391,
         round_inst_S_13__sbox_inst_com_z_inst_n390,
         round_inst_S_14__sbox_inst_n6, round_inst_S_14__sbox_inst_n5,
         round_inst_S_14__sbox_inst_n4, round_inst_S_14__sbox_inst_n3,
         round_inst_S_14__sbox_inst_n2, round_inst_S_14__sbox_inst_n1,
         round_inst_S_14__sbox_inst_com_w_inst_n529,
         round_inst_S_14__sbox_inst_com_w_inst_n528,
         round_inst_S_14__sbox_inst_com_w_inst_n527,
         round_inst_S_14__sbox_inst_com_w_inst_n526,
         round_inst_S_14__sbox_inst_com_w_inst_n525,
         round_inst_S_14__sbox_inst_com_w_inst_n524,
         round_inst_S_14__sbox_inst_com_w_inst_n523,
         round_inst_S_14__sbox_inst_com_w_inst_n522,
         round_inst_S_14__sbox_inst_com_w_inst_n521,
         round_inst_S_14__sbox_inst_com_w_inst_n520,
         round_inst_S_14__sbox_inst_com_w_inst_n519,
         round_inst_S_14__sbox_inst_com_w_inst_n518,
         round_inst_S_14__sbox_inst_com_w_inst_n517,
         round_inst_S_14__sbox_inst_com_w_inst_n516,
         round_inst_S_14__sbox_inst_com_w_inst_n515,
         round_inst_S_14__sbox_inst_com_w_inst_n514,
         round_inst_S_14__sbox_inst_com_w_inst_n513,
         round_inst_S_14__sbox_inst_com_w_inst_n512,
         round_inst_S_14__sbox_inst_com_w_inst_n511,
         round_inst_S_14__sbox_inst_com_w_inst_n510,
         round_inst_S_14__sbox_inst_com_w_inst_n509,
         round_inst_S_14__sbox_inst_com_w_inst_n508,
         round_inst_S_14__sbox_inst_com_w_inst_n507,
         round_inst_S_14__sbox_inst_com_w_inst_n506,
         round_inst_S_14__sbox_inst_com_w_inst_n505,
         round_inst_S_14__sbox_inst_com_w_inst_n504,
         round_inst_S_14__sbox_inst_com_w_inst_n503,
         round_inst_S_14__sbox_inst_com_w_inst_n502,
         round_inst_S_14__sbox_inst_com_w_inst_n501,
         round_inst_S_14__sbox_inst_com_w_inst_n500,
         round_inst_S_14__sbox_inst_com_w_inst_n499,
         round_inst_S_14__sbox_inst_com_w_inst_n498,
         round_inst_S_14__sbox_inst_com_w_inst_n497,
         round_inst_S_14__sbox_inst_com_w_inst_n496,
         round_inst_S_14__sbox_inst_com_w_inst_n495,
         round_inst_S_14__sbox_inst_com_w_inst_n494,
         round_inst_S_14__sbox_inst_com_w_inst_n493,
         round_inst_S_14__sbox_inst_com_w_inst_n492,
         round_inst_S_14__sbox_inst_com_w_inst_n491,
         round_inst_S_14__sbox_inst_com_w_inst_n490,
         round_inst_S_14__sbox_inst_com_w_inst_n489,
         round_inst_S_14__sbox_inst_com_w_inst_n488,
         round_inst_S_14__sbox_inst_com_w_inst_n487,
         round_inst_S_14__sbox_inst_com_w_inst_n486,
         round_inst_S_14__sbox_inst_com_w_inst_n485,
         round_inst_S_14__sbox_inst_com_w_inst_n484,
         round_inst_S_14__sbox_inst_com_w_inst_n483,
         round_inst_S_14__sbox_inst_com_w_inst_n482,
         round_inst_S_14__sbox_inst_com_w_inst_n481,
         round_inst_S_14__sbox_inst_com_w_inst_n480,
         round_inst_S_14__sbox_inst_com_w_inst_n479,
         round_inst_S_14__sbox_inst_com_w_inst_n478,
         round_inst_S_14__sbox_inst_com_w_inst_n477,
         round_inst_S_14__sbox_inst_com_w_inst_n476,
         round_inst_S_14__sbox_inst_com_w_inst_n475,
         round_inst_S_14__sbox_inst_com_w_inst_n474,
         round_inst_S_14__sbox_inst_com_w_inst_n473,
         round_inst_S_14__sbox_inst_com_w_inst_n472,
         round_inst_S_14__sbox_inst_com_w_inst_n471,
         round_inst_S_14__sbox_inst_com_w_inst_n470,
         round_inst_S_14__sbox_inst_com_w_inst_n469,
         round_inst_S_14__sbox_inst_com_w_inst_n468,
         round_inst_S_14__sbox_inst_com_w_inst_n467,
         round_inst_S_14__sbox_inst_com_w_inst_n466,
         round_inst_S_14__sbox_inst_com_w_inst_n465,
         round_inst_S_14__sbox_inst_com_w_inst_n464,
         round_inst_S_14__sbox_inst_com_w_inst_n463,
         round_inst_S_14__sbox_inst_com_w_inst_n462,
         round_inst_S_14__sbox_inst_com_w_inst_n461,
         round_inst_S_14__sbox_inst_com_w_inst_n460,
         round_inst_S_14__sbox_inst_com_w_inst_n459,
         round_inst_S_14__sbox_inst_com_w_inst_n458,
         round_inst_S_14__sbox_inst_com_w_inst_n457,
         round_inst_S_14__sbox_inst_com_w_inst_n456,
         round_inst_S_14__sbox_inst_com_w_inst_n455,
         round_inst_S_14__sbox_inst_com_w_inst_n454,
         round_inst_S_14__sbox_inst_com_w_inst_n453,
         round_inst_S_14__sbox_inst_com_w_inst_n452,
         round_inst_S_14__sbox_inst_com_w_inst_n451,
         round_inst_S_14__sbox_inst_com_w_inst_n450,
         round_inst_S_14__sbox_inst_com_w_inst_n449,
         round_inst_S_14__sbox_inst_com_w_inst_n448,
         round_inst_S_14__sbox_inst_com_w_inst_n447,
         round_inst_S_14__sbox_inst_com_w_inst_n446,
         round_inst_S_14__sbox_inst_com_w_inst_n445,
         round_inst_S_14__sbox_inst_com_w_inst_n444,
         round_inst_S_14__sbox_inst_com_w_inst_n443,
         round_inst_S_14__sbox_inst_com_w_inst_n442,
         round_inst_S_14__sbox_inst_com_w_inst_n441,
         round_inst_S_14__sbox_inst_com_w_inst_n440,
         round_inst_S_14__sbox_inst_com_w_inst_n439,
         round_inst_S_14__sbox_inst_com_w_inst_n438,
         round_inst_S_14__sbox_inst_com_w_inst_n437,
         round_inst_S_14__sbox_inst_com_w_inst_n436,
         round_inst_S_14__sbox_inst_com_w_inst_n435,
         round_inst_S_14__sbox_inst_com_w_inst_n434,
         round_inst_S_14__sbox_inst_com_w_inst_n433,
         round_inst_S_14__sbox_inst_com_w_inst_n432,
         round_inst_S_14__sbox_inst_com_w_inst_n431,
         round_inst_S_14__sbox_inst_com_w_inst_n430,
         round_inst_S_14__sbox_inst_com_w_inst_n429,
         round_inst_S_14__sbox_inst_com_w_inst_n428,
         round_inst_S_14__sbox_inst_com_w_inst_n427,
         round_inst_S_14__sbox_inst_com_w_inst_n426,
         round_inst_S_14__sbox_inst_com_w_inst_n425,
         round_inst_S_14__sbox_inst_com_w_inst_n424,
         round_inst_S_14__sbox_inst_com_w_inst_n423,
         round_inst_S_14__sbox_inst_com_w_inst_n422,
         round_inst_S_14__sbox_inst_com_w_inst_n421,
         round_inst_S_14__sbox_inst_com_w_inst_n420,
         round_inst_S_14__sbox_inst_com_w_inst_n419,
         round_inst_S_14__sbox_inst_com_w_inst_n418,
         round_inst_S_14__sbox_inst_com_w_inst_n417,
         round_inst_S_14__sbox_inst_com_w_inst_n416,
         round_inst_S_14__sbox_inst_com_w_inst_n415,
         round_inst_S_14__sbox_inst_com_w_inst_n414,
         round_inst_S_14__sbox_inst_com_w_inst_n413,
         round_inst_S_14__sbox_inst_com_w_inst_n412,
         round_inst_S_14__sbox_inst_com_w_inst_n411,
         round_inst_S_14__sbox_inst_com_w_inst_n410,
         round_inst_S_14__sbox_inst_com_w_inst_n409,
         round_inst_S_14__sbox_inst_com_w_inst_n408,
         round_inst_S_14__sbox_inst_com_w_inst_n407,
         round_inst_S_14__sbox_inst_com_w_inst_n406,
         round_inst_S_14__sbox_inst_com_w_inst_n405,
         round_inst_S_14__sbox_inst_com_w_inst_n404,
         round_inst_S_14__sbox_inst_com_w_inst_n403,
         round_inst_S_14__sbox_inst_com_w_inst_n402,
         round_inst_S_14__sbox_inst_com_w_inst_n401,
         round_inst_S_14__sbox_inst_com_w_inst_n400,
         round_inst_S_14__sbox_inst_com_w_inst_n399,
         round_inst_S_14__sbox_inst_com_w_inst_n398,
         round_inst_S_14__sbox_inst_com_w_inst_n397,
         round_inst_S_14__sbox_inst_com_w_inst_n396,
         round_inst_S_14__sbox_inst_com_x_inst_n512,
         round_inst_S_14__sbox_inst_com_x_inst_n511,
         round_inst_S_14__sbox_inst_com_x_inst_n510,
         round_inst_S_14__sbox_inst_com_x_inst_n509,
         round_inst_S_14__sbox_inst_com_x_inst_n508,
         round_inst_S_14__sbox_inst_com_x_inst_n507,
         round_inst_S_14__sbox_inst_com_x_inst_n506,
         round_inst_S_14__sbox_inst_com_x_inst_n505,
         round_inst_S_14__sbox_inst_com_x_inst_n504,
         round_inst_S_14__sbox_inst_com_x_inst_n503,
         round_inst_S_14__sbox_inst_com_x_inst_n502,
         round_inst_S_14__sbox_inst_com_x_inst_n501,
         round_inst_S_14__sbox_inst_com_x_inst_n500,
         round_inst_S_14__sbox_inst_com_x_inst_n499,
         round_inst_S_14__sbox_inst_com_x_inst_n498,
         round_inst_S_14__sbox_inst_com_x_inst_n497,
         round_inst_S_14__sbox_inst_com_x_inst_n496,
         round_inst_S_14__sbox_inst_com_x_inst_n495,
         round_inst_S_14__sbox_inst_com_x_inst_n494,
         round_inst_S_14__sbox_inst_com_x_inst_n493,
         round_inst_S_14__sbox_inst_com_x_inst_n492,
         round_inst_S_14__sbox_inst_com_x_inst_n491,
         round_inst_S_14__sbox_inst_com_x_inst_n490,
         round_inst_S_14__sbox_inst_com_x_inst_n489,
         round_inst_S_14__sbox_inst_com_x_inst_n488,
         round_inst_S_14__sbox_inst_com_x_inst_n487,
         round_inst_S_14__sbox_inst_com_x_inst_n486,
         round_inst_S_14__sbox_inst_com_x_inst_n485,
         round_inst_S_14__sbox_inst_com_x_inst_n484,
         round_inst_S_14__sbox_inst_com_x_inst_n483,
         round_inst_S_14__sbox_inst_com_x_inst_n482,
         round_inst_S_14__sbox_inst_com_x_inst_n481,
         round_inst_S_14__sbox_inst_com_x_inst_n480,
         round_inst_S_14__sbox_inst_com_x_inst_n479,
         round_inst_S_14__sbox_inst_com_x_inst_n478,
         round_inst_S_14__sbox_inst_com_x_inst_n477,
         round_inst_S_14__sbox_inst_com_x_inst_n476,
         round_inst_S_14__sbox_inst_com_x_inst_n475,
         round_inst_S_14__sbox_inst_com_x_inst_n474,
         round_inst_S_14__sbox_inst_com_x_inst_n473,
         round_inst_S_14__sbox_inst_com_x_inst_n472,
         round_inst_S_14__sbox_inst_com_x_inst_n471,
         round_inst_S_14__sbox_inst_com_x_inst_n470,
         round_inst_S_14__sbox_inst_com_x_inst_n469,
         round_inst_S_14__sbox_inst_com_x_inst_n468,
         round_inst_S_14__sbox_inst_com_x_inst_n467,
         round_inst_S_14__sbox_inst_com_x_inst_n466,
         round_inst_S_14__sbox_inst_com_x_inst_n465,
         round_inst_S_14__sbox_inst_com_x_inst_n464,
         round_inst_S_14__sbox_inst_com_x_inst_n463,
         round_inst_S_14__sbox_inst_com_x_inst_n462,
         round_inst_S_14__sbox_inst_com_x_inst_n461,
         round_inst_S_14__sbox_inst_com_x_inst_n460,
         round_inst_S_14__sbox_inst_com_x_inst_n459,
         round_inst_S_14__sbox_inst_com_x_inst_n458,
         round_inst_S_14__sbox_inst_com_x_inst_n457,
         round_inst_S_14__sbox_inst_com_x_inst_n456,
         round_inst_S_14__sbox_inst_com_x_inst_n455,
         round_inst_S_14__sbox_inst_com_x_inst_n454,
         round_inst_S_14__sbox_inst_com_x_inst_n453,
         round_inst_S_14__sbox_inst_com_x_inst_n452,
         round_inst_S_14__sbox_inst_com_x_inst_n451,
         round_inst_S_14__sbox_inst_com_x_inst_n450,
         round_inst_S_14__sbox_inst_com_x_inst_n449,
         round_inst_S_14__sbox_inst_com_x_inst_n448,
         round_inst_S_14__sbox_inst_com_x_inst_n447,
         round_inst_S_14__sbox_inst_com_x_inst_n446,
         round_inst_S_14__sbox_inst_com_x_inst_n445,
         round_inst_S_14__sbox_inst_com_x_inst_n444,
         round_inst_S_14__sbox_inst_com_x_inst_n443,
         round_inst_S_14__sbox_inst_com_x_inst_n442,
         round_inst_S_14__sbox_inst_com_x_inst_n441,
         round_inst_S_14__sbox_inst_com_x_inst_n440,
         round_inst_S_14__sbox_inst_com_x_inst_n439,
         round_inst_S_14__sbox_inst_com_x_inst_n438,
         round_inst_S_14__sbox_inst_com_x_inst_n437,
         round_inst_S_14__sbox_inst_com_x_inst_n436,
         round_inst_S_14__sbox_inst_com_x_inst_n435,
         round_inst_S_14__sbox_inst_com_x_inst_n434,
         round_inst_S_14__sbox_inst_com_x_inst_n433,
         round_inst_S_14__sbox_inst_com_x_inst_n432,
         round_inst_S_14__sbox_inst_com_x_inst_n431,
         round_inst_S_14__sbox_inst_com_x_inst_n430,
         round_inst_S_14__sbox_inst_com_x_inst_n429,
         round_inst_S_14__sbox_inst_com_x_inst_n428,
         round_inst_S_14__sbox_inst_com_x_inst_n427,
         round_inst_S_14__sbox_inst_com_x_inst_n426,
         round_inst_S_14__sbox_inst_com_x_inst_n425,
         round_inst_S_14__sbox_inst_com_x_inst_n424,
         round_inst_S_14__sbox_inst_com_x_inst_n423,
         round_inst_S_14__sbox_inst_com_x_inst_n422,
         round_inst_S_14__sbox_inst_com_x_inst_n421,
         round_inst_S_14__sbox_inst_com_x_inst_n420,
         round_inst_S_14__sbox_inst_com_x_inst_n419,
         round_inst_S_14__sbox_inst_com_x_inst_n418,
         round_inst_S_14__sbox_inst_com_x_inst_n417,
         round_inst_S_14__sbox_inst_com_x_inst_n416,
         round_inst_S_14__sbox_inst_com_x_inst_n415,
         round_inst_S_14__sbox_inst_com_x_inst_n414,
         round_inst_S_14__sbox_inst_com_x_inst_n413,
         round_inst_S_14__sbox_inst_com_x_inst_n412,
         round_inst_S_14__sbox_inst_com_x_inst_n411,
         round_inst_S_14__sbox_inst_com_x_inst_n410,
         round_inst_S_14__sbox_inst_com_x_inst_n409,
         round_inst_S_14__sbox_inst_com_x_inst_n408,
         round_inst_S_14__sbox_inst_com_x_inst_n407,
         round_inst_S_14__sbox_inst_com_x_inst_n406,
         round_inst_S_14__sbox_inst_com_x_inst_n405,
         round_inst_S_14__sbox_inst_com_x_inst_n404,
         round_inst_S_14__sbox_inst_com_x_inst_n403,
         round_inst_S_14__sbox_inst_com_x_inst_n402,
         round_inst_S_14__sbox_inst_com_x_inst_n401,
         round_inst_S_14__sbox_inst_com_x_inst_n400,
         round_inst_S_14__sbox_inst_com_x_inst_n399,
         round_inst_S_14__sbox_inst_com_x_inst_n398,
         round_inst_S_14__sbox_inst_com_x_inst_n397,
         round_inst_S_14__sbox_inst_com_x_inst_n396,
         round_inst_S_14__sbox_inst_com_x_inst_n395,
         round_inst_S_14__sbox_inst_com_x_inst_n394,
         round_inst_S_14__sbox_inst_com_x_inst_n393,
         round_inst_S_14__sbox_inst_com_x_inst_n392,
         round_inst_S_14__sbox_inst_com_x_inst_n391,
         round_inst_S_14__sbox_inst_com_x_inst_n390,
         round_inst_S_14__sbox_inst_com_x_inst_n389,
         round_inst_S_14__sbox_inst_com_x_inst_n388,
         round_inst_S_14__sbox_inst_com_x_inst_n387,
         round_inst_S_14__sbox_inst_com_x_inst_n386,
         round_inst_S_14__sbox_inst_com_x_inst_n385,
         round_inst_S_14__sbox_inst_com_x_inst_n384,
         round_inst_S_14__sbox_inst_com_x_inst_n383,
         round_inst_S_14__sbox_inst_com_x_inst_n382,
         round_inst_S_14__sbox_inst_com_x_inst_n381,
         round_inst_S_14__sbox_inst_com_y_inst_n519,
         round_inst_S_14__sbox_inst_com_y_inst_n518,
         round_inst_S_14__sbox_inst_com_y_inst_n517,
         round_inst_S_14__sbox_inst_com_y_inst_n516,
         round_inst_S_14__sbox_inst_com_y_inst_n515,
         round_inst_S_14__sbox_inst_com_y_inst_n514,
         round_inst_S_14__sbox_inst_com_y_inst_n513,
         round_inst_S_14__sbox_inst_com_y_inst_n512,
         round_inst_S_14__sbox_inst_com_y_inst_n511,
         round_inst_S_14__sbox_inst_com_y_inst_n510,
         round_inst_S_14__sbox_inst_com_y_inst_n509,
         round_inst_S_14__sbox_inst_com_y_inst_n508,
         round_inst_S_14__sbox_inst_com_y_inst_n507,
         round_inst_S_14__sbox_inst_com_y_inst_n506,
         round_inst_S_14__sbox_inst_com_y_inst_n505,
         round_inst_S_14__sbox_inst_com_y_inst_n504,
         round_inst_S_14__sbox_inst_com_y_inst_n503,
         round_inst_S_14__sbox_inst_com_y_inst_n502,
         round_inst_S_14__sbox_inst_com_y_inst_n501,
         round_inst_S_14__sbox_inst_com_y_inst_n500,
         round_inst_S_14__sbox_inst_com_y_inst_n499,
         round_inst_S_14__sbox_inst_com_y_inst_n498,
         round_inst_S_14__sbox_inst_com_y_inst_n497,
         round_inst_S_14__sbox_inst_com_y_inst_n496,
         round_inst_S_14__sbox_inst_com_y_inst_n495,
         round_inst_S_14__sbox_inst_com_y_inst_n494,
         round_inst_S_14__sbox_inst_com_y_inst_n493,
         round_inst_S_14__sbox_inst_com_y_inst_n492,
         round_inst_S_14__sbox_inst_com_y_inst_n491,
         round_inst_S_14__sbox_inst_com_y_inst_n490,
         round_inst_S_14__sbox_inst_com_y_inst_n489,
         round_inst_S_14__sbox_inst_com_y_inst_n488,
         round_inst_S_14__sbox_inst_com_y_inst_n487,
         round_inst_S_14__sbox_inst_com_y_inst_n486,
         round_inst_S_14__sbox_inst_com_y_inst_n485,
         round_inst_S_14__sbox_inst_com_y_inst_n484,
         round_inst_S_14__sbox_inst_com_y_inst_n483,
         round_inst_S_14__sbox_inst_com_y_inst_n482,
         round_inst_S_14__sbox_inst_com_y_inst_n481,
         round_inst_S_14__sbox_inst_com_y_inst_n480,
         round_inst_S_14__sbox_inst_com_y_inst_n479,
         round_inst_S_14__sbox_inst_com_y_inst_n478,
         round_inst_S_14__sbox_inst_com_y_inst_n477,
         round_inst_S_14__sbox_inst_com_y_inst_n476,
         round_inst_S_14__sbox_inst_com_y_inst_n475,
         round_inst_S_14__sbox_inst_com_y_inst_n474,
         round_inst_S_14__sbox_inst_com_y_inst_n473,
         round_inst_S_14__sbox_inst_com_y_inst_n472,
         round_inst_S_14__sbox_inst_com_y_inst_n471,
         round_inst_S_14__sbox_inst_com_y_inst_n470,
         round_inst_S_14__sbox_inst_com_y_inst_n469,
         round_inst_S_14__sbox_inst_com_y_inst_n468,
         round_inst_S_14__sbox_inst_com_y_inst_n467,
         round_inst_S_14__sbox_inst_com_y_inst_n466,
         round_inst_S_14__sbox_inst_com_y_inst_n465,
         round_inst_S_14__sbox_inst_com_y_inst_n464,
         round_inst_S_14__sbox_inst_com_y_inst_n463,
         round_inst_S_14__sbox_inst_com_y_inst_n462,
         round_inst_S_14__sbox_inst_com_y_inst_n461,
         round_inst_S_14__sbox_inst_com_y_inst_n460,
         round_inst_S_14__sbox_inst_com_y_inst_n459,
         round_inst_S_14__sbox_inst_com_y_inst_n458,
         round_inst_S_14__sbox_inst_com_y_inst_n457,
         round_inst_S_14__sbox_inst_com_y_inst_n456,
         round_inst_S_14__sbox_inst_com_y_inst_n455,
         round_inst_S_14__sbox_inst_com_y_inst_n454,
         round_inst_S_14__sbox_inst_com_y_inst_n453,
         round_inst_S_14__sbox_inst_com_y_inst_n452,
         round_inst_S_14__sbox_inst_com_y_inst_n451,
         round_inst_S_14__sbox_inst_com_y_inst_n450,
         round_inst_S_14__sbox_inst_com_y_inst_n449,
         round_inst_S_14__sbox_inst_com_y_inst_n448,
         round_inst_S_14__sbox_inst_com_y_inst_n447,
         round_inst_S_14__sbox_inst_com_y_inst_n446,
         round_inst_S_14__sbox_inst_com_y_inst_n445,
         round_inst_S_14__sbox_inst_com_y_inst_n444,
         round_inst_S_14__sbox_inst_com_y_inst_n443,
         round_inst_S_14__sbox_inst_com_y_inst_n442,
         round_inst_S_14__sbox_inst_com_y_inst_n441,
         round_inst_S_14__sbox_inst_com_y_inst_n440,
         round_inst_S_14__sbox_inst_com_y_inst_n439,
         round_inst_S_14__sbox_inst_com_y_inst_n438,
         round_inst_S_14__sbox_inst_com_y_inst_n437,
         round_inst_S_14__sbox_inst_com_y_inst_n436,
         round_inst_S_14__sbox_inst_com_y_inst_n435,
         round_inst_S_14__sbox_inst_com_y_inst_n434,
         round_inst_S_14__sbox_inst_com_y_inst_n433,
         round_inst_S_14__sbox_inst_com_y_inst_n432,
         round_inst_S_14__sbox_inst_com_y_inst_n431,
         round_inst_S_14__sbox_inst_com_y_inst_n430,
         round_inst_S_14__sbox_inst_com_y_inst_n429,
         round_inst_S_14__sbox_inst_com_y_inst_n428,
         round_inst_S_14__sbox_inst_com_y_inst_n427,
         round_inst_S_14__sbox_inst_com_y_inst_n426,
         round_inst_S_14__sbox_inst_com_y_inst_n425,
         round_inst_S_14__sbox_inst_com_y_inst_n424,
         round_inst_S_14__sbox_inst_com_y_inst_n423,
         round_inst_S_14__sbox_inst_com_y_inst_n422,
         round_inst_S_14__sbox_inst_com_y_inst_n421,
         round_inst_S_14__sbox_inst_com_y_inst_n420,
         round_inst_S_14__sbox_inst_com_y_inst_n419,
         round_inst_S_14__sbox_inst_com_y_inst_n418,
         round_inst_S_14__sbox_inst_com_y_inst_n417,
         round_inst_S_14__sbox_inst_com_y_inst_n416,
         round_inst_S_14__sbox_inst_com_y_inst_n415,
         round_inst_S_14__sbox_inst_com_y_inst_n414,
         round_inst_S_14__sbox_inst_com_y_inst_n413,
         round_inst_S_14__sbox_inst_com_y_inst_n412,
         round_inst_S_14__sbox_inst_com_y_inst_n411,
         round_inst_S_14__sbox_inst_com_y_inst_n410,
         round_inst_S_14__sbox_inst_com_y_inst_n409,
         round_inst_S_14__sbox_inst_com_y_inst_n408,
         round_inst_S_14__sbox_inst_com_y_inst_n407,
         round_inst_S_14__sbox_inst_com_y_inst_n406,
         round_inst_S_14__sbox_inst_com_y_inst_n405,
         round_inst_S_14__sbox_inst_com_y_inst_n404,
         round_inst_S_14__sbox_inst_com_y_inst_n403,
         round_inst_S_14__sbox_inst_com_y_inst_n402,
         round_inst_S_14__sbox_inst_com_y_inst_n401,
         round_inst_S_14__sbox_inst_com_y_inst_n400,
         round_inst_S_14__sbox_inst_com_y_inst_n399,
         round_inst_S_14__sbox_inst_com_y_inst_n398,
         round_inst_S_14__sbox_inst_com_y_inst_n397,
         round_inst_S_14__sbox_inst_com_y_inst_n396,
         round_inst_S_14__sbox_inst_com_y_inst_n395,
         round_inst_S_14__sbox_inst_com_y_inst_n394,
         round_inst_S_14__sbox_inst_com_y_inst_n393,
         round_inst_S_14__sbox_inst_com_y_inst_n392,
         round_inst_S_14__sbox_inst_com_y_inst_n391,
         round_inst_S_14__sbox_inst_com_y_inst_n390,
         round_inst_S_14__sbox_inst_com_y_inst_n389,
         round_inst_S_14__sbox_inst_com_y_inst_n388,
         round_inst_S_14__sbox_inst_com_y_inst_n387,
         round_inst_S_14__sbox_inst_com_y_inst_n386,
         round_inst_S_14__sbox_inst_com_z_inst_n517,
         round_inst_S_14__sbox_inst_com_z_inst_n516,
         round_inst_S_14__sbox_inst_com_z_inst_n515,
         round_inst_S_14__sbox_inst_com_z_inst_n514,
         round_inst_S_14__sbox_inst_com_z_inst_n513,
         round_inst_S_14__sbox_inst_com_z_inst_n512,
         round_inst_S_14__sbox_inst_com_z_inst_n511,
         round_inst_S_14__sbox_inst_com_z_inst_n510,
         round_inst_S_14__sbox_inst_com_z_inst_n509,
         round_inst_S_14__sbox_inst_com_z_inst_n508,
         round_inst_S_14__sbox_inst_com_z_inst_n507,
         round_inst_S_14__sbox_inst_com_z_inst_n506,
         round_inst_S_14__sbox_inst_com_z_inst_n505,
         round_inst_S_14__sbox_inst_com_z_inst_n504,
         round_inst_S_14__sbox_inst_com_z_inst_n503,
         round_inst_S_14__sbox_inst_com_z_inst_n502,
         round_inst_S_14__sbox_inst_com_z_inst_n501,
         round_inst_S_14__sbox_inst_com_z_inst_n500,
         round_inst_S_14__sbox_inst_com_z_inst_n499,
         round_inst_S_14__sbox_inst_com_z_inst_n498,
         round_inst_S_14__sbox_inst_com_z_inst_n497,
         round_inst_S_14__sbox_inst_com_z_inst_n496,
         round_inst_S_14__sbox_inst_com_z_inst_n495,
         round_inst_S_14__sbox_inst_com_z_inst_n494,
         round_inst_S_14__sbox_inst_com_z_inst_n493,
         round_inst_S_14__sbox_inst_com_z_inst_n492,
         round_inst_S_14__sbox_inst_com_z_inst_n491,
         round_inst_S_14__sbox_inst_com_z_inst_n490,
         round_inst_S_14__sbox_inst_com_z_inst_n489,
         round_inst_S_14__sbox_inst_com_z_inst_n488,
         round_inst_S_14__sbox_inst_com_z_inst_n487,
         round_inst_S_14__sbox_inst_com_z_inst_n486,
         round_inst_S_14__sbox_inst_com_z_inst_n485,
         round_inst_S_14__sbox_inst_com_z_inst_n484,
         round_inst_S_14__sbox_inst_com_z_inst_n483,
         round_inst_S_14__sbox_inst_com_z_inst_n482,
         round_inst_S_14__sbox_inst_com_z_inst_n481,
         round_inst_S_14__sbox_inst_com_z_inst_n480,
         round_inst_S_14__sbox_inst_com_z_inst_n479,
         round_inst_S_14__sbox_inst_com_z_inst_n478,
         round_inst_S_14__sbox_inst_com_z_inst_n477,
         round_inst_S_14__sbox_inst_com_z_inst_n476,
         round_inst_S_14__sbox_inst_com_z_inst_n475,
         round_inst_S_14__sbox_inst_com_z_inst_n474,
         round_inst_S_14__sbox_inst_com_z_inst_n473,
         round_inst_S_14__sbox_inst_com_z_inst_n472,
         round_inst_S_14__sbox_inst_com_z_inst_n471,
         round_inst_S_14__sbox_inst_com_z_inst_n470,
         round_inst_S_14__sbox_inst_com_z_inst_n469,
         round_inst_S_14__sbox_inst_com_z_inst_n468,
         round_inst_S_14__sbox_inst_com_z_inst_n467,
         round_inst_S_14__sbox_inst_com_z_inst_n466,
         round_inst_S_14__sbox_inst_com_z_inst_n465,
         round_inst_S_14__sbox_inst_com_z_inst_n464,
         round_inst_S_14__sbox_inst_com_z_inst_n463,
         round_inst_S_14__sbox_inst_com_z_inst_n462,
         round_inst_S_14__sbox_inst_com_z_inst_n461,
         round_inst_S_14__sbox_inst_com_z_inst_n460,
         round_inst_S_14__sbox_inst_com_z_inst_n459,
         round_inst_S_14__sbox_inst_com_z_inst_n458,
         round_inst_S_14__sbox_inst_com_z_inst_n457,
         round_inst_S_14__sbox_inst_com_z_inst_n456,
         round_inst_S_14__sbox_inst_com_z_inst_n455,
         round_inst_S_14__sbox_inst_com_z_inst_n454,
         round_inst_S_14__sbox_inst_com_z_inst_n453,
         round_inst_S_14__sbox_inst_com_z_inst_n452,
         round_inst_S_14__sbox_inst_com_z_inst_n451,
         round_inst_S_14__sbox_inst_com_z_inst_n450,
         round_inst_S_14__sbox_inst_com_z_inst_n449,
         round_inst_S_14__sbox_inst_com_z_inst_n448,
         round_inst_S_14__sbox_inst_com_z_inst_n447,
         round_inst_S_14__sbox_inst_com_z_inst_n446,
         round_inst_S_14__sbox_inst_com_z_inst_n445,
         round_inst_S_14__sbox_inst_com_z_inst_n444,
         round_inst_S_14__sbox_inst_com_z_inst_n443,
         round_inst_S_14__sbox_inst_com_z_inst_n442,
         round_inst_S_14__sbox_inst_com_z_inst_n441,
         round_inst_S_14__sbox_inst_com_z_inst_n440,
         round_inst_S_14__sbox_inst_com_z_inst_n439,
         round_inst_S_14__sbox_inst_com_z_inst_n438,
         round_inst_S_14__sbox_inst_com_z_inst_n437,
         round_inst_S_14__sbox_inst_com_z_inst_n436,
         round_inst_S_14__sbox_inst_com_z_inst_n435,
         round_inst_S_14__sbox_inst_com_z_inst_n434,
         round_inst_S_14__sbox_inst_com_z_inst_n433,
         round_inst_S_14__sbox_inst_com_z_inst_n432,
         round_inst_S_14__sbox_inst_com_z_inst_n431,
         round_inst_S_14__sbox_inst_com_z_inst_n430,
         round_inst_S_14__sbox_inst_com_z_inst_n429,
         round_inst_S_14__sbox_inst_com_z_inst_n428,
         round_inst_S_14__sbox_inst_com_z_inst_n427,
         round_inst_S_14__sbox_inst_com_z_inst_n426,
         round_inst_S_14__sbox_inst_com_z_inst_n425,
         round_inst_S_14__sbox_inst_com_z_inst_n424,
         round_inst_S_14__sbox_inst_com_z_inst_n423,
         round_inst_S_14__sbox_inst_com_z_inst_n422,
         round_inst_S_14__sbox_inst_com_z_inst_n421,
         round_inst_S_14__sbox_inst_com_z_inst_n420,
         round_inst_S_14__sbox_inst_com_z_inst_n419,
         round_inst_S_14__sbox_inst_com_z_inst_n418,
         round_inst_S_14__sbox_inst_com_z_inst_n417,
         round_inst_S_14__sbox_inst_com_z_inst_n416,
         round_inst_S_14__sbox_inst_com_z_inst_n415,
         round_inst_S_14__sbox_inst_com_z_inst_n414,
         round_inst_S_14__sbox_inst_com_z_inst_n413,
         round_inst_S_14__sbox_inst_com_z_inst_n412,
         round_inst_S_14__sbox_inst_com_z_inst_n411,
         round_inst_S_14__sbox_inst_com_z_inst_n410,
         round_inst_S_14__sbox_inst_com_z_inst_n409,
         round_inst_S_14__sbox_inst_com_z_inst_n408,
         round_inst_S_14__sbox_inst_com_z_inst_n407,
         round_inst_S_14__sbox_inst_com_z_inst_n406,
         round_inst_S_14__sbox_inst_com_z_inst_n405,
         round_inst_S_14__sbox_inst_com_z_inst_n404,
         round_inst_S_14__sbox_inst_com_z_inst_n403,
         round_inst_S_14__sbox_inst_com_z_inst_n402,
         round_inst_S_14__sbox_inst_com_z_inst_n401,
         round_inst_S_14__sbox_inst_com_z_inst_n400,
         round_inst_S_14__sbox_inst_com_z_inst_n399,
         round_inst_S_14__sbox_inst_com_z_inst_n398,
         round_inst_S_14__sbox_inst_com_z_inst_n397,
         round_inst_S_14__sbox_inst_com_z_inst_n396,
         round_inst_S_14__sbox_inst_com_z_inst_n395,
         round_inst_S_14__sbox_inst_com_z_inst_n394,
         round_inst_S_14__sbox_inst_com_z_inst_n393,
         round_inst_S_14__sbox_inst_com_z_inst_n392,
         round_inst_S_14__sbox_inst_com_z_inst_n391,
         round_inst_S_14__sbox_inst_com_z_inst_n390,
         round_inst_S_15__sbox_inst_n6, round_inst_S_15__sbox_inst_n5,
         round_inst_S_15__sbox_inst_n4, round_inst_S_15__sbox_inst_n3,
         round_inst_S_15__sbox_inst_n2, round_inst_S_15__sbox_inst_n1,
         round_inst_S_15__sbox_inst_com_w_inst_n532,
         round_inst_S_15__sbox_inst_com_w_inst_n531,
         round_inst_S_15__sbox_inst_com_w_inst_n530,
         round_inst_S_15__sbox_inst_com_w_inst_n529,
         round_inst_S_15__sbox_inst_com_w_inst_n528,
         round_inst_S_15__sbox_inst_com_w_inst_n527,
         round_inst_S_15__sbox_inst_com_w_inst_n526,
         round_inst_S_15__sbox_inst_com_w_inst_n525,
         round_inst_S_15__sbox_inst_com_w_inst_n524,
         round_inst_S_15__sbox_inst_com_w_inst_n523,
         round_inst_S_15__sbox_inst_com_w_inst_n522,
         round_inst_S_15__sbox_inst_com_w_inst_n521,
         round_inst_S_15__sbox_inst_com_w_inst_n520,
         round_inst_S_15__sbox_inst_com_w_inst_n519,
         round_inst_S_15__sbox_inst_com_w_inst_n518,
         round_inst_S_15__sbox_inst_com_w_inst_n517,
         round_inst_S_15__sbox_inst_com_w_inst_n516,
         round_inst_S_15__sbox_inst_com_w_inst_n515,
         round_inst_S_15__sbox_inst_com_w_inst_n514,
         round_inst_S_15__sbox_inst_com_w_inst_n513,
         round_inst_S_15__sbox_inst_com_w_inst_n512,
         round_inst_S_15__sbox_inst_com_w_inst_n511,
         round_inst_S_15__sbox_inst_com_w_inst_n510,
         round_inst_S_15__sbox_inst_com_w_inst_n509,
         round_inst_S_15__sbox_inst_com_w_inst_n508,
         round_inst_S_15__sbox_inst_com_w_inst_n507,
         round_inst_S_15__sbox_inst_com_w_inst_n506,
         round_inst_S_15__sbox_inst_com_w_inst_n505,
         round_inst_S_15__sbox_inst_com_w_inst_n504,
         round_inst_S_15__sbox_inst_com_w_inst_n503,
         round_inst_S_15__sbox_inst_com_w_inst_n502,
         round_inst_S_15__sbox_inst_com_w_inst_n501,
         round_inst_S_15__sbox_inst_com_w_inst_n500,
         round_inst_S_15__sbox_inst_com_w_inst_n499,
         round_inst_S_15__sbox_inst_com_w_inst_n498,
         round_inst_S_15__sbox_inst_com_w_inst_n497,
         round_inst_S_15__sbox_inst_com_w_inst_n496,
         round_inst_S_15__sbox_inst_com_w_inst_n495,
         round_inst_S_15__sbox_inst_com_w_inst_n494,
         round_inst_S_15__sbox_inst_com_w_inst_n493,
         round_inst_S_15__sbox_inst_com_w_inst_n492,
         round_inst_S_15__sbox_inst_com_w_inst_n491,
         round_inst_S_15__sbox_inst_com_w_inst_n490,
         round_inst_S_15__sbox_inst_com_w_inst_n489,
         round_inst_S_15__sbox_inst_com_w_inst_n488,
         round_inst_S_15__sbox_inst_com_w_inst_n487,
         round_inst_S_15__sbox_inst_com_w_inst_n486,
         round_inst_S_15__sbox_inst_com_w_inst_n485,
         round_inst_S_15__sbox_inst_com_w_inst_n484,
         round_inst_S_15__sbox_inst_com_w_inst_n483,
         round_inst_S_15__sbox_inst_com_w_inst_n482,
         round_inst_S_15__sbox_inst_com_w_inst_n481,
         round_inst_S_15__sbox_inst_com_w_inst_n480,
         round_inst_S_15__sbox_inst_com_w_inst_n479,
         round_inst_S_15__sbox_inst_com_w_inst_n478,
         round_inst_S_15__sbox_inst_com_w_inst_n477,
         round_inst_S_15__sbox_inst_com_w_inst_n476,
         round_inst_S_15__sbox_inst_com_w_inst_n475,
         round_inst_S_15__sbox_inst_com_w_inst_n474,
         round_inst_S_15__sbox_inst_com_w_inst_n473,
         round_inst_S_15__sbox_inst_com_w_inst_n472,
         round_inst_S_15__sbox_inst_com_w_inst_n471,
         round_inst_S_15__sbox_inst_com_w_inst_n470,
         round_inst_S_15__sbox_inst_com_w_inst_n469,
         round_inst_S_15__sbox_inst_com_w_inst_n468,
         round_inst_S_15__sbox_inst_com_w_inst_n467,
         round_inst_S_15__sbox_inst_com_w_inst_n466,
         round_inst_S_15__sbox_inst_com_w_inst_n465,
         round_inst_S_15__sbox_inst_com_w_inst_n464,
         round_inst_S_15__sbox_inst_com_w_inst_n463,
         round_inst_S_15__sbox_inst_com_w_inst_n462,
         round_inst_S_15__sbox_inst_com_w_inst_n461,
         round_inst_S_15__sbox_inst_com_w_inst_n460,
         round_inst_S_15__sbox_inst_com_w_inst_n459,
         round_inst_S_15__sbox_inst_com_w_inst_n458,
         round_inst_S_15__sbox_inst_com_w_inst_n457,
         round_inst_S_15__sbox_inst_com_w_inst_n456,
         round_inst_S_15__sbox_inst_com_w_inst_n455,
         round_inst_S_15__sbox_inst_com_w_inst_n454,
         round_inst_S_15__sbox_inst_com_w_inst_n453,
         round_inst_S_15__sbox_inst_com_w_inst_n452,
         round_inst_S_15__sbox_inst_com_w_inst_n451,
         round_inst_S_15__sbox_inst_com_w_inst_n450,
         round_inst_S_15__sbox_inst_com_w_inst_n449,
         round_inst_S_15__sbox_inst_com_w_inst_n448,
         round_inst_S_15__sbox_inst_com_w_inst_n447,
         round_inst_S_15__sbox_inst_com_w_inst_n446,
         round_inst_S_15__sbox_inst_com_w_inst_n445,
         round_inst_S_15__sbox_inst_com_w_inst_n444,
         round_inst_S_15__sbox_inst_com_w_inst_n443,
         round_inst_S_15__sbox_inst_com_w_inst_n442,
         round_inst_S_15__sbox_inst_com_w_inst_n441,
         round_inst_S_15__sbox_inst_com_w_inst_n440,
         round_inst_S_15__sbox_inst_com_w_inst_n439,
         round_inst_S_15__sbox_inst_com_w_inst_n438,
         round_inst_S_15__sbox_inst_com_w_inst_n437,
         round_inst_S_15__sbox_inst_com_w_inst_n436,
         round_inst_S_15__sbox_inst_com_w_inst_n435,
         round_inst_S_15__sbox_inst_com_w_inst_n434,
         round_inst_S_15__sbox_inst_com_w_inst_n433,
         round_inst_S_15__sbox_inst_com_w_inst_n432,
         round_inst_S_15__sbox_inst_com_w_inst_n431,
         round_inst_S_15__sbox_inst_com_w_inst_n430,
         round_inst_S_15__sbox_inst_com_w_inst_n429,
         round_inst_S_15__sbox_inst_com_w_inst_n428,
         round_inst_S_15__sbox_inst_com_w_inst_n427,
         round_inst_S_15__sbox_inst_com_w_inst_n426,
         round_inst_S_15__sbox_inst_com_w_inst_n425,
         round_inst_S_15__sbox_inst_com_w_inst_n424,
         round_inst_S_15__sbox_inst_com_w_inst_n423,
         round_inst_S_15__sbox_inst_com_w_inst_n422,
         round_inst_S_15__sbox_inst_com_w_inst_n421,
         round_inst_S_15__sbox_inst_com_w_inst_n420,
         round_inst_S_15__sbox_inst_com_w_inst_n419,
         round_inst_S_15__sbox_inst_com_w_inst_n418,
         round_inst_S_15__sbox_inst_com_w_inst_n417,
         round_inst_S_15__sbox_inst_com_w_inst_n416,
         round_inst_S_15__sbox_inst_com_w_inst_n415,
         round_inst_S_15__sbox_inst_com_w_inst_n414,
         round_inst_S_15__sbox_inst_com_w_inst_n413,
         round_inst_S_15__sbox_inst_com_w_inst_n412,
         round_inst_S_15__sbox_inst_com_w_inst_n411,
         round_inst_S_15__sbox_inst_com_w_inst_n410,
         round_inst_S_15__sbox_inst_com_w_inst_n409,
         round_inst_S_15__sbox_inst_com_w_inst_n408,
         round_inst_S_15__sbox_inst_com_w_inst_n407,
         round_inst_S_15__sbox_inst_com_w_inst_n406,
         round_inst_S_15__sbox_inst_com_w_inst_n405,
         round_inst_S_15__sbox_inst_com_w_inst_n404,
         round_inst_S_15__sbox_inst_com_w_inst_n403,
         round_inst_S_15__sbox_inst_com_w_inst_n402,
         round_inst_S_15__sbox_inst_com_w_inst_n401,
         round_inst_S_15__sbox_inst_com_w_inst_n400,
         round_inst_S_15__sbox_inst_com_w_inst_n399,
         round_inst_S_15__sbox_inst_com_w_inst_n398,
         round_inst_S_15__sbox_inst_com_w_inst_n397,
         round_inst_S_15__sbox_inst_com_w_inst_n396,
         round_inst_S_15__sbox_inst_com_x_inst_n511,
         round_inst_S_15__sbox_inst_com_x_inst_n510,
         round_inst_S_15__sbox_inst_com_x_inst_n509,
         round_inst_S_15__sbox_inst_com_x_inst_n508,
         round_inst_S_15__sbox_inst_com_x_inst_n507,
         round_inst_S_15__sbox_inst_com_x_inst_n506,
         round_inst_S_15__sbox_inst_com_x_inst_n505,
         round_inst_S_15__sbox_inst_com_x_inst_n504,
         round_inst_S_15__sbox_inst_com_x_inst_n503,
         round_inst_S_15__sbox_inst_com_x_inst_n502,
         round_inst_S_15__sbox_inst_com_x_inst_n501,
         round_inst_S_15__sbox_inst_com_x_inst_n500,
         round_inst_S_15__sbox_inst_com_x_inst_n499,
         round_inst_S_15__sbox_inst_com_x_inst_n498,
         round_inst_S_15__sbox_inst_com_x_inst_n497,
         round_inst_S_15__sbox_inst_com_x_inst_n496,
         round_inst_S_15__sbox_inst_com_x_inst_n495,
         round_inst_S_15__sbox_inst_com_x_inst_n494,
         round_inst_S_15__sbox_inst_com_x_inst_n493,
         round_inst_S_15__sbox_inst_com_x_inst_n492,
         round_inst_S_15__sbox_inst_com_x_inst_n491,
         round_inst_S_15__sbox_inst_com_x_inst_n490,
         round_inst_S_15__sbox_inst_com_x_inst_n489,
         round_inst_S_15__sbox_inst_com_x_inst_n488,
         round_inst_S_15__sbox_inst_com_x_inst_n487,
         round_inst_S_15__sbox_inst_com_x_inst_n486,
         round_inst_S_15__sbox_inst_com_x_inst_n485,
         round_inst_S_15__sbox_inst_com_x_inst_n484,
         round_inst_S_15__sbox_inst_com_x_inst_n483,
         round_inst_S_15__sbox_inst_com_x_inst_n482,
         round_inst_S_15__sbox_inst_com_x_inst_n481,
         round_inst_S_15__sbox_inst_com_x_inst_n480,
         round_inst_S_15__sbox_inst_com_x_inst_n479,
         round_inst_S_15__sbox_inst_com_x_inst_n478,
         round_inst_S_15__sbox_inst_com_x_inst_n477,
         round_inst_S_15__sbox_inst_com_x_inst_n476,
         round_inst_S_15__sbox_inst_com_x_inst_n475,
         round_inst_S_15__sbox_inst_com_x_inst_n474,
         round_inst_S_15__sbox_inst_com_x_inst_n473,
         round_inst_S_15__sbox_inst_com_x_inst_n472,
         round_inst_S_15__sbox_inst_com_x_inst_n471,
         round_inst_S_15__sbox_inst_com_x_inst_n470,
         round_inst_S_15__sbox_inst_com_x_inst_n469,
         round_inst_S_15__sbox_inst_com_x_inst_n468,
         round_inst_S_15__sbox_inst_com_x_inst_n467,
         round_inst_S_15__sbox_inst_com_x_inst_n466,
         round_inst_S_15__sbox_inst_com_x_inst_n465,
         round_inst_S_15__sbox_inst_com_x_inst_n464,
         round_inst_S_15__sbox_inst_com_x_inst_n463,
         round_inst_S_15__sbox_inst_com_x_inst_n462,
         round_inst_S_15__sbox_inst_com_x_inst_n461,
         round_inst_S_15__sbox_inst_com_x_inst_n460,
         round_inst_S_15__sbox_inst_com_x_inst_n459,
         round_inst_S_15__sbox_inst_com_x_inst_n458,
         round_inst_S_15__sbox_inst_com_x_inst_n457,
         round_inst_S_15__sbox_inst_com_x_inst_n456,
         round_inst_S_15__sbox_inst_com_x_inst_n455,
         round_inst_S_15__sbox_inst_com_x_inst_n454,
         round_inst_S_15__sbox_inst_com_x_inst_n453,
         round_inst_S_15__sbox_inst_com_x_inst_n452,
         round_inst_S_15__sbox_inst_com_x_inst_n451,
         round_inst_S_15__sbox_inst_com_x_inst_n450,
         round_inst_S_15__sbox_inst_com_x_inst_n449,
         round_inst_S_15__sbox_inst_com_x_inst_n448,
         round_inst_S_15__sbox_inst_com_x_inst_n447,
         round_inst_S_15__sbox_inst_com_x_inst_n446,
         round_inst_S_15__sbox_inst_com_x_inst_n445,
         round_inst_S_15__sbox_inst_com_x_inst_n444,
         round_inst_S_15__sbox_inst_com_x_inst_n443,
         round_inst_S_15__sbox_inst_com_x_inst_n442,
         round_inst_S_15__sbox_inst_com_x_inst_n441,
         round_inst_S_15__sbox_inst_com_x_inst_n440,
         round_inst_S_15__sbox_inst_com_x_inst_n439,
         round_inst_S_15__sbox_inst_com_x_inst_n438,
         round_inst_S_15__sbox_inst_com_x_inst_n437,
         round_inst_S_15__sbox_inst_com_x_inst_n436,
         round_inst_S_15__sbox_inst_com_x_inst_n435,
         round_inst_S_15__sbox_inst_com_x_inst_n434,
         round_inst_S_15__sbox_inst_com_x_inst_n433,
         round_inst_S_15__sbox_inst_com_x_inst_n432,
         round_inst_S_15__sbox_inst_com_x_inst_n431,
         round_inst_S_15__sbox_inst_com_x_inst_n430,
         round_inst_S_15__sbox_inst_com_x_inst_n429,
         round_inst_S_15__sbox_inst_com_x_inst_n428,
         round_inst_S_15__sbox_inst_com_x_inst_n427,
         round_inst_S_15__sbox_inst_com_x_inst_n426,
         round_inst_S_15__sbox_inst_com_x_inst_n425,
         round_inst_S_15__sbox_inst_com_x_inst_n424,
         round_inst_S_15__sbox_inst_com_x_inst_n423,
         round_inst_S_15__sbox_inst_com_x_inst_n422,
         round_inst_S_15__sbox_inst_com_x_inst_n421,
         round_inst_S_15__sbox_inst_com_x_inst_n420,
         round_inst_S_15__sbox_inst_com_x_inst_n419,
         round_inst_S_15__sbox_inst_com_x_inst_n418,
         round_inst_S_15__sbox_inst_com_x_inst_n417,
         round_inst_S_15__sbox_inst_com_x_inst_n416,
         round_inst_S_15__sbox_inst_com_x_inst_n415,
         round_inst_S_15__sbox_inst_com_x_inst_n414,
         round_inst_S_15__sbox_inst_com_x_inst_n413,
         round_inst_S_15__sbox_inst_com_x_inst_n412,
         round_inst_S_15__sbox_inst_com_x_inst_n411,
         round_inst_S_15__sbox_inst_com_x_inst_n410,
         round_inst_S_15__sbox_inst_com_x_inst_n409,
         round_inst_S_15__sbox_inst_com_x_inst_n408,
         round_inst_S_15__sbox_inst_com_x_inst_n407,
         round_inst_S_15__sbox_inst_com_x_inst_n406,
         round_inst_S_15__sbox_inst_com_x_inst_n405,
         round_inst_S_15__sbox_inst_com_x_inst_n404,
         round_inst_S_15__sbox_inst_com_x_inst_n403,
         round_inst_S_15__sbox_inst_com_x_inst_n402,
         round_inst_S_15__sbox_inst_com_x_inst_n401,
         round_inst_S_15__sbox_inst_com_x_inst_n400,
         round_inst_S_15__sbox_inst_com_x_inst_n399,
         round_inst_S_15__sbox_inst_com_x_inst_n398,
         round_inst_S_15__sbox_inst_com_x_inst_n397,
         round_inst_S_15__sbox_inst_com_x_inst_n396,
         round_inst_S_15__sbox_inst_com_x_inst_n395,
         round_inst_S_15__sbox_inst_com_x_inst_n394,
         round_inst_S_15__sbox_inst_com_x_inst_n393,
         round_inst_S_15__sbox_inst_com_x_inst_n392,
         round_inst_S_15__sbox_inst_com_x_inst_n391,
         round_inst_S_15__sbox_inst_com_x_inst_n390,
         round_inst_S_15__sbox_inst_com_x_inst_n389,
         round_inst_S_15__sbox_inst_com_x_inst_n388,
         round_inst_S_15__sbox_inst_com_x_inst_n387,
         round_inst_S_15__sbox_inst_com_x_inst_n386,
         round_inst_S_15__sbox_inst_com_x_inst_n385,
         round_inst_S_15__sbox_inst_com_x_inst_n384,
         round_inst_S_15__sbox_inst_com_x_inst_n383,
         round_inst_S_15__sbox_inst_com_x_inst_n382,
         round_inst_S_15__sbox_inst_com_x_inst_n381,
         round_inst_S_15__sbox_inst_com_y_inst_n518,
         round_inst_S_15__sbox_inst_com_y_inst_n517,
         round_inst_S_15__sbox_inst_com_y_inst_n516,
         round_inst_S_15__sbox_inst_com_y_inst_n515,
         round_inst_S_15__sbox_inst_com_y_inst_n514,
         round_inst_S_15__sbox_inst_com_y_inst_n513,
         round_inst_S_15__sbox_inst_com_y_inst_n512,
         round_inst_S_15__sbox_inst_com_y_inst_n511,
         round_inst_S_15__sbox_inst_com_y_inst_n510,
         round_inst_S_15__sbox_inst_com_y_inst_n509,
         round_inst_S_15__sbox_inst_com_y_inst_n508,
         round_inst_S_15__sbox_inst_com_y_inst_n507,
         round_inst_S_15__sbox_inst_com_y_inst_n506,
         round_inst_S_15__sbox_inst_com_y_inst_n505,
         round_inst_S_15__sbox_inst_com_y_inst_n504,
         round_inst_S_15__sbox_inst_com_y_inst_n503,
         round_inst_S_15__sbox_inst_com_y_inst_n502,
         round_inst_S_15__sbox_inst_com_y_inst_n501,
         round_inst_S_15__sbox_inst_com_y_inst_n500,
         round_inst_S_15__sbox_inst_com_y_inst_n499,
         round_inst_S_15__sbox_inst_com_y_inst_n498,
         round_inst_S_15__sbox_inst_com_y_inst_n497,
         round_inst_S_15__sbox_inst_com_y_inst_n496,
         round_inst_S_15__sbox_inst_com_y_inst_n495,
         round_inst_S_15__sbox_inst_com_y_inst_n494,
         round_inst_S_15__sbox_inst_com_y_inst_n493,
         round_inst_S_15__sbox_inst_com_y_inst_n492,
         round_inst_S_15__sbox_inst_com_y_inst_n491,
         round_inst_S_15__sbox_inst_com_y_inst_n490,
         round_inst_S_15__sbox_inst_com_y_inst_n489,
         round_inst_S_15__sbox_inst_com_y_inst_n488,
         round_inst_S_15__sbox_inst_com_y_inst_n487,
         round_inst_S_15__sbox_inst_com_y_inst_n486,
         round_inst_S_15__sbox_inst_com_y_inst_n485,
         round_inst_S_15__sbox_inst_com_y_inst_n484,
         round_inst_S_15__sbox_inst_com_y_inst_n483,
         round_inst_S_15__sbox_inst_com_y_inst_n482,
         round_inst_S_15__sbox_inst_com_y_inst_n481,
         round_inst_S_15__sbox_inst_com_y_inst_n480,
         round_inst_S_15__sbox_inst_com_y_inst_n479,
         round_inst_S_15__sbox_inst_com_y_inst_n478,
         round_inst_S_15__sbox_inst_com_y_inst_n477,
         round_inst_S_15__sbox_inst_com_y_inst_n476,
         round_inst_S_15__sbox_inst_com_y_inst_n475,
         round_inst_S_15__sbox_inst_com_y_inst_n474,
         round_inst_S_15__sbox_inst_com_y_inst_n473,
         round_inst_S_15__sbox_inst_com_y_inst_n472,
         round_inst_S_15__sbox_inst_com_y_inst_n471,
         round_inst_S_15__sbox_inst_com_y_inst_n470,
         round_inst_S_15__sbox_inst_com_y_inst_n469,
         round_inst_S_15__sbox_inst_com_y_inst_n468,
         round_inst_S_15__sbox_inst_com_y_inst_n467,
         round_inst_S_15__sbox_inst_com_y_inst_n466,
         round_inst_S_15__sbox_inst_com_y_inst_n465,
         round_inst_S_15__sbox_inst_com_y_inst_n464,
         round_inst_S_15__sbox_inst_com_y_inst_n463,
         round_inst_S_15__sbox_inst_com_y_inst_n462,
         round_inst_S_15__sbox_inst_com_y_inst_n461,
         round_inst_S_15__sbox_inst_com_y_inst_n460,
         round_inst_S_15__sbox_inst_com_y_inst_n459,
         round_inst_S_15__sbox_inst_com_y_inst_n458,
         round_inst_S_15__sbox_inst_com_y_inst_n457,
         round_inst_S_15__sbox_inst_com_y_inst_n456,
         round_inst_S_15__sbox_inst_com_y_inst_n455,
         round_inst_S_15__sbox_inst_com_y_inst_n454,
         round_inst_S_15__sbox_inst_com_y_inst_n453,
         round_inst_S_15__sbox_inst_com_y_inst_n452,
         round_inst_S_15__sbox_inst_com_y_inst_n451,
         round_inst_S_15__sbox_inst_com_y_inst_n450,
         round_inst_S_15__sbox_inst_com_y_inst_n449,
         round_inst_S_15__sbox_inst_com_y_inst_n448,
         round_inst_S_15__sbox_inst_com_y_inst_n447,
         round_inst_S_15__sbox_inst_com_y_inst_n446,
         round_inst_S_15__sbox_inst_com_y_inst_n445,
         round_inst_S_15__sbox_inst_com_y_inst_n444,
         round_inst_S_15__sbox_inst_com_y_inst_n443,
         round_inst_S_15__sbox_inst_com_y_inst_n442,
         round_inst_S_15__sbox_inst_com_y_inst_n441,
         round_inst_S_15__sbox_inst_com_y_inst_n440,
         round_inst_S_15__sbox_inst_com_y_inst_n439,
         round_inst_S_15__sbox_inst_com_y_inst_n438,
         round_inst_S_15__sbox_inst_com_y_inst_n437,
         round_inst_S_15__sbox_inst_com_y_inst_n436,
         round_inst_S_15__sbox_inst_com_y_inst_n435,
         round_inst_S_15__sbox_inst_com_y_inst_n434,
         round_inst_S_15__sbox_inst_com_y_inst_n433,
         round_inst_S_15__sbox_inst_com_y_inst_n432,
         round_inst_S_15__sbox_inst_com_y_inst_n431,
         round_inst_S_15__sbox_inst_com_y_inst_n430,
         round_inst_S_15__sbox_inst_com_y_inst_n429,
         round_inst_S_15__sbox_inst_com_y_inst_n428,
         round_inst_S_15__sbox_inst_com_y_inst_n427,
         round_inst_S_15__sbox_inst_com_y_inst_n426,
         round_inst_S_15__sbox_inst_com_y_inst_n425,
         round_inst_S_15__sbox_inst_com_y_inst_n424,
         round_inst_S_15__sbox_inst_com_y_inst_n423,
         round_inst_S_15__sbox_inst_com_y_inst_n422,
         round_inst_S_15__sbox_inst_com_y_inst_n421,
         round_inst_S_15__sbox_inst_com_y_inst_n420,
         round_inst_S_15__sbox_inst_com_y_inst_n419,
         round_inst_S_15__sbox_inst_com_y_inst_n418,
         round_inst_S_15__sbox_inst_com_y_inst_n417,
         round_inst_S_15__sbox_inst_com_y_inst_n416,
         round_inst_S_15__sbox_inst_com_y_inst_n415,
         round_inst_S_15__sbox_inst_com_y_inst_n414,
         round_inst_S_15__sbox_inst_com_y_inst_n413,
         round_inst_S_15__sbox_inst_com_y_inst_n412,
         round_inst_S_15__sbox_inst_com_y_inst_n411,
         round_inst_S_15__sbox_inst_com_y_inst_n410,
         round_inst_S_15__sbox_inst_com_y_inst_n409,
         round_inst_S_15__sbox_inst_com_y_inst_n408,
         round_inst_S_15__sbox_inst_com_y_inst_n407,
         round_inst_S_15__sbox_inst_com_y_inst_n406,
         round_inst_S_15__sbox_inst_com_y_inst_n405,
         round_inst_S_15__sbox_inst_com_y_inst_n404,
         round_inst_S_15__sbox_inst_com_y_inst_n403,
         round_inst_S_15__sbox_inst_com_y_inst_n402,
         round_inst_S_15__sbox_inst_com_y_inst_n401,
         round_inst_S_15__sbox_inst_com_y_inst_n400,
         round_inst_S_15__sbox_inst_com_y_inst_n399,
         round_inst_S_15__sbox_inst_com_y_inst_n398,
         round_inst_S_15__sbox_inst_com_y_inst_n397,
         round_inst_S_15__sbox_inst_com_y_inst_n396,
         round_inst_S_15__sbox_inst_com_y_inst_n395,
         round_inst_S_15__sbox_inst_com_y_inst_n394,
         round_inst_S_15__sbox_inst_com_y_inst_n393,
         round_inst_S_15__sbox_inst_com_y_inst_n392,
         round_inst_S_15__sbox_inst_com_y_inst_n391,
         round_inst_S_15__sbox_inst_com_y_inst_n390,
         round_inst_S_15__sbox_inst_com_y_inst_n389,
         round_inst_S_15__sbox_inst_com_y_inst_n388,
         round_inst_S_15__sbox_inst_com_y_inst_n387,
         round_inst_S_15__sbox_inst_com_y_inst_n386,
         round_inst_S_15__sbox_inst_com_z_inst_n517,
         round_inst_S_15__sbox_inst_com_z_inst_n516,
         round_inst_S_15__sbox_inst_com_z_inst_n515,
         round_inst_S_15__sbox_inst_com_z_inst_n514,
         round_inst_S_15__sbox_inst_com_z_inst_n513,
         round_inst_S_15__sbox_inst_com_z_inst_n512,
         round_inst_S_15__sbox_inst_com_z_inst_n511,
         round_inst_S_15__sbox_inst_com_z_inst_n510,
         round_inst_S_15__sbox_inst_com_z_inst_n509,
         round_inst_S_15__sbox_inst_com_z_inst_n508,
         round_inst_S_15__sbox_inst_com_z_inst_n507,
         round_inst_S_15__sbox_inst_com_z_inst_n506,
         round_inst_S_15__sbox_inst_com_z_inst_n505,
         round_inst_S_15__sbox_inst_com_z_inst_n504,
         round_inst_S_15__sbox_inst_com_z_inst_n503,
         round_inst_S_15__sbox_inst_com_z_inst_n502,
         round_inst_S_15__sbox_inst_com_z_inst_n501,
         round_inst_S_15__sbox_inst_com_z_inst_n500,
         round_inst_S_15__sbox_inst_com_z_inst_n499,
         round_inst_S_15__sbox_inst_com_z_inst_n498,
         round_inst_S_15__sbox_inst_com_z_inst_n497,
         round_inst_S_15__sbox_inst_com_z_inst_n496,
         round_inst_S_15__sbox_inst_com_z_inst_n495,
         round_inst_S_15__sbox_inst_com_z_inst_n494,
         round_inst_S_15__sbox_inst_com_z_inst_n493,
         round_inst_S_15__sbox_inst_com_z_inst_n492,
         round_inst_S_15__sbox_inst_com_z_inst_n491,
         round_inst_S_15__sbox_inst_com_z_inst_n490,
         round_inst_S_15__sbox_inst_com_z_inst_n489,
         round_inst_S_15__sbox_inst_com_z_inst_n488,
         round_inst_S_15__sbox_inst_com_z_inst_n487,
         round_inst_S_15__sbox_inst_com_z_inst_n486,
         round_inst_S_15__sbox_inst_com_z_inst_n485,
         round_inst_S_15__sbox_inst_com_z_inst_n484,
         round_inst_S_15__sbox_inst_com_z_inst_n483,
         round_inst_S_15__sbox_inst_com_z_inst_n482,
         round_inst_S_15__sbox_inst_com_z_inst_n481,
         round_inst_S_15__sbox_inst_com_z_inst_n480,
         round_inst_S_15__sbox_inst_com_z_inst_n479,
         round_inst_S_15__sbox_inst_com_z_inst_n478,
         round_inst_S_15__sbox_inst_com_z_inst_n477,
         round_inst_S_15__sbox_inst_com_z_inst_n476,
         round_inst_S_15__sbox_inst_com_z_inst_n475,
         round_inst_S_15__sbox_inst_com_z_inst_n474,
         round_inst_S_15__sbox_inst_com_z_inst_n473,
         round_inst_S_15__sbox_inst_com_z_inst_n472,
         round_inst_S_15__sbox_inst_com_z_inst_n471,
         round_inst_S_15__sbox_inst_com_z_inst_n470,
         round_inst_S_15__sbox_inst_com_z_inst_n469,
         round_inst_S_15__sbox_inst_com_z_inst_n468,
         round_inst_S_15__sbox_inst_com_z_inst_n467,
         round_inst_S_15__sbox_inst_com_z_inst_n466,
         round_inst_S_15__sbox_inst_com_z_inst_n465,
         round_inst_S_15__sbox_inst_com_z_inst_n464,
         round_inst_S_15__sbox_inst_com_z_inst_n463,
         round_inst_S_15__sbox_inst_com_z_inst_n462,
         round_inst_S_15__sbox_inst_com_z_inst_n461,
         round_inst_S_15__sbox_inst_com_z_inst_n460,
         round_inst_S_15__sbox_inst_com_z_inst_n459,
         round_inst_S_15__sbox_inst_com_z_inst_n458,
         round_inst_S_15__sbox_inst_com_z_inst_n457,
         round_inst_S_15__sbox_inst_com_z_inst_n456,
         round_inst_S_15__sbox_inst_com_z_inst_n455,
         round_inst_S_15__sbox_inst_com_z_inst_n454,
         round_inst_S_15__sbox_inst_com_z_inst_n453,
         round_inst_S_15__sbox_inst_com_z_inst_n452,
         round_inst_S_15__sbox_inst_com_z_inst_n451,
         round_inst_S_15__sbox_inst_com_z_inst_n450,
         round_inst_S_15__sbox_inst_com_z_inst_n449,
         round_inst_S_15__sbox_inst_com_z_inst_n448,
         round_inst_S_15__sbox_inst_com_z_inst_n447,
         round_inst_S_15__sbox_inst_com_z_inst_n446,
         round_inst_S_15__sbox_inst_com_z_inst_n445,
         round_inst_S_15__sbox_inst_com_z_inst_n444,
         round_inst_S_15__sbox_inst_com_z_inst_n443,
         round_inst_S_15__sbox_inst_com_z_inst_n442,
         round_inst_S_15__sbox_inst_com_z_inst_n441,
         round_inst_S_15__sbox_inst_com_z_inst_n440,
         round_inst_S_15__sbox_inst_com_z_inst_n439,
         round_inst_S_15__sbox_inst_com_z_inst_n438,
         round_inst_S_15__sbox_inst_com_z_inst_n437,
         round_inst_S_15__sbox_inst_com_z_inst_n436,
         round_inst_S_15__sbox_inst_com_z_inst_n435,
         round_inst_S_15__sbox_inst_com_z_inst_n434,
         round_inst_S_15__sbox_inst_com_z_inst_n433,
         round_inst_S_15__sbox_inst_com_z_inst_n432,
         round_inst_S_15__sbox_inst_com_z_inst_n431,
         round_inst_S_15__sbox_inst_com_z_inst_n430,
         round_inst_S_15__sbox_inst_com_z_inst_n429,
         round_inst_S_15__sbox_inst_com_z_inst_n428,
         round_inst_S_15__sbox_inst_com_z_inst_n427,
         round_inst_S_15__sbox_inst_com_z_inst_n426,
         round_inst_S_15__sbox_inst_com_z_inst_n425,
         round_inst_S_15__sbox_inst_com_z_inst_n424,
         round_inst_S_15__sbox_inst_com_z_inst_n423,
         round_inst_S_15__sbox_inst_com_z_inst_n422,
         round_inst_S_15__sbox_inst_com_z_inst_n421,
         round_inst_S_15__sbox_inst_com_z_inst_n420,
         round_inst_S_15__sbox_inst_com_z_inst_n419,
         round_inst_S_15__sbox_inst_com_z_inst_n418,
         round_inst_S_15__sbox_inst_com_z_inst_n417,
         round_inst_S_15__sbox_inst_com_z_inst_n416,
         round_inst_S_15__sbox_inst_com_z_inst_n415,
         round_inst_S_15__sbox_inst_com_z_inst_n414,
         round_inst_S_15__sbox_inst_com_z_inst_n413,
         round_inst_S_15__sbox_inst_com_z_inst_n412,
         round_inst_S_15__sbox_inst_com_z_inst_n411,
         round_inst_S_15__sbox_inst_com_z_inst_n410,
         round_inst_S_15__sbox_inst_com_z_inst_n409,
         round_inst_S_15__sbox_inst_com_z_inst_n408,
         round_inst_S_15__sbox_inst_com_z_inst_n407,
         round_inst_S_15__sbox_inst_com_z_inst_n406,
         round_inst_S_15__sbox_inst_com_z_inst_n405,
         round_inst_S_15__sbox_inst_com_z_inst_n404,
         round_inst_S_15__sbox_inst_com_z_inst_n403,
         round_inst_S_15__sbox_inst_com_z_inst_n402,
         round_inst_S_15__sbox_inst_com_z_inst_n401,
         round_inst_S_15__sbox_inst_com_z_inst_n400,
         round_inst_S_15__sbox_inst_com_z_inst_n399,
         round_inst_S_15__sbox_inst_com_z_inst_n398,
         round_inst_S_15__sbox_inst_com_z_inst_n397,
         round_inst_S_15__sbox_inst_com_z_inst_n396,
         round_inst_S_15__sbox_inst_com_z_inst_n395,
         round_inst_S_15__sbox_inst_com_z_inst_n394,
         round_inst_S_15__sbox_inst_com_z_inst_n393,
         round_inst_S_15__sbox_inst_com_z_inst_n392,
         round_inst_S_15__sbox_inst_com_z_inst_n391,
         round_inst_S_15__sbox_inst_com_z_inst_n390, round_inst_A2_0__aw2_n5,
         round_inst_A2_0__ax2_n3, round_inst_A2_0__ay2_n3,
         round_inst_A2_0__az2_n3, round_inst_A2_1__aw2_n5,
         round_inst_A2_1__ax2_n3, round_inst_A2_1__ay2_n3,
         round_inst_A2_1__az2_n3, round_inst_A2_2__aw2_n5,
         round_inst_A2_2__ax2_n3, round_inst_A2_2__ay2_n3,
         round_inst_A2_2__az2_n3, round_inst_A2_3__aw2_n5,
         round_inst_A2_3__ax2_n3, round_inst_A2_3__ay2_n3,
         round_inst_A2_3__az2_n3, round_inst_A2_4__aw2_n5,
         round_inst_A2_4__ax2_n3, round_inst_A2_4__ay2_n3,
         round_inst_A2_4__az2_n3, round_inst_A2_5__aw2_n5,
         round_inst_A2_5__ax2_n3, round_inst_A2_5__ay2_n3,
         round_inst_A2_5__az2_n3, round_inst_A2_6__aw2_n5,
         round_inst_A2_6__ax2_n3, round_inst_A2_6__ay2_n3,
         round_inst_A2_6__az2_n3, round_inst_A2_7__aw2_n5,
         round_inst_A2_7__ax2_n3, round_inst_A2_7__ay2_n3,
         round_inst_A2_7__az2_n3, round_inst_A2_8__aw2_n5,
         round_inst_A2_8__ax2_n3, round_inst_A2_8__ay2_n3,
         round_inst_A2_8__az2_n3, round_inst_A2_9__aw2_n5,
         round_inst_A2_9__ax2_n3, round_inst_A2_9__ay2_n3,
         round_inst_A2_9__az2_n3, round_inst_A2_10__aw2_n5,
         round_inst_A2_10__ax2_n3, round_inst_A2_10__ay2_n3,
         round_inst_A2_10__az2_n3, round_inst_A2_11__aw2_n5,
         round_inst_A2_11__ax2_n3, round_inst_A2_11__ay2_n3,
         round_inst_A2_11__az2_n3, round_inst_A2_12__aw2_n5,
         round_inst_A2_12__ax2_n3, round_inst_A2_12__ay2_n3,
         round_inst_A2_12__az2_n3, round_inst_A2_13__aw2_n5,
         round_inst_A2_13__ax2_n3, round_inst_A2_13__ay2_n3,
         round_inst_A2_13__az2_n3, round_inst_A2_14__aw2_n5,
         round_inst_A2_14__ax2_n3, round_inst_A2_14__ay2_n3,
         round_inst_A2_14__az2_n3, round_inst_A2_15__aw2_n5,
         round_inst_A2_15__ax2_n3, round_inst_A2_15__ay2_n3,
         round_inst_A2_15__az2_n3, round_inst_mux_inv_w2_n266,
         round_inst_mux_inv_w2_n265, round_inst_mux_inv_w2_n264,
         round_inst_mux_inv_w2_n263, round_inst_mux_inv_x2_n267,
         round_inst_mux_inv_x2_n266, round_inst_mux_inv_x2_n265,
         round_inst_mux_inv_x2_n264, round_inst_mux_inv_x2_n263,
         round_inst_mux_inv_y2_n267, round_inst_mux_inv_y2_n266,
         round_inst_mux_inv_y2_n265, round_inst_mux_inv_y2_n264,
         round_inst_mux_inv_y2_n263, round_inst_mux_inv_z2_n267,
         round_inst_mux_inv_z2_n266, round_inst_mux_inv_z2_n265,
         round_inst_mux_inv_z2_n264, round_inst_mux_inv_z2_n263,
         round_inst_mw_inst_n32, round_inst_mw_inst_n31,
         round_inst_mw_inst_n30, round_inst_mw_inst_n29,
         round_inst_mw_inst_n28, round_inst_mw_inst_n27,
         round_inst_mw_inst_n26, round_inst_mw_inst_n25,
         round_inst_mw_inst_n24, round_inst_mw_inst_n23,
         round_inst_mw_inst_n22, round_inst_mw_inst_n21,
         round_inst_mw_inst_n20, round_inst_mw_inst_n19,
         round_inst_mw_inst_n18, round_inst_mw_inst_n17,
         round_inst_mw_inst_n16, round_inst_mw_inst_n15,
         round_inst_mw_inst_n14, round_inst_mw_inst_n13,
         round_inst_mw_inst_n12, round_inst_mw_inst_n11,
         round_inst_mw_inst_n10, round_inst_mw_inst_n9, round_inst_mw_inst_n8,
         round_inst_mw_inst_n7, round_inst_mw_inst_n6, round_inst_mw_inst_n5,
         round_inst_mw_inst_n4, round_inst_mw_inst_n3, round_inst_mw_inst_n2,
         round_inst_mw_inst_n1, round_inst_mx_inst_n96, round_inst_mx_inst_n95,
         round_inst_mx_inst_n94, round_inst_mx_inst_n93,
         round_inst_mx_inst_n92, round_inst_mx_inst_n91,
         round_inst_mx_inst_n90, round_inst_mx_inst_n89,
         round_inst_mx_inst_n88, round_inst_mx_inst_n87,
         round_inst_mx_inst_n86, round_inst_mx_inst_n85,
         round_inst_mx_inst_n84, round_inst_mx_inst_n83,
         round_inst_mx_inst_n82, round_inst_mx_inst_n81,
         round_inst_mx_inst_n80, round_inst_mx_inst_n79,
         round_inst_mx_inst_n78, round_inst_mx_inst_n77,
         round_inst_mx_inst_n76, round_inst_mx_inst_n75,
         round_inst_mx_inst_n74, round_inst_mx_inst_n73,
         round_inst_mx_inst_n72, round_inst_mx_inst_n71,
         round_inst_mx_inst_n70, round_inst_mx_inst_n69,
         round_inst_mx_inst_n68, round_inst_mx_inst_n67,
         round_inst_mx_inst_n66, round_inst_mx_inst_n65,
         round_inst_my_inst_n96, round_inst_my_inst_n95,
         round_inst_my_inst_n94, round_inst_my_inst_n93,
         round_inst_my_inst_n92, round_inst_my_inst_n91,
         round_inst_my_inst_n90, round_inst_my_inst_n89,
         round_inst_my_inst_n88, round_inst_my_inst_n87,
         round_inst_my_inst_n86, round_inst_my_inst_n85,
         round_inst_my_inst_n84, round_inst_my_inst_n83,
         round_inst_my_inst_n82, round_inst_my_inst_n81,
         round_inst_my_inst_n80, round_inst_my_inst_n79,
         round_inst_my_inst_n78, round_inst_my_inst_n77,
         round_inst_my_inst_n76, round_inst_my_inst_n75,
         round_inst_my_inst_n74, round_inst_my_inst_n73,
         round_inst_my_inst_n72, round_inst_my_inst_n71,
         round_inst_my_inst_n70, round_inst_my_inst_n69,
         round_inst_my_inst_n68, round_inst_my_inst_n67,
         round_inst_my_inst_n66, round_inst_my_inst_n65,
         round_inst_mz_inst_n96, round_inst_mz_inst_n95,
         round_inst_mz_inst_n94, round_inst_mz_inst_n93,
         round_inst_mz_inst_n92, round_inst_mz_inst_n91,
         round_inst_mz_inst_n90, round_inst_mz_inst_n89,
         round_inst_mz_inst_n88, round_inst_mz_inst_n87,
         round_inst_mz_inst_n86, round_inst_mz_inst_n85,
         round_inst_mz_inst_n84, round_inst_mz_inst_n83,
         round_inst_mz_inst_n82, round_inst_mz_inst_n81,
         round_inst_mz_inst_n80, round_inst_mz_inst_n79,
         round_inst_mz_inst_n78, round_inst_mz_inst_n77,
         round_inst_mz_inst_n76, round_inst_mz_inst_n75,
         round_inst_mz_inst_n74, round_inst_mz_inst_n73,
         round_inst_mz_inst_n72, round_inst_mz_inst_n71,
         round_inst_mz_inst_n70, round_inst_mz_inst_n69,
         round_inst_mz_inst_n68, round_inst_mz_inst_n67,
         round_inst_mz_inst_n66, round_inst_mz_inst_n65, mux_c0_n265,
         mux_c0_n264, mux_c0_n263, mux_c1_n265, mux_c1_n264, mux_c1_n263,
         mux_c2_n264, mux_c2_n263, mux_c3_n264, mux_c3_n263, mux_c3_n262;
  wire   [63:0] init_w;
  wire   [63:0] rout_w;
  wire   [63:0] state_w;
  wire   [63:0] rout_x;
  wire   [63:0] state_x;
  wire   [63:0] rout_y;
  wire   [63:0] state_y;
  wire   [63:0] rout_z;
  wire   [63:0] state_z;
  wire   [3:0] bout;
  wire   [3:0] state_b;
  wire   [3:0] cout;
  wire   [3:0] state_c;
  wire   [3:0] dout;
  wire   [3:0] state_d;
  wire   [3:0] bin;
  wire   [3:0] cin;
  wire   [3:0] din;
  wire   [63:0] final_w_k;
  wire   [2:0] cntrl_inst_counter;
  wire   [63:0] round_inst_min_z;
  wire   [63:0] round_inst_min_y;
  wire   [63:0] round_inst_min_x;
  wire   [63:0] round_inst_min_w;
  wire   [63:0] round_inst_srout2_z;
  wire   [63:0] round_inst_srout2_y;
  wire   [63:0] round_inst_srout2_x;
  wire   [63:0] round_inst_srout2_w;
  wire   [63:0] round_inst_xin_w;
  wire   [60:0] round_inst_sout_z;
  wire   [60:0] round_inst_sout_y;
  wire   [60:0] round_inst_sout_x;
  wire   [63:0] round_inst_sout_w;
  wire   [59:0] round_inst_sin_z;
  wire   [59:0] round_inst_sin_y;
  wire   [59:0] round_inst_sin_x;
  wire   [63:0] round_inst_sin_w;
  wire   [63:0] round_inst_aout_z;
  wire   [63:0] round_inst_aout_y;
  wire   [63:0] round_inst_aout_x;
  wire   [63:0] round_inst_aout_w;
  wire   [63:0] round_inst_xout_w;
  wire   [60:0] round_inst_srout_z;
  wire   [60:0] round_inst_srout_y;
  wire   [60:0] round_inst_srout_x;
  wire   [63:0] round_inst_srout_w;

  MUX2_X1 U773 ( .A(k[74]), .B(k[73]), .S(enc), .Z(n526) );
  XOR2_X1 U774 ( .A(p0[9]), .B(n526), .Z(init_w[57]) );
  MUX2_X1 U775 ( .A(k[73]), .B(k[72]), .S(enc), .Z(n527) );
  XOR2_X1 U776 ( .A(p0[8]), .B(n527), .Z(init_w[56]) );
  MUX2_X1 U777 ( .A(k[72]), .B(k[71]), .S(enc), .Z(n528) );
  XOR2_X1 U778 ( .A(p0[7]), .B(n528), .Z(init_w[39]) );
  MUX2_X1 U779 ( .A(k[71]), .B(k[70]), .S(enc), .Z(n529) );
  XOR2_X1 U780 ( .A(p0[6]), .B(n529), .Z(init_w[38]) );
  MUX2_X1 U781 ( .A(k[64]), .B(k[127]), .S(enc), .Z(n530) );
  XOR2_X1 U782 ( .A(p0[63]), .B(n530), .Z(init_w[63]) );
  MUX2_X1 U783 ( .A(k[127]), .B(k[126]), .S(enc), .Z(n531) );
  XOR2_X1 U784 ( .A(p0[62]), .B(n531), .Z(init_w[62]) );
  MUX2_X1 U785 ( .A(k[126]), .B(k[125]), .S(enc), .Z(n532) );
  XOR2_X1 U786 ( .A(p0[61]), .B(n532), .Z(init_w[61]) );
  MUX2_X1 U787 ( .A(k[125]), .B(k[124]), .S(enc), .Z(n533) );
  XOR2_X1 U788 ( .A(p0[60]), .B(n533), .Z(init_w[60]) );
  MUX2_X1 U789 ( .A(k[70]), .B(k[69]), .S(enc), .Z(n534) );
  XOR2_X1 U790 ( .A(p0[5]), .B(n534), .Z(init_w[37]) );
  MUX2_X1 U791 ( .A(k[124]), .B(k[123]), .S(enc), .Z(n535) );
  XOR2_X1 U792 ( .A(p0[59]), .B(n535), .Z(init_w[43]) );
  MUX2_X1 U793 ( .A(k[123]), .B(k[122]), .S(enc), .Z(n536) );
  XOR2_X1 U794 ( .A(p0[58]), .B(n536), .Z(init_w[42]) );
  MUX2_X1 U795 ( .A(k[122]), .B(k[121]), .S(enc), .Z(n537) );
  XOR2_X1 U796 ( .A(p0[57]), .B(n537), .Z(init_w[41]) );
  MUX2_X1 U797 ( .A(k[121]), .B(k[120]), .S(enc), .Z(n538) );
  XOR2_X1 U798 ( .A(p0[56]), .B(n538), .Z(init_w[40]) );
  MUX2_X1 U799 ( .A(k[120]), .B(k[119]), .S(enc), .Z(n539) );
  XOR2_X1 U800 ( .A(p0[55]), .B(n539), .Z(init_w[23]) );
  MUX2_X1 U801 ( .A(k[119]), .B(k[118]), .S(enc), .Z(n540) );
  XOR2_X1 U802 ( .A(p0[54]), .B(n540), .Z(init_w[22]) );
  MUX2_X1 U803 ( .A(k[118]), .B(k[117]), .S(enc), .Z(n541) );
  XOR2_X1 U804 ( .A(p0[53]), .B(n541), .Z(init_w[21]) );
  MUX2_X1 U805 ( .A(k[117]), .B(k[116]), .S(enc), .Z(n542) );
  XOR2_X1 U806 ( .A(p0[52]), .B(n542), .Z(init_w[20]) );
  MUX2_X1 U807 ( .A(k[116]), .B(k[115]), .S(enc), .Z(n543) );
  XOR2_X1 U808 ( .A(p0[51]), .B(n543), .Z(init_w[3]) );
  MUX2_X1 U809 ( .A(k[115]), .B(k[114]), .S(enc), .Z(n544) );
  XOR2_X1 U810 ( .A(p0[50]), .B(n544), .Z(init_w[2]) );
  MUX2_X1 U811 ( .A(k[69]), .B(k[68]), .S(enc), .Z(n545) );
  XOR2_X1 U812 ( .A(p0[4]), .B(n545), .Z(init_w[36]) );
  MUX2_X1 U813 ( .A(k[114]), .B(k[113]), .S(enc), .Z(n546) );
  XOR2_X1 U814 ( .A(p0[49]), .B(n546), .Z(init_w[1]) );
  MUX2_X1 U815 ( .A(k[113]), .B(k[112]), .S(enc), .Z(n547) );
  XOR2_X1 U816 ( .A(p0[48]), .B(n547), .Z(init_w[0]) );
  MUX2_X1 U817 ( .A(k[112]), .B(k[111]), .S(enc), .Z(n548) );
  XOR2_X1 U818 ( .A(p0[47]), .B(n548), .Z(init_w[47]) );
  MUX2_X1 U819 ( .A(k[111]), .B(k[110]), .S(enc), .Z(n549) );
  XOR2_X1 U820 ( .A(p0[46]), .B(n549), .Z(init_w[46]) );
  MUX2_X1 U821 ( .A(k[110]), .B(k[109]), .S(enc), .Z(n550) );
  XOR2_X1 U822 ( .A(p0[45]), .B(n550), .Z(init_w[45]) );
  MUX2_X1 U823 ( .A(k[109]), .B(k[108]), .S(enc), .Z(n551) );
  XOR2_X1 U824 ( .A(p0[44]), .B(n551), .Z(init_w[44]) );
  MUX2_X1 U825 ( .A(k[108]), .B(k[107]), .S(enc), .Z(n552) );
  XOR2_X1 U826 ( .A(p0[43]), .B(n552), .Z(init_w[27]) );
  MUX2_X1 U827 ( .A(k[107]), .B(k[106]), .S(enc), .Z(n553) );
  XOR2_X1 U828 ( .A(p0[42]), .B(n553), .Z(init_w[26]) );
  MUX2_X1 U829 ( .A(k[106]), .B(k[105]), .S(enc), .Z(n554) );
  XOR2_X1 U830 ( .A(p0[41]), .B(n554), .Z(init_w[25]) );
  MUX2_X1 U831 ( .A(k[105]), .B(k[104]), .S(enc), .Z(n555) );
  XOR2_X1 U832 ( .A(p0[40]), .B(n555), .Z(init_w[24]) );
  MUX2_X1 U833 ( .A(k[68]), .B(k[67]), .S(enc), .Z(n556) );
  XOR2_X1 U834 ( .A(p0[3]), .B(n556), .Z(init_w[19]) );
  MUX2_X1 U835 ( .A(k[104]), .B(k[103]), .S(enc), .Z(n557) );
  XOR2_X1 U836 ( .A(p0[39]), .B(n557), .Z(init_w[7]) );
  MUX2_X1 U837 ( .A(k[103]), .B(k[102]), .S(enc), .Z(n558) );
  XOR2_X1 U838 ( .A(p0[38]), .B(n558), .Z(init_w[6]) );
  MUX2_X1 U839 ( .A(k[102]), .B(k[101]), .S(enc), .Z(n559) );
  XOR2_X1 U840 ( .A(p0[37]), .B(n559), .Z(init_w[5]) );
  MUX2_X1 U841 ( .A(k[101]), .B(k[100]), .S(enc), .Z(n560) );
  XOR2_X1 U842 ( .A(p0[36]), .B(n560), .Z(init_w[4]) );
  MUX2_X1 U843 ( .A(k[100]), .B(k[99]), .S(enc), .Z(n561) );
  XOR2_X1 U844 ( .A(p0[35]), .B(n561), .Z(init_w[51]) );
  MUX2_X1 U845 ( .A(k[99]), .B(k[98]), .S(enc), .Z(n562) );
  XOR2_X1 U846 ( .A(p0[34]), .B(n562), .Z(init_w[50]) );
  MUX2_X1 U847 ( .A(k[98]), .B(k[97]), .S(enc), .Z(n563) );
  XOR2_X1 U848 ( .A(p0[33]), .B(n563), .Z(init_w[49]) );
  MUX2_X1 U849 ( .A(k[97]), .B(k[96]), .S(enc), .Z(n564) );
  XOR2_X1 U850 ( .A(p0[32]), .B(n564), .Z(init_w[48]) );
  MUX2_X1 U851 ( .A(k[96]), .B(k[95]), .S(enc), .Z(n565) );
  XOR2_X1 U852 ( .A(p0[31]), .B(n565), .Z(init_w[31]) );
  MUX2_X1 U853 ( .A(k[95]), .B(k[94]), .S(enc), .Z(n566) );
  XOR2_X1 U854 ( .A(p0[30]), .B(n566), .Z(init_w[30]) );
  MUX2_X1 U855 ( .A(k[67]), .B(k[66]), .S(enc), .Z(n567) );
  XOR2_X1 U856 ( .A(p0[2]), .B(n567), .Z(init_w[18]) );
  MUX2_X1 U857 ( .A(k[94]), .B(k[93]), .S(enc), .Z(n568) );
  XOR2_X1 U858 ( .A(p0[29]), .B(n568), .Z(init_w[29]) );
  MUX2_X1 U859 ( .A(k[93]), .B(k[92]), .S(enc), .Z(n569) );
  XOR2_X1 U860 ( .A(p0[28]), .B(n569), .Z(init_w[28]) );
  MUX2_X1 U861 ( .A(k[92]), .B(k[91]), .S(enc), .Z(n570) );
  XOR2_X1 U862 ( .A(p0[27]), .B(n570), .Z(init_w[11]) );
  MUX2_X1 U863 ( .A(k[91]), .B(k[90]), .S(enc), .Z(n571) );
  XOR2_X1 U864 ( .A(p0[26]), .B(n571), .Z(init_w[10]) );
  MUX2_X1 U865 ( .A(k[90]), .B(k[89]), .S(enc), .Z(n572) );
  XOR2_X1 U866 ( .A(p0[25]), .B(n572), .Z(init_w[9]) );
  MUX2_X1 U867 ( .A(k[89]), .B(k[88]), .S(enc), .Z(n573) );
  XOR2_X1 U868 ( .A(p0[24]), .B(n573), .Z(init_w[8]) );
  MUX2_X1 U869 ( .A(k[88]), .B(k[87]), .S(enc), .Z(n574) );
  XOR2_X1 U870 ( .A(p0[23]), .B(n574), .Z(init_w[55]) );
  MUX2_X1 U871 ( .A(k[87]), .B(k[86]), .S(enc), .Z(n575) );
  XOR2_X1 U872 ( .A(p0[22]), .B(n575), .Z(init_w[54]) );
  MUX2_X1 U873 ( .A(k[86]), .B(k[85]), .S(enc), .Z(n576) );
  XOR2_X1 U874 ( .A(p0[21]), .B(n576), .Z(init_w[53]) );
  MUX2_X1 U875 ( .A(k[85]), .B(k[84]), .S(enc), .Z(n577) );
  XOR2_X1 U876 ( .A(p0[20]), .B(n577), .Z(init_w[52]) );
  MUX2_X1 U877 ( .A(k[66]), .B(k[65]), .S(enc), .Z(n578) );
  XOR2_X1 U878 ( .A(p0[1]), .B(n578), .Z(init_w[17]) );
  MUX2_X1 U879 ( .A(k[84]), .B(k[83]), .S(enc), .Z(n579) );
  XOR2_X1 U880 ( .A(p0[19]), .B(n579), .Z(init_w[35]) );
  MUX2_X1 U881 ( .A(k[83]), .B(k[82]), .S(enc), .Z(n580) );
  XOR2_X1 U882 ( .A(p0[18]), .B(n580), .Z(init_w[34]) );
  MUX2_X1 U883 ( .A(k[82]), .B(k[81]), .S(enc), .Z(n581) );
  XOR2_X1 U884 ( .A(p0[17]), .B(n581), .Z(init_w[33]) );
  MUX2_X1 U885 ( .A(k[81]), .B(k[80]), .S(enc), .Z(n582) );
  XOR2_X1 U886 ( .A(p0[16]), .B(n582), .Z(init_w[32]) );
  MUX2_X1 U887 ( .A(k[80]), .B(k[79]), .S(enc), .Z(n583) );
  XOR2_X1 U888 ( .A(p0[15]), .B(n583), .Z(init_w[15]) );
  MUX2_X1 U889 ( .A(k[79]), .B(k[78]), .S(enc), .Z(n584) );
  XOR2_X1 U890 ( .A(p0[14]), .B(n584), .Z(init_w[14]) );
  MUX2_X1 U891 ( .A(k[78]), .B(k[77]), .S(enc), .Z(n585) );
  XOR2_X1 U892 ( .A(p0[13]), .B(n585), .Z(init_w[13]) );
  MUX2_X1 U893 ( .A(k[77]), .B(k[76]), .S(enc), .Z(n586) );
  XOR2_X1 U894 ( .A(p0[12]), .B(n586), .Z(init_w[12]) );
  MUX2_X1 U895 ( .A(k[76]), .B(k[75]), .S(enc), .Z(n587) );
  XOR2_X1 U896 ( .A(p0[11]), .B(n587), .Z(init_w[59]) );
  MUX2_X1 U897 ( .A(k[75]), .B(k[74]), .S(enc), .Z(n588) );
  XOR2_X1 U898 ( .A(p0[10]), .B(n588), .Z(init_w[58]) );
  MUX2_X1 U899 ( .A(kext_64_), .B(k[64]), .S(enc), .Z(n589) );
  XOR2_X1 U900 ( .A(p0[0]), .B(n589), .Z(init_w[16]) );
  MUX2_X1 U901 ( .A(k[73]), .B(k[74]), .S(enc), .Z(n590) );
  XOR2_X1 U902 ( .A(round_inst_srout2_w[57]), .B(n590), .Z(final_w_k[9]) );
  MUX2_X1 U903 ( .A(k[72]), .B(k[73]), .S(enc), .Z(n591) );
  XOR2_X1 U904 ( .A(round_inst_srout2_w[56]), .B(n591), .Z(final_w_k[8]) );
  MUX2_X1 U905 ( .A(k[71]), .B(k[72]), .S(enc), .Z(n592) );
  XOR2_X1 U906 ( .A(round_inst_srout2_w[39]), .B(n592), .Z(final_w_k[7]) );
  MUX2_X1 U907 ( .A(k[70]), .B(k[71]), .S(enc), .Z(n593) );
  XOR2_X1 U908 ( .A(round_inst_srout2_w[38]), .B(n593), .Z(final_w_k[6]) );
  MUX2_X1 U909 ( .A(k[127]), .B(k[64]), .S(enc), .Z(n594) );
  XOR2_X1 U910 ( .A(round_inst_srout2_w[63]), .B(n594), .Z(final_w_k[63]) );
  MUX2_X1 U911 ( .A(k[126]), .B(k[127]), .S(enc), .Z(n595) );
  XOR2_X1 U912 ( .A(round_inst_srout2_w[62]), .B(n595), .Z(final_w_k[62]) );
  MUX2_X1 U913 ( .A(k[125]), .B(k[126]), .S(enc), .Z(n596) );
  XOR2_X1 U914 ( .A(round_inst_srout2_w[61]), .B(n596), .Z(final_w_k[61]) );
  MUX2_X1 U915 ( .A(k[124]), .B(k[125]), .S(enc), .Z(n597) );
  XOR2_X1 U916 ( .A(round_inst_srout2_w[60]), .B(n597), .Z(final_w_k[60]) );
  MUX2_X1 U917 ( .A(k[69]), .B(k[70]), .S(enc), .Z(n598) );
  XOR2_X1 U918 ( .A(round_inst_srout2_w[37]), .B(n598), .Z(final_w_k[5]) );
  MUX2_X1 U919 ( .A(k[123]), .B(k[124]), .S(enc), .Z(n599) );
  XOR2_X1 U920 ( .A(round_inst_srout2_w[43]), .B(n599), .Z(final_w_k[59]) );
  MUX2_X1 U921 ( .A(k[122]), .B(k[123]), .S(enc), .Z(n600) );
  XOR2_X1 U922 ( .A(round_inst_srout2_w[42]), .B(n600), .Z(final_w_k[58]) );
  MUX2_X1 U923 ( .A(k[121]), .B(k[122]), .S(enc), .Z(n601) );
  XOR2_X1 U924 ( .A(round_inst_srout2_w[41]), .B(n601), .Z(final_w_k[57]) );
  MUX2_X1 U925 ( .A(k[120]), .B(k[121]), .S(enc), .Z(n602) );
  XOR2_X1 U926 ( .A(round_inst_srout2_w[40]), .B(n602), .Z(final_w_k[56]) );
  MUX2_X1 U927 ( .A(k[119]), .B(k[120]), .S(enc), .Z(n603) );
  XOR2_X1 U928 ( .A(round_inst_srout2_w[23]), .B(n603), .Z(final_w_k[55]) );
  MUX2_X1 U929 ( .A(k[118]), .B(k[119]), .S(enc), .Z(n604) );
  XOR2_X1 U930 ( .A(round_inst_srout2_w[22]), .B(n604), .Z(final_w_k[54]) );
  MUX2_X1 U931 ( .A(k[117]), .B(k[118]), .S(enc), .Z(n605) );
  XOR2_X1 U932 ( .A(round_inst_srout2_w[21]), .B(n605), .Z(final_w_k[53]) );
  MUX2_X1 U933 ( .A(k[116]), .B(k[117]), .S(enc), .Z(n606) );
  XOR2_X1 U934 ( .A(round_inst_srout2_w[20]), .B(n606), .Z(final_w_k[52]) );
  MUX2_X1 U935 ( .A(k[115]), .B(k[116]), .S(enc), .Z(n607) );
  XOR2_X1 U936 ( .A(round_inst_srout2_w[3]), .B(n607), .Z(final_w_k[51]) );
  MUX2_X1 U937 ( .A(k[114]), .B(k[115]), .S(enc), .Z(n608) );
  XOR2_X1 U938 ( .A(round_inst_srout2_w[2]), .B(n608), .Z(final_w_k[50]) );
  MUX2_X1 U939 ( .A(k[68]), .B(k[69]), .S(enc), .Z(n609) );
  XOR2_X1 U940 ( .A(round_inst_srout2_w[36]), .B(n609), .Z(final_w_k[4]) );
  MUX2_X1 U941 ( .A(k[113]), .B(k[114]), .S(enc), .Z(n610) );
  XOR2_X1 U942 ( .A(round_inst_srout2_w[1]), .B(n610), .Z(final_w_k[49]) );
  MUX2_X1 U943 ( .A(k[112]), .B(k[113]), .S(enc), .Z(n611) );
  XOR2_X1 U944 ( .A(round_inst_srout2_w[0]), .B(n611), .Z(final_w_k[48]) );
  MUX2_X1 U945 ( .A(k[111]), .B(k[112]), .S(enc), .Z(n612) );
  XOR2_X1 U946 ( .A(round_inst_srout2_w[47]), .B(n612), .Z(final_w_k[47]) );
  MUX2_X1 U947 ( .A(k[110]), .B(k[111]), .S(enc), .Z(n613) );
  XOR2_X1 U948 ( .A(round_inst_srout2_w[46]), .B(n613), .Z(final_w_k[46]) );
  MUX2_X1 U949 ( .A(k[109]), .B(k[110]), .S(enc), .Z(n614) );
  XOR2_X1 U950 ( .A(round_inst_srout2_w[45]), .B(n614), .Z(final_w_k[45]) );
  MUX2_X1 U951 ( .A(k[108]), .B(k[109]), .S(enc), .Z(n615) );
  XOR2_X1 U952 ( .A(round_inst_srout2_w[44]), .B(n615), .Z(final_w_k[44]) );
  MUX2_X1 U953 ( .A(k[107]), .B(k[108]), .S(enc), .Z(n616) );
  XOR2_X1 U954 ( .A(round_inst_srout2_w[27]), .B(n616), .Z(final_w_k[43]) );
  MUX2_X1 U955 ( .A(k[106]), .B(k[107]), .S(enc), .Z(n617) );
  XOR2_X1 U956 ( .A(round_inst_srout2_w[26]), .B(n617), .Z(final_w_k[42]) );
  MUX2_X1 U957 ( .A(k[105]), .B(k[106]), .S(enc), .Z(n618) );
  XOR2_X1 U958 ( .A(round_inst_srout2_w[25]), .B(n618), .Z(final_w_k[41]) );
  MUX2_X1 U959 ( .A(k[104]), .B(k[105]), .S(enc), .Z(n619) );
  XOR2_X1 U960 ( .A(round_inst_srout2_w[24]), .B(n619), .Z(final_w_k[40]) );
  MUX2_X1 U961 ( .A(k[67]), .B(k[68]), .S(enc), .Z(n620) );
  XOR2_X1 U962 ( .A(round_inst_srout2_w[19]), .B(n620), .Z(final_w_k[3]) );
  MUX2_X1 U963 ( .A(k[103]), .B(k[104]), .S(enc), .Z(n621) );
  XOR2_X1 U964 ( .A(round_inst_srout2_w[7]), .B(n621), .Z(final_w_k[39]) );
  MUX2_X1 U965 ( .A(k[102]), .B(k[103]), .S(enc), .Z(n622) );
  XOR2_X1 U966 ( .A(round_inst_srout2_w[6]), .B(n622), .Z(final_w_k[38]) );
  MUX2_X1 U967 ( .A(k[101]), .B(k[102]), .S(enc), .Z(n623) );
  XOR2_X1 U968 ( .A(round_inst_srout2_w[5]), .B(n623), .Z(final_w_k[37]) );
  MUX2_X1 U969 ( .A(k[100]), .B(k[101]), .S(enc), .Z(n624) );
  XOR2_X1 U970 ( .A(round_inst_srout2_w[4]), .B(n624), .Z(final_w_k[36]) );
  MUX2_X1 U971 ( .A(k[99]), .B(k[100]), .S(enc), .Z(n625) );
  XOR2_X1 U972 ( .A(round_inst_srout2_w[51]), .B(n625), .Z(final_w_k[35]) );
  MUX2_X1 U973 ( .A(k[98]), .B(k[99]), .S(enc), .Z(n626) );
  XOR2_X1 U974 ( .A(round_inst_srout2_w[50]), .B(n626), .Z(final_w_k[34]) );
  MUX2_X1 U975 ( .A(k[97]), .B(k[98]), .S(enc), .Z(n627) );
  XOR2_X1 U976 ( .A(round_inst_srout2_w[49]), .B(n627), .Z(final_w_k[33]) );
  MUX2_X1 U977 ( .A(k[96]), .B(k[97]), .S(enc), .Z(n628) );
  XOR2_X1 U978 ( .A(round_inst_srout2_w[48]), .B(n628), .Z(final_w_k[32]) );
  MUX2_X1 U979 ( .A(k[95]), .B(k[96]), .S(enc), .Z(n629) );
  XOR2_X1 U980 ( .A(round_inst_srout2_w[31]), .B(n629), .Z(final_w_k[31]) );
  MUX2_X1 U981 ( .A(k[94]), .B(k[95]), .S(enc), .Z(n630) );
  XOR2_X1 U982 ( .A(round_inst_srout2_w[30]), .B(n630), .Z(final_w_k[30]) );
  MUX2_X1 U983 ( .A(k[66]), .B(k[67]), .S(enc), .Z(n631) );
  XOR2_X1 U984 ( .A(round_inst_srout2_w[18]), .B(n631), .Z(final_w_k[2]) );
  MUX2_X1 U985 ( .A(k[93]), .B(k[94]), .S(enc), .Z(n632) );
  XOR2_X1 U986 ( .A(round_inst_srout2_w[29]), .B(n632), .Z(final_w_k[29]) );
  MUX2_X1 U987 ( .A(k[92]), .B(k[93]), .S(enc), .Z(n633) );
  XOR2_X1 U988 ( .A(round_inst_srout2_w[28]), .B(n633), .Z(final_w_k[28]) );
  MUX2_X1 U989 ( .A(k[91]), .B(k[92]), .S(enc), .Z(n634) );
  XOR2_X1 U990 ( .A(round_inst_srout2_w[11]), .B(n634), .Z(final_w_k[27]) );
  MUX2_X1 U991 ( .A(k[90]), .B(k[91]), .S(enc), .Z(n635) );
  XOR2_X1 U992 ( .A(round_inst_srout2_w[10]), .B(n635), .Z(final_w_k[26]) );
  MUX2_X1 U993 ( .A(k[89]), .B(k[90]), .S(enc), .Z(n636) );
  XOR2_X1 U994 ( .A(round_inst_srout2_w[9]), .B(n636), .Z(final_w_k[25]) );
  MUX2_X1 U995 ( .A(k[88]), .B(k[89]), .S(enc), .Z(n637) );
  XOR2_X1 U996 ( .A(round_inst_srout2_w[8]), .B(n637), .Z(final_w_k[24]) );
  MUX2_X1 U997 ( .A(k[87]), .B(k[88]), .S(enc), .Z(n638) );
  XOR2_X1 U998 ( .A(round_inst_srout2_w[55]), .B(n638), .Z(final_w_k[23]) );
  MUX2_X1 U999 ( .A(k[86]), .B(k[87]), .S(enc), .Z(n639) );
  XOR2_X1 U1000 ( .A(round_inst_srout2_w[54]), .B(n639), .Z(final_w_k[22]) );
  MUX2_X1 U1001 ( .A(k[85]), .B(k[86]), .S(enc), .Z(n640) );
  XOR2_X1 U1002 ( .A(round_inst_srout2_w[53]), .B(n640), .Z(final_w_k[21]) );
  MUX2_X1 U1003 ( .A(k[84]), .B(k[85]), .S(enc), .Z(n641) );
  XOR2_X1 U1004 ( .A(round_inst_srout2_w[52]), .B(n641), .Z(final_w_k[20]) );
  MUX2_X1 U1005 ( .A(k[65]), .B(k[66]), .S(enc), .Z(n642) );
  XOR2_X1 U1006 ( .A(round_inst_srout2_w[17]), .B(n642), .Z(final_w_k[1]) );
  MUX2_X1 U1007 ( .A(k[83]), .B(k[84]), .S(enc), .Z(n643) );
  XOR2_X1 U1008 ( .A(round_inst_srout2_w[35]), .B(n643), .Z(final_w_k[19]) );
  MUX2_X1 U1009 ( .A(k[82]), .B(k[83]), .S(enc), .Z(n644) );
  XOR2_X1 U1010 ( .A(round_inst_srout2_w[34]), .B(n644), .Z(final_w_k[18]) );
  MUX2_X1 U1011 ( .A(k[81]), .B(k[82]), .S(enc), .Z(n645) );
  XOR2_X1 U1012 ( .A(round_inst_srout2_w[33]), .B(n645), .Z(final_w_k[17]) );
  MUX2_X1 U1013 ( .A(k[80]), .B(k[81]), .S(enc), .Z(n646) );
  XOR2_X1 U1014 ( .A(round_inst_srout2_w[32]), .B(n646), .Z(final_w_k[16]) );
  MUX2_X1 U1015 ( .A(k[79]), .B(k[80]), .S(enc), .Z(n647) );
  XOR2_X1 U1016 ( .A(round_inst_srout2_w[15]), .B(n647), .Z(final_w_k[15]) );
  MUX2_X1 U1017 ( .A(k[78]), .B(k[79]), .S(enc), .Z(n648) );
  XOR2_X1 U1018 ( .A(round_inst_srout2_w[14]), .B(n648), .Z(final_w_k[14]) );
  MUX2_X1 U1019 ( .A(k[77]), .B(k[78]), .S(enc), .Z(n649) );
  XOR2_X1 U1020 ( .A(round_inst_srout2_w[13]), .B(n649), .Z(final_w_k[13]) );
  MUX2_X1 U1021 ( .A(k[76]), .B(k[77]), .S(enc), .Z(n650) );
  XOR2_X1 U1022 ( .A(round_inst_srout2_w[12]), .B(n650), .Z(final_w_k[12]) );
  MUX2_X1 U1023 ( .A(k[75]), .B(k[76]), .S(enc), .Z(n651) );
  XOR2_X1 U1024 ( .A(round_inst_srout2_w[59]), .B(n651), .Z(final_w_k[11]) );
  MUX2_X1 U1025 ( .A(k[74]), .B(k[75]), .S(enc), .Z(n652) );
  XOR2_X1 U1026 ( .A(round_inst_srout2_w[58]), .B(n652), .Z(final_w_k[10]) );
  MUX2_X1 U1027 ( .A(k[64]), .B(kext_64_), .S(enc), .Z(n653) );
  XOR2_X1 U1028 ( .A(round_inst_srout2_w[16]), .B(n653), .Z(final_w_k[0]) );
  XOR2_X1 k_inst_U1 ( .A(k[65]), .B(k[127]), .Z(kext_64_) );
  MUX2_X1 mux_w_U68 ( .A(rout_w[35]), .B(init_w[35]), .S(mux_w_n138), .Z(
        state_w[35]) );
  MUX2_X1 mux_w_U67 ( .A(rout_w[34]), .B(init_w[34]), .S(mux_w_n137), .Z(
        state_w[34]) );
  MUX2_X1 mux_w_U66 ( .A(rout_w[33]), .B(init_w[33]), .S(mux_w_n136), .Z(
        state_w[33]) );
  MUX2_X1 mux_w_U65 ( .A(rout_w[32]), .B(init_w[32]), .S(mux_w_n136), .Z(
        state_w[32]) );
  MUX2_X1 mux_w_U64 ( .A(rout_w[31]), .B(init_w[31]), .S(mux_w_n136), .Z(
        state_w[31]) );
  MUX2_X1 mux_w_U63 ( .A(rout_w[30]), .B(init_w[30]), .S(mux_w_n138), .Z(
        state_w[30]) );
  MUX2_X1 mux_w_U62 ( .A(rout_w[29]), .B(init_w[29]), .S(mux_w_n137), .Z(
        state_w[29]) );
  MUX2_X1 mux_w_U61 ( .A(rout_w[28]), .B(init_w[28]), .S(mux_w_n136), .Z(
        state_w[28]) );
  MUX2_X1 mux_w_U60 ( .A(rout_w[27]), .B(init_w[27]), .S(mux_w_n138), .Z(
        state_w[27]) );
  MUX2_X1 mux_w_U59 ( .A(rout_w[26]), .B(init_w[26]), .S(mux_w_n137), .Z(
        state_w[26]) );
  MUX2_X1 mux_w_U58 ( .A(rout_w[25]), .B(init_w[25]), .S(mux_w_n136), .Z(
        state_w[25]) );
  MUX2_X1 mux_w_U57 ( .A(rout_w[24]), .B(init_w[24]), .S(mux_w_n138), .Z(
        state_w[24]) );
  MUX2_X1 mux_w_U56 ( .A(rout_w[23]), .B(init_w[23]), .S(mux_w_n137), .Z(
        state_w[23]) );
  MUX2_X1 mux_w_U55 ( .A(rout_w[22]), .B(init_w[22]), .S(mux_w_n136), .Z(
        state_w[22]) );
  MUX2_X1 mux_w_U54 ( .A(rout_w[21]), .B(init_w[21]), .S(mux_w_n138), .Z(
        state_w[21]) );
  MUX2_X1 mux_w_U53 ( .A(rout_w[20]), .B(init_w[20]), .S(mux_w_n137), .Z(
        state_w[20]) );
  MUX2_X1 mux_w_U52 ( .A(rout_w[19]), .B(init_w[19]), .S(start_sig), .Z(
        state_w[19]) );
  MUX2_X1 mux_w_U51 ( .A(rout_w[18]), .B(init_w[18]), .S(mux_w_n138), .Z(
        state_w[18]) );
  MUX2_X1 mux_w_U50 ( .A(rout_w[17]), .B(init_w[17]), .S(mux_w_n137), .Z(
        state_w[17]) );
  MUX2_X1 mux_w_U49 ( .A(rout_w[16]), .B(init_w[16]), .S(mux_w_n136), .Z(
        state_w[16]) );
  MUX2_X1 mux_w_U48 ( .A(rout_w[15]), .B(init_w[15]), .S(start_sig), .Z(
        state_w[15]) );
  MUX2_X1 mux_w_U47 ( .A(rout_w[14]), .B(init_w[14]), .S(start_sig), .Z(
        state_w[14]) );
  MUX2_X1 mux_w_U46 ( .A(rout_w[13]), .B(init_w[13]), .S(mux_w_n138), .Z(
        state_w[13]) );
  MUX2_X1 mux_w_U45 ( .A(rout_w[12]), .B(init_w[12]), .S(mux_w_n137), .Z(
        state_w[12]) );
  MUX2_X1 mux_w_U44 ( .A(rout_w[11]), .B(init_w[11]), .S(mux_w_n138), .Z(
        state_w[11]) );
  MUX2_X1 mux_w_U43 ( .A(rout_w[10]), .B(init_w[10]), .S(mux_w_n137), .Z(
        state_w[10]) );
  MUX2_X1 mux_w_U42 ( .A(rout_w[9]), .B(init_w[9]), .S(mux_w_n136), .Z(
        state_w[9]) );
  MUX2_X1 mux_w_U41 ( .A(rout_w[8]), .B(init_w[8]), .S(start_sig), .Z(
        state_w[8]) );
  MUX2_X1 mux_w_U40 ( .A(rout_w[7]), .B(init_w[7]), .S(mux_w_n136), .Z(
        state_w[7]) );
  MUX2_X1 mux_w_U39 ( .A(rout_w[4]), .B(init_w[4]), .S(mux_w_n136), .Z(
        state_w[4]) );
  MUX2_X1 mux_w_U38 ( .A(rout_w[3]), .B(init_w[3]), .S(mux_w_n136), .Z(
        state_w[3]) );
  MUX2_X1 mux_w_U37 ( .A(rout_w[2]), .B(init_w[2]), .S(mux_w_n136), .Z(
        state_w[2]) );
  MUX2_X1 mux_w_U36 ( .A(rout_w[1]), .B(init_w[1]), .S(mux_w_n136), .Z(
        state_w[1]) );
  MUX2_X1 mux_w_U35 ( .A(rout_w[0]), .B(init_w[0]), .S(mux_w_n136), .Z(
        state_w[0]) );
  MUX2_X1 mux_w_U34 ( .A(rout_w[59]), .B(init_w[59]), .S(mux_w_n136), .Z(
        state_w[59]) );
  MUX2_X1 mux_w_U33 ( .A(rout_w[58]), .B(init_w[58]), .S(mux_w_n136), .Z(
        state_w[58]) );
  MUX2_X1 mux_w_U32 ( .A(rout_w[57]), .B(init_w[57]), .S(mux_w_n136), .Z(
        state_w[57]) );
  MUX2_X1 mux_w_U31 ( .A(rout_w[56]), .B(init_w[56]), .S(mux_w_n136), .Z(
        state_w[56]) );
  MUX2_X1 mux_w_U30 ( .A(rout_w[55]), .B(init_w[55]), .S(mux_w_n136), .Z(
        state_w[55]) );
  MUX2_X1 mux_w_U29 ( .A(rout_w[54]), .B(init_w[54]), .S(mux_w_n136), .Z(
        state_w[54]) );
  INV_X1 mux_w_U28 ( .A(mux_w_n135), .ZN(mux_w_n136) );
  MUX2_X1 mux_w_U27 ( .A(rout_w[53]), .B(init_w[53]), .S(mux_w_n137), .Z(
        state_w[53]) );
  MUX2_X1 mux_w_U26 ( .A(rout_w[52]), .B(init_w[52]), .S(mux_w_n137), .Z(
        state_w[52]) );
  MUX2_X1 mux_w_U25 ( .A(rout_w[51]), .B(init_w[51]), .S(mux_w_n137), .Z(
        state_w[51]) );
  MUX2_X1 mux_w_U24 ( .A(rout_w[50]), .B(init_w[50]), .S(mux_w_n137), .Z(
        state_w[50]) );
  MUX2_X1 mux_w_U23 ( .A(rout_w[49]), .B(init_w[49]), .S(mux_w_n137), .Z(
        state_w[49]) );
  MUX2_X1 mux_w_U22 ( .A(rout_w[48]), .B(init_w[48]), .S(mux_w_n137), .Z(
        state_w[48]) );
  MUX2_X1 mux_w_U21 ( .A(rout_w[47]), .B(init_w[47]), .S(mux_w_n137), .Z(
        state_w[47]) );
  MUX2_X1 mux_w_U20 ( .A(rout_w[46]), .B(init_w[46]), .S(mux_w_n137), .Z(
        state_w[46]) );
  MUX2_X1 mux_w_U19 ( .A(rout_w[45]), .B(init_w[45]), .S(mux_w_n137), .Z(
        state_w[45]) );
  MUX2_X1 mux_w_U18 ( .A(rout_w[44]), .B(init_w[44]), .S(mux_w_n137), .Z(
        state_w[44]) );
  MUX2_X1 mux_w_U17 ( .A(rout_w[43]), .B(init_w[43]), .S(mux_w_n137), .Z(
        state_w[43]) );
  MUX2_X1 mux_w_U16 ( .A(rout_w[42]), .B(init_w[42]), .S(mux_w_n137), .Z(
        state_w[42]) );
  INV_X1 mux_w_U15 ( .A(mux_w_n135), .ZN(mux_w_n137) );
  MUX2_X1 mux_w_U14 ( .A(rout_w[41]), .B(init_w[41]), .S(mux_w_n138), .Z(
        state_w[41]) );
  MUX2_X1 mux_w_U13 ( .A(rout_w[40]), .B(init_w[40]), .S(mux_w_n138), .Z(
        state_w[40]) );
  MUX2_X1 mux_w_U12 ( .A(rout_w[39]), .B(init_w[39]), .S(mux_w_n138), .Z(
        state_w[39]) );
  MUX2_X1 mux_w_U11 ( .A(rout_w[38]), .B(init_w[38]), .S(mux_w_n138), .Z(
        state_w[38]) );
  MUX2_X1 mux_w_U10 ( .A(rout_w[37]), .B(init_w[37]), .S(mux_w_n138), .Z(
        state_w[37]) );
  MUX2_X1 mux_w_U9 ( .A(rout_w[36]), .B(init_w[36]), .S(mux_w_n138), .Z(
        state_w[36]) );
  MUX2_X1 mux_w_U8 ( .A(rout_w[63]), .B(init_w[63]), .S(mux_w_n138), .Z(
        state_w[63]) );
  MUX2_X1 mux_w_U7 ( .A(rout_w[62]), .B(init_w[62]), .S(mux_w_n138), .Z(
        state_w[62]) );
  MUX2_X1 mux_w_U6 ( .A(rout_w[61]), .B(init_w[61]), .S(mux_w_n138), .Z(
        state_w[61]) );
  MUX2_X1 mux_w_U5 ( .A(rout_w[60]), .B(init_w[60]), .S(mux_w_n138), .Z(
        state_w[60]) );
  MUX2_X1 mux_w_U4 ( .A(rout_w[6]), .B(init_w[6]), .S(mux_w_n138), .Z(
        state_w[6]) );
  MUX2_X1 mux_w_U3 ( .A(rout_w[5]), .B(init_w[5]), .S(mux_w_n138), .Z(
        state_w[5]) );
  INV_X1 mux_w_U2 ( .A(mux_w_n135), .ZN(mux_w_n138) );
  INV_X1 mux_w_U1 ( .A(start_sig), .ZN(mux_w_n135) );
  MUX2_X1 mux_x_U68 ( .A(rout_x[34]), .B(p1[18]), .S(mux_x_n266), .Z(
        state_x[34]) );
  MUX2_X1 mux_x_U67 ( .A(rout_x[33]), .B(p1[17]), .S(mux_x_n265), .Z(
        state_x[33]) );
  MUX2_X1 mux_x_U66 ( .A(rout_x[32]), .B(p1[16]), .S(mux_x_n265), .Z(
        state_x[32]) );
  MUX2_X1 mux_x_U65 ( .A(rout_x[30]), .B(p1[30]), .S(mux_x_n264), .Z(
        state_x[30]) );
  MUX2_X1 mux_x_U64 ( .A(rout_x[29]), .B(p1[29]), .S(mux_x_n264), .Z(
        state_x[29]) );
  MUX2_X1 mux_x_U63 ( .A(rout_x[28]), .B(p1[28]), .S(mux_x_n264), .Z(
        state_x[28]) );
  MUX2_X1 mux_x_U62 ( .A(rout_x[27]), .B(p1[43]), .S(mux_x_n264), .Z(
        state_x[27]) );
  MUX2_X1 mux_x_U61 ( .A(rout_x[26]), .B(p1[42]), .S(mux_x_n264), .Z(
        state_x[26]) );
  MUX2_X1 mux_x_U60 ( .A(rout_x[25]), .B(p1[41]), .S(mux_x_n264), .Z(
        state_x[25]) );
  MUX2_X1 mux_x_U59 ( .A(rout_x[24]), .B(p1[40]), .S(mux_x_n264), .Z(
        state_x[24]) );
  MUX2_X1 mux_x_U58 ( .A(rout_x[23]), .B(p1[55]), .S(mux_x_n264), .Z(
        state_x[23]) );
  MUX2_X1 mux_x_U57 ( .A(rout_x[22]), .B(p1[54]), .S(mux_x_n264), .Z(
        state_x[22]) );
  MUX2_X1 mux_x_U56 ( .A(rout_x[21]), .B(p1[53]), .S(mux_x_n264), .Z(
        state_x[21]) );
  MUX2_X1 mux_x_U55 ( .A(rout_x[20]), .B(p1[52]), .S(mux_x_n264), .Z(
        state_x[20]) );
  MUX2_X1 mux_x_U54 ( .A(rout_x[18]), .B(p1[2]), .S(mux_x_n264), .Z(
        state_x[18]) );
  MUX2_X1 mux_x_U53 ( .A(rout_x[17]), .B(p1[1]), .S(mux_x_n264), .Z(
        state_x[17]) );
  MUX2_X1 mux_x_U52 ( .A(rout_x[16]), .B(p1[0]), .S(mux_x_n264), .Z(
        state_x[16]) );
  MUX2_X1 mux_x_U51 ( .A(rout_x[14]), .B(p1[14]), .S(mux_x_n264), .Z(
        state_x[14]) );
  MUX2_X1 mux_x_U50 ( .A(rout_x[13]), .B(p1[13]), .S(mux_x_n264), .Z(
        state_x[13]) );
  MUX2_X1 mux_x_U49 ( .A(rout_x[12]), .B(p1[12]), .S(mux_x_n264), .Z(
        state_x[12]) );
  MUX2_X1 mux_x_U48 ( .A(rout_x[11]), .B(p1[27]), .S(mux_x_n265), .Z(
        state_x[11]) );
  MUX2_X1 mux_x_U47 ( .A(rout_x[10]), .B(p1[26]), .S(mux_x_n266), .Z(
        state_x[10]) );
  MUX2_X1 mux_x_U46 ( .A(rout_x[9]), .B(p1[25]), .S(mux_x_n264), .Z(state_x[9]) );
  MUX2_X1 mux_x_U45 ( .A(rout_x[7]), .B(p1[39]), .S(mux_x_n264), .Z(state_x[7]) );
  MUX2_X1 mux_x_U44 ( .A(rout_x[6]), .B(p1[38]), .S(mux_x_n264), .Z(state_x[6]) );
  MUX2_X1 mux_x_U43 ( .A(rout_x[3]), .B(p1[51]), .S(mux_x_n264), .Z(state_x[3]) );
  MUX2_X1 mux_x_U42 ( .A(rout_x[2]), .B(p1[50]), .S(mux_x_n264), .Z(state_x[2]) );
  MUX2_X1 mux_x_U41 ( .A(rout_x[1]), .B(p1[49]), .S(mux_x_n266), .Z(state_x[1]) );
  MUX2_X1 mux_x_U40 ( .A(rout_x[0]), .B(p1[48]), .S(mux_x_n265), .Z(state_x[0]) );
  MUX2_X1 mux_x_U39 ( .A(rout_x[59]), .B(p1[11]), .S(mux_x_n264), .Z(
        state_x[59]) );
  MUX2_X1 mux_x_U38 ( .A(rout_x[58]), .B(p1[10]), .S(mux_x_n264), .Z(
        state_x[58]) );
  MUX2_X1 mux_x_U37 ( .A(rout_x[57]), .B(p1[9]), .S(mux_x_n266), .Z(
        state_x[57]) );
  MUX2_X1 mux_x_U36 ( .A(rout_x[56]), .B(p1[8]), .S(mux_x_n265), .Z(
        state_x[56]) );
  MUX2_X1 mux_x_U35 ( .A(rout_x[55]), .B(p1[23]), .S(mux_x_n264), .Z(
        state_x[55]) );
  MUX2_X1 mux_x_U34 ( .A(rout_x[54]), .B(p1[22]), .S(mux_x_n264), .Z(
        state_x[54]) );
  MUX2_X1 mux_x_U33 ( .A(rout_x[53]), .B(p1[21]), .S(mux_x_n266), .Z(
        state_x[53]) );
  MUX2_X1 mux_x_U32 ( .A(rout_x[52]), .B(p1[20]), .S(mux_x_n265), .Z(
        state_x[52]) );
  MUX2_X1 mux_x_U31 ( .A(rout_x[51]), .B(p1[35]), .S(mux_x_n264), .Z(
        state_x[51]) );
  MUX2_X1 mux_x_U30 ( .A(rout_x[50]), .B(p1[34]), .S(mux_x_n264), .Z(
        state_x[50]) );
  MUX2_X1 mux_x_U29 ( .A(rout_x[49]), .B(p1[33]), .S(mux_x_n266), .Z(
        state_x[49]) );
  MUX2_X1 mux_x_U28 ( .A(rout_x[48]), .B(p1[32]), .S(mux_x_n265), .Z(
        state_x[48]) );
  MUX2_X1 mux_x_U27 ( .A(rout_x[47]), .B(p1[47]), .S(mux_x_n265), .Z(
        state_x[47]) );
  MUX2_X1 mux_x_U26 ( .A(rout_x[46]), .B(p1[46]), .S(mux_x_n265), .Z(
        state_x[46]) );
  MUX2_X1 mux_x_U25 ( .A(rout_x[45]), .B(p1[45]), .S(mux_x_n265), .Z(
        state_x[45]) );
  MUX2_X1 mux_x_U24 ( .A(rout_x[44]), .B(p1[44]), .S(mux_x_n265), .Z(
        state_x[44]) );
  MUX2_X1 mux_x_U23 ( .A(rout_x[43]), .B(p1[59]), .S(mux_x_n265), .Z(
        state_x[43]) );
  MUX2_X1 mux_x_U22 ( .A(rout_x[42]), .B(p1[58]), .S(mux_x_n265), .Z(
        state_x[42]) );
  MUX2_X1 mux_x_U21 ( .A(rout_x[41]), .B(p1[57]), .S(mux_x_n265), .Z(
        state_x[41]) );
  MUX2_X1 mux_x_U20 ( .A(rout_x[40]), .B(p1[56]), .S(mux_x_n265), .Z(
        state_x[40]) );
  MUX2_X1 mux_x_U19 ( .A(rout_x[39]), .B(p1[7]), .S(mux_x_n265), .Z(
        state_x[39]) );
  MUX2_X1 mux_x_U18 ( .A(rout_x[38]), .B(p1[6]), .S(mux_x_n265), .Z(
        state_x[38]) );
  MUX2_X1 mux_x_U17 ( .A(rout_x[37]), .B(p1[5]), .S(mux_x_n265), .Z(
        state_x[37]) );
  INV_X1 mux_x_U16 ( .A(mux_x_n263), .ZN(mux_x_n265) );
  MUX2_X1 mux_x_U15 ( .A(rout_x[36]), .B(p1[4]), .S(mux_x_n266), .Z(
        state_x[36]) );
  MUX2_X1 mux_x_U14 ( .A(rout_x[63]), .B(p1[63]), .S(mux_x_n266), .Z(
        state_x[63]) );
  MUX2_X1 mux_x_U13 ( .A(rout_x[62]), .B(p1[62]), .S(mux_x_n266), .Z(
        state_x[62]) );
  MUX2_X1 mux_x_U12 ( .A(rout_x[61]), .B(p1[61]), .S(mux_x_n266), .Z(
        state_x[61]) );
  MUX2_X1 mux_x_U11 ( .A(rout_x[60]), .B(p1[60]), .S(mux_x_n266), .Z(
        state_x[60]) );
  MUX2_X1 mux_x_U10 ( .A(rout_x[35]), .B(p1[19]), .S(mux_x_n266), .Z(
        state_x[35]) );
  MUX2_X1 mux_x_U9 ( .A(rout_x[31]), .B(p1[31]), .S(mux_x_n266), .Z(
        state_x[31]) );
  MUX2_X1 mux_x_U8 ( .A(rout_x[19]), .B(p1[3]), .S(mux_x_n266), .Z(state_x[19]) );
  MUX2_X1 mux_x_U7 ( .A(rout_x[15]), .B(p1[15]), .S(mux_x_n266), .Z(
        state_x[15]) );
  MUX2_X1 mux_x_U6 ( .A(rout_x[8]), .B(p1[24]), .S(mux_x_n266), .Z(state_x[8])
         );
  MUX2_X1 mux_x_U5 ( .A(rout_x[5]), .B(p1[37]), .S(mux_x_n266), .Z(state_x[5])
         );
  MUX2_X1 mux_x_U4 ( .A(rout_x[4]), .B(p1[36]), .S(mux_x_n266), .Z(state_x[4])
         );
  INV_X1 mux_x_U3 ( .A(mux_x_n263), .ZN(mux_x_n266) );
  INV_X1 mux_x_U2 ( .A(start_sig), .ZN(mux_x_n263) );
  INV_X2 mux_x_U1 ( .A(mux_x_n263), .ZN(mux_x_n264) );
  MUX2_X1 mux_y_U68 ( .A(rout_y[35]), .B(p2[19]), .S(mux_y_n266), .Z(
        state_y[35]) );
  MUX2_X1 mux_y_U67 ( .A(rout_y[34]), .B(p2[18]), .S(mux_y_n265), .Z(
        state_y[34]) );
  MUX2_X1 mux_y_U66 ( .A(rout_y[33]), .B(p2[17]), .S(mux_y_n265), .Z(
        state_y[33]) );
  MUX2_X1 mux_y_U65 ( .A(rout_y[32]), .B(p2[16]), .S(mux_y_n264), .Z(
        state_y[32]) );
  MUX2_X1 mux_y_U64 ( .A(rout_y[31]), .B(p2[31]), .S(mux_y_n264), .Z(
        state_y[31]) );
  MUX2_X1 mux_y_U63 ( .A(rout_y[30]), .B(p2[30]), .S(mux_y_n264), .Z(
        state_y[30]) );
  MUX2_X1 mux_y_U62 ( .A(rout_y[28]), .B(p2[28]), .S(mux_y_n264), .Z(
        state_y[28]) );
  MUX2_X1 mux_y_U61 ( .A(rout_y[27]), .B(p2[43]), .S(mux_y_n264), .Z(
        state_y[27]) );
  MUX2_X1 mux_y_U60 ( .A(rout_y[26]), .B(p2[42]), .S(mux_y_n264), .Z(
        state_y[26]) );
  MUX2_X1 mux_y_U59 ( .A(rout_y[24]), .B(p2[40]), .S(mux_y_n264), .Z(
        state_y[24]) );
  MUX2_X1 mux_y_U58 ( .A(rout_y[23]), .B(p2[55]), .S(mux_y_n264), .Z(
        state_y[23]) );
  MUX2_X1 mux_y_U57 ( .A(rout_y[22]), .B(p2[54]), .S(mux_y_n264), .Z(
        state_y[22]) );
  MUX2_X1 mux_y_U56 ( .A(rout_y[21]), .B(p2[53]), .S(mux_y_n264), .Z(
        state_y[21]) );
  MUX2_X1 mux_y_U55 ( .A(rout_y[20]), .B(p2[52]), .S(mux_y_n264), .Z(
        state_y[20]) );
  MUX2_X1 mux_y_U54 ( .A(rout_y[19]), .B(p2[3]), .S(mux_y_n264), .Z(
        state_y[19]) );
  MUX2_X1 mux_y_U53 ( .A(rout_y[18]), .B(p2[2]), .S(mux_y_n264), .Z(
        state_y[18]) );
  MUX2_X1 mux_y_U52 ( .A(rout_y[17]), .B(p2[1]), .S(mux_y_n264), .Z(
        state_y[17]) );
  MUX2_X1 mux_y_U51 ( .A(rout_y[16]), .B(p2[0]), .S(mux_y_n264), .Z(
        state_y[16]) );
  MUX2_X1 mux_y_U50 ( .A(rout_y[14]), .B(p2[14]), .S(mux_y_n264), .Z(
        state_y[14]) );
  MUX2_X1 mux_y_U49 ( .A(rout_y[13]), .B(p2[13]), .S(mux_y_n264), .Z(
        state_y[13]) );
  MUX2_X1 mux_y_U48 ( .A(rout_y[12]), .B(p2[12]), .S(mux_y_n264), .Z(
        state_y[12]) );
  MUX2_X1 mux_y_U47 ( .A(rout_y[10]), .B(p2[26]), .S(mux_y_n264), .Z(
        state_y[10]) );
  MUX2_X1 mux_y_U46 ( .A(rout_y[9]), .B(p2[25]), .S(mux_y_n264), .Z(state_y[9]) );
  MUX2_X1 mux_y_U45 ( .A(rout_y[8]), .B(p2[24]), .S(mux_y_n264), .Z(state_y[8]) );
  MUX2_X1 mux_y_U44 ( .A(rout_y[5]), .B(p2[37]), .S(mux_y_n266), .Z(state_y[5]) );
  MUX2_X1 mux_y_U43 ( .A(rout_y[4]), .B(p2[36]), .S(mux_y_n265), .Z(state_y[4]) );
  MUX2_X1 mux_y_U42 ( .A(rout_y[3]), .B(p2[51]), .S(mux_y_n266), .Z(state_y[3]) );
  MUX2_X1 mux_y_U41 ( .A(rout_y[2]), .B(p2[50]), .S(mux_y_n264), .Z(state_y[2]) );
  MUX2_X1 mux_y_U40 ( .A(rout_y[1]), .B(p2[49]), .S(mux_y_n265), .Z(state_y[1]) );
  MUX2_X1 mux_y_U39 ( .A(rout_y[0]), .B(p2[48]), .S(mux_y_n264), .Z(state_y[0]) );
  MUX2_X1 mux_y_U38 ( .A(rout_y[59]), .B(p2[11]), .S(mux_y_n264), .Z(
        state_y[59]) );
  MUX2_X1 mux_y_U37 ( .A(rout_y[58]), .B(p2[10]), .S(mux_y_n266), .Z(
        state_y[58]) );
  MUX2_X1 mux_y_U36 ( .A(rout_y[57]), .B(p2[9]), .S(mux_y_n265), .Z(
        state_y[57]) );
  MUX2_X1 mux_y_U35 ( .A(rout_y[56]), .B(p2[8]), .S(mux_y_n264), .Z(
        state_y[56]) );
  MUX2_X1 mux_y_U34 ( .A(rout_y[55]), .B(p2[23]), .S(mux_y_n264), .Z(
        state_y[55]) );
  MUX2_X1 mux_y_U33 ( .A(rout_y[54]), .B(p2[22]), .S(mux_y_n266), .Z(
        state_y[54]) );
  MUX2_X1 mux_y_U32 ( .A(rout_y[53]), .B(p2[21]), .S(mux_y_n265), .Z(
        state_y[53]) );
  MUX2_X1 mux_y_U31 ( .A(rout_y[52]), .B(p2[20]), .S(mux_y_n264), .Z(
        state_y[52]) );
  MUX2_X1 mux_y_U30 ( .A(rout_y[51]), .B(p2[35]), .S(mux_y_n264), .Z(
        state_y[51]) );
  MUX2_X1 mux_y_U29 ( .A(rout_y[50]), .B(p2[34]), .S(mux_y_n266), .Z(
        state_y[50]) );
  MUX2_X1 mux_y_U28 ( .A(rout_y[49]), .B(p2[33]), .S(mux_y_n265), .Z(
        state_y[49]) );
  MUX2_X1 mux_y_U27 ( .A(rout_y[48]), .B(p2[32]), .S(mux_y_n265), .Z(
        state_y[48]) );
  MUX2_X1 mux_y_U26 ( .A(rout_y[47]), .B(p2[47]), .S(mux_y_n265), .Z(
        state_y[47]) );
  MUX2_X1 mux_y_U25 ( .A(rout_y[46]), .B(p2[46]), .S(mux_y_n265), .Z(
        state_y[46]) );
  MUX2_X1 mux_y_U24 ( .A(rout_y[45]), .B(p2[45]), .S(mux_y_n265), .Z(
        state_y[45]) );
  MUX2_X1 mux_y_U23 ( .A(rout_y[44]), .B(p2[44]), .S(mux_y_n265), .Z(
        state_y[44]) );
  MUX2_X1 mux_y_U22 ( .A(rout_y[43]), .B(p2[59]), .S(mux_y_n265), .Z(
        state_y[43]) );
  MUX2_X1 mux_y_U21 ( .A(rout_y[42]), .B(p2[58]), .S(mux_y_n265), .Z(
        state_y[42]) );
  MUX2_X1 mux_y_U20 ( .A(rout_y[41]), .B(p2[57]), .S(mux_y_n265), .Z(
        state_y[41]) );
  MUX2_X1 mux_y_U19 ( .A(rout_y[40]), .B(p2[56]), .S(mux_y_n265), .Z(
        state_y[40]) );
  MUX2_X1 mux_y_U18 ( .A(rout_y[39]), .B(p2[7]), .S(mux_y_n265), .Z(
        state_y[39]) );
  MUX2_X1 mux_y_U17 ( .A(rout_y[38]), .B(p2[6]), .S(mux_y_n265), .Z(
        state_y[38]) );
  INV_X1 mux_y_U16 ( .A(mux_y_n263), .ZN(mux_y_n265) );
  MUX2_X1 mux_y_U15 ( .A(rout_y[37]), .B(p2[5]), .S(mux_y_n266), .Z(
        state_y[37]) );
  MUX2_X1 mux_y_U14 ( .A(rout_y[36]), .B(p2[4]), .S(mux_y_n266), .Z(
        state_y[36]) );
  MUX2_X1 mux_y_U13 ( .A(rout_y[63]), .B(p2[63]), .S(mux_y_n266), .Z(
        state_y[63]) );
  MUX2_X1 mux_y_U12 ( .A(rout_y[62]), .B(p2[62]), .S(mux_y_n266), .Z(
        state_y[62]) );
  MUX2_X1 mux_y_U11 ( .A(rout_y[61]), .B(p2[61]), .S(mux_y_n266), .Z(
        state_y[61]) );
  MUX2_X1 mux_y_U10 ( .A(rout_y[60]), .B(p2[60]), .S(mux_y_n266), .Z(
        state_y[60]) );
  MUX2_X1 mux_y_U9 ( .A(rout_y[29]), .B(p2[29]), .S(mux_y_n266), .Z(
        state_y[29]) );
  MUX2_X1 mux_y_U8 ( .A(rout_y[25]), .B(p2[41]), .S(mux_y_n266), .Z(
        state_y[25]) );
  MUX2_X1 mux_y_U7 ( .A(rout_y[15]), .B(p2[15]), .S(mux_y_n266), .Z(
        state_y[15]) );
  MUX2_X1 mux_y_U6 ( .A(rout_y[11]), .B(p2[27]), .S(mux_y_n266), .Z(
        state_y[11]) );
  MUX2_X1 mux_y_U5 ( .A(rout_y[7]), .B(p2[39]), .S(mux_y_n266), .Z(state_y[7])
         );
  MUX2_X1 mux_y_U4 ( .A(rout_y[6]), .B(p2[38]), .S(mux_y_n266), .Z(state_y[6])
         );
  INV_X1 mux_y_U3 ( .A(mux_y_n263), .ZN(mux_y_n266) );
  INV_X1 mux_y_U2 ( .A(start_sig), .ZN(mux_y_n263) );
  INV_X2 mux_y_U1 ( .A(mux_y_n263), .ZN(mux_y_n264) );
  MUX2_X1 mux_z_U68 ( .A(rout_z[34]), .B(p3[18]), .S(mux_z_n266), .Z(
        state_z[34]) );
  MUX2_X1 mux_z_U67 ( .A(rout_z[33]), .B(p3[17]), .S(mux_z_n265), .Z(
        state_z[33]) );
  MUX2_X1 mux_z_U66 ( .A(rout_z[30]), .B(p3[30]), .S(mux_z_n265), .Z(
        state_z[30]) );
  MUX2_X1 mux_z_U65 ( .A(rout_z[29]), .B(p3[29]), .S(mux_z_n264), .Z(
        state_z[29]) );
  MUX2_X1 mux_z_U64 ( .A(rout_z[28]), .B(p3[28]), .S(mux_z_n264), .Z(
        state_z[28]) );
  MUX2_X1 mux_z_U63 ( .A(rout_z[27]), .B(p3[43]), .S(mux_z_n264), .Z(
        state_z[27]) );
  MUX2_X1 mux_z_U62 ( .A(rout_z[26]), .B(p3[42]), .S(mux_z_n264), .Z(
        state_z[26]) );
  MUX2_X1 mux_z_U61 ( .A(rout_z[25]), .B(p3[41]), .S(mux_z_n264), .Z(
        state_z[25]) );
  MUX2_X1 mux_z_U60 ( .A(rout_z[24]), .B(p3[40]), .S(mux_z_n264), .Z(
        state_z[24]) );
  MUX2_X1 mux_z_U59 ( .A(rout_z[23]), .B(p3[55]), .S(mux_z_n264), .Z(
        state_z[23]) );
  MUX2_X1 mux_z_U58 ( .A(rout_z[21]), .B(p3[53]), .S(mux_z_n264), .Z(
        state_z[21]) );
  MUX2_X1 mux_z_U57 ( .A(rout_z[19]), .B(p3[3]), .S(mux_z_n264), .Z(
        state_z[19]) );
  MUX2_X1 mux_z_U56 ( .A(rout_z[18]), .B(p3[2]), .S(mux_z_n264), .Z(
        state_z[18]) );
  MUX2_X1 mux_z_U55 ( .A(rout_z[17]), .B(p3[1]), .S(mux_z_n264), .Z(
        state_z[17]) );
  MUX2_X1 mux_z_U54 ( .A(rout_z[15]), .B(p3[15]), .S(mux_z_n264), .Z(
        state_z[15]) );
  MUX2_X1 mux_z_U53 ( .A(rout_z[14]), .B(p3[14]), .S(mux_z_n264), .Z(
        state_z[14]) );
  MUX2_X1 mux_z_U52 ( .A(rout_z[13]), .B(p3[13]), .S(mux_z_n264), .Z(
        state_z[13]) );
  MUX2_X1 mux_z_U51 ( .A(rout_z[12]), .B(p3[12]), .S(mux_z_n264), .Z(
        state_z[12]) );
  MUX2_X1 mux_z_U50 ( .A(rout_z[11]), .B(p3[27]), .S(mux_z_n264), .Z(
        state_z[11]) );
  MUX2_X1 mux_z_U49 ( .A(rout_z[10]), .B(p3[26]), .S(mux_z_n264), .Z(
        state_z[10]) );
  MUX2_X1 mux_z_U48 ( .A(rout_z[9]), .B(p3[25]), .S(mux_z_n264), .Z(state_z[9]) );
  MUX2_X1 mux_z_U47 ( .A(rout_z[8]), .B(p3[24]), .S(mux_z_n264), .Z(state_z[8]) );
  MUX2_X1 mux_z_U46 ( .A(rout_z[7]), .B(p3[39]), .S(mux_z_n264), .Z(state_z[7]) );
  MUX2_X1 mux_z_U45 ( .A(rout_z[6]), .B(p3[38]), .S(mux_z_n266), .Z(state_z[6]) );
  MUX2_X1 mux_z_U44 ( .A(rout_z[5]), .B(p3[37]), .S(mux_z_n265), .Z(state_z[5]) );
  MUX2_X1 mux_z_U43 ( .A(rout_z[4]), .B(p3[36]), .S(mux_z_n266), .Z(state_z[4]) );
  MUX2_X1 mux_z_U42 ( .A(rout_z[3]), .B(p3[51]), .S(mux_z_n264), .Z(state_z[3]) );
  MUX2_X1 mux_z_U41 ( .A(rout_z[2]), .B(p3[50]), .S(mux_z_n264), .Z(state_z[2]) );
  MUX2_X1 mux_z_U40 ( .A(rout_z[0]), .B(p3[48]), .S(mux_z_n265), .Z(state_z[0]) );
  MUX2_X1 mux_z_U39 ( .A(rout_z[59]), .B(p3[11]), .S(mux_z_n264), .Z(
        state_z[59]) );
  MUX2_X1 mux_z_U38 ( .A(rout_z[58]), .B(p3[10]), .S(mux_z_n264), .Z(
        state_z[58]) );
  MUX2_X1 mux_z_U37 ( .A(rout_z[57]), .B(p3[9]), .S(mux_z_n266), .Z(
        state_z[57]) );
  MUX2_X1 mux_z_U36 ( .A(rout_z[56]), .B(p3[8]), .S(mux_z_n265), .Z(
        state_z[56]) );
  MUX2_X1 mux_z_U35 ( .A(rout_z[55]), .B(p3[23]), .S(mux_z_n264), .Z(
        state_z[55]) );
  MUX2_X1 mux_z_U34 ( .A(rout_z[54]), .B(p3[22]), .S(mux_z_n264), .Z(
        state_z[54]) );
  MUX2_X1 mux_z_U33 ( .A(rout_z[53]), .B(p3[21]), .S(mux_z_n266), .Z(
        state_z[53]) );
  MUX2_X1 mux_z_U32 ( .A(rout_z[52]), .B(p3[20]), .S(mux_z_n265), .Z(
        state_z[52]) );
  MUX2_X1 mux_z_U31 ( .A(rout_z[51]), .B(p3[35]), .S(mux_z_n264), .Z(
        state_z[51]) );
  MUX2_X1 mux_z_U30 ( .A(rout_z[50]), .B(p3[34]), .S(mux_z_n264), .Z(
        state_z[50]) );
  MUX2_X1 mux_z_U29 ( .A(rout_z[49]), .B(p3[33]), .S(mux_z_n266), .Z(
        state_z[49]) );
  MUX2_X1 mux_z_U28 ( .A(rout_z[48]), .B(p3[32]), .S(mux_z_n265), .Z(
        state_z[48]) );
  MUX2_X1 mux_z_U27 ( .A(rout_z[47]), .B(p3[47]), .S(mux_z_n265), .Z(
        state_z[47]) );
  MUX2_X1 mux_z_U26 ( .A(rout_z[46]), .B(p3[46]), .S(mux_z_n265), .Z(
        state_z[46]) );
  MUX2_X1 mux_z_U25 ( .A(rout_z[45]), .B(p3[45]), .S(mux_z_n265), .Z(
        state_z[45]) );
  MUX2_X1 mux_z_U24 ( .A(rout_z[44]), .B(p3[44]), .S(mux_z_n265), .Z(
        state_z[44]) );
  MUX2_X1 mux_z_U23 ( .A(rout_z[43]), .B(p3[59]), .S(mux_z_n265), .Z(
        state_z[43]) );
  MUX2_X1 mux_z_U22 ( .A(rout_z[42]), .B(p3[58]), .S(mux_z_n265), .Z(
        state_z[42]) );
  MUX2_X1 mux_z_U21 ( .A(rout_z[41]), .B(p3[57]), .S(mux_z_n265), .Z(
        state_z[41]) );
  MUX2_X1 mux_z_U20 ( .A(rout_z[40]), .B(p3[56]), .S(mux_z_n265), .Z(
        state_z[40]) );
  MUX2_X1 mux_z_U19 ( .A(rout_z[39]), .B(p3[7]), .S(mux_z_n265), .Z(
        state_z[39]) );
  MUX2_X1 mux_z_U18 ( .A(rout_z[38]), .B(p3[6]), .S(mux_z_n265), .Z(
        state_z[38]) );
  MUX2_X1 mux_z_U17 ( .A(rout_z[37]), .B(p3[5]), .S(mux_z_n265), .Z(
        state_z[37]) );
  INV_X1 mux_z_U16 ( .A(mux_z_n263), .ZN(mux_z_n265) );
  MUX2_X1 mux_z_U15 ( .A(rout_z[36]), .B(p3[4]), .S(mux_z_n266), .Z(
        state_z[36]) );
  MUX2_X1 mux_z_U14 ( .A(rout_z[63]), .B(p3[63]), .S(mux_z_n266), .Z(
        state_z[63]) );
  MUX2_X1 mux_z_U13 ( .A(rout_z[62]), .B(p3[62]), .S(mux_z_n266), .Z(
        state_z[62]) );
  MUX2_X1 mux_z_U12 ( .A(rout_z[61]), .B(p3[61]), .S(mux_z_n266), .Z(
        state_z[61]) );
  MUX2_X1 mux_z_U11 ( .A(rout_z[60]), .B(p3[60]), .S(mux_z_n266), .Z(
        state_z[60]) );
  MUX2_X1 mux_z_U10 ( .A(rout_z[35]), .B(p3[19]), .S(mux_z_n266), .Z(
        state_z[35]) );
  MUX2_X1 mux_z_U9 ( .A(rout_z[32]), .B(p3[16]), .S(mux_z_n266), .Z(
        state_z[32]) );
  MUX2_X1 mux_z_U8 ( .A(rout_z[31]), .B(p3[31]), .S(mux_z_n266), .Z(
        state_z[31]) );
  MUX2_X1 mux_z_U7 ( .A(rout_z[22]), .B(p3[54]), .S(mux_z_n266), .Z(
        state_z[22]) );
  MUX2_X1 mux_z_U6 ( .A(rout_z[20]), .B(p3[52]), .S(mux_z_n266), .Z(
        state_z[20]) );
  MUX2_X1 mux_z_U5 ( .A(rout_z[16]), .B(p3[0]), .S(mux_z_n266), .Z(state_z[16]) );
  MUX2_X1 mux_z_U4 ( .A(rout_z[1]), .B(p3[49]), .S(mux_z_n266), .Z(state_z[1])
         );
  INV_X1 mux_z_U3 ( .A(mux_z_n263), .ZN(mux_z_n266) );
  INV_X1 mux_z_U2 ( .A(start_sig), .ZN(mux_z_n263) );
  INV_X2 mux_z_U1 ( .A(mux_z_n263), .ZN(mux_z_n264) );
  MUX2_X1 mux_b_U4 ( .A(bout[3]), .B(b_guard[3]), .S(start_sig), .Z(state_b[3]) );
  MUX2_X1 mux_b_U3 ( .A(bout[2]), .B(b_guard[2]), .S(start_sig), .Z(state_b[2]) );
  MUX2_X1 mux_b_U2 ( .A(bout[1]), .B(b_guard[1]), .S(start_sig), .Z(state_b[1]) );
  MUX2_X1 mux_b_U1 ( .A(bout[0]), .B(b_guard[0]), .S(start_sig), .Z(state_b[0]) );
  MUX2_X1 mux_c_U4 ( .A(cout[2]), .B(c_guard[2]), .S(start_sig), .Z(state_c[2]) );
  MUX2_X1 mux_c_U3 ( .A(cout[1]), .B(c_guard[1]), .S(start_sig), .Z(state_c[1]) );
  MUX2_X1 mux_c_U2 ( .A(cout[0]), .B(c_guard[0]), .S(start_sig), .Z(state_c[0]) );
  MUX2_X1 mux_c_U1 ( .A(cout[3]), .B(c_guard[3]), .S(start_sig), .Z(state_c[3]) );
  MUX2_X1 mux_d_U4 ( .A(dout[3]), .B(d_guard[3]), .S(start_sig), .Z(state_d[3]) );
  MUX2_X1 mux_d_U3 ( .A(dout[2]), .B(d_guard[2]), .S(start_sig), .Z(state_d[2]) );
  MUX2_X1 mux_d_U2 ( .A(dout[1]), .B(d_guard[1]), .S(start_sig), .Z(state_d[1]) );
  MUX2_X1 mux_d_U1 ( .A(dout[0]), .B(d_guard[0]), .S(start_sig), .Z(state_d[0]) );
  NAND2_X1 reg_w_U204 ( .A1(reg_w_n339), .A2(reg_w_n338), .ZN(reg_w_n167) );
  NAND2_X1 reg_w_U203 ( .A1(state_w[35]), .A2(reg_w_n337), .ZN(reg_w_n338) );
  NAND2_X1 reg_w_U202 ( .A1(round_inst_srout_w[19]), .A2(reg_w_n336), .ZN(
        reg_w_n339) );
  NAND2_X1 reg_w_U201 ( .A1(reg_w_n335), .A2(reg_w_n334), .ZN(reg_w_n166) );
  NAND2_X1 reg_w_U200 ( .A1(state_w[34]), .A2(reg_w_n337), .ZN(reg_w_n334) );
  NAND2_X1 reg_w_U199 ( .A1(round_inst_aout_w[35]), .A2(reg_w_n336), .ZN(
        reg_w_n335) );
  NAND2_X1 reg_w_U198 ( .A1(reg_w_n333), .A2(reg_w_n332), .ZN(reg_w_n165) );
  NAND2_X1 reg_w_U197 ( .A1(state_w[33]), .A2(reg_w_n337), .ZN(reg_w_n332) );
  NAND2_X1 reg_w_U196 ( .A1(round_inst_srout_w[17]), .A2(reg_w_n336), .ZN(
        reg_w_n333) );
  NAND2_X1 reg_w_U195 ( .A1(reg_w_n331), .A2(reg_w_n330), .ZN(reg_w_n164) );
  NAND2_X1 reg_w_U194 ( .A1(state_w[32]), .A2(reg_w_n337), .ZN(reg_w_n330) );
  NAND2_X1 reg_w_U193 ( .A1(round_inst_srout_w[16]), .A2(reg_w_n336), .ZN(
        reg_w_n331) );
  NAND2_X1 reg_w_U192 ( .A1(reg_w_n329), .A2(reg_w_n328), .ZN(reg_w_n163) );
  NAND2_X1 reg_w_U191 ( .A1(state_w[31]), .A2(reg_w_n337), .ZN(reg_w_n328) );
  NAND2_X1 reg_w_U190 ( .A1(round_inst_srout_w[31]), .A2(reg_w_n336), .ZN(
        reg_w_n329) );
  NAND2_X1 reg_w_U189 ( .A1(reg_w_n327), .A2(reg_w_n326), .ZN(reg_w_n162) );
  NAND2_X1 reg_w_U188 ( .A1(state_w[30]), .A2(reg_w_n337), .ZN(reg_w_n326) );
  NAND2_X1 reg_w_U187 ( .A1(round_inst_aout_w[31]), .A2(reg_w_n336), .ZN(
        reg_w_n327) );
  NAND2_X1 reg_w_U186 ( .A1(reg_w_n325), .A2(reg_w_n324), .ZN(reg_w_n161) );
  NAND2_X1 reg_w_U185 ( .A1(state_w[29]), .A2(reg_w_n337), .ZN(reg_w_n324) );
  NAND2_X1 reg_w_U184 ( .A1(round_inst_srout_w[29]), .A2(reg_w_n336), .ZN(
        reg_w_n325) );
  NAND2_X1 reg_w_U183 ( .A1(reg_w_n323), .A2(reg_w_n322), .ZN(reg_w_n160) );
  NAND2_X1 reg_w_U182 ( .A1(state_w[28]), .A2(reg_w_n337), .ZN(reg_w_n322) );
  NAND2_X1 reg_w_U181 ( .A1(round_inst_srout_w[28]), .A2(reg_w_n336), .ZN(
        reg_w_n323) );
  NAND2_X1 reg_w_U180 ( .A1(reg_w_n321), .A2(reg_w_n320), .ZN(reg_w_n159) );
  NAND2_X1 reg_w_U179 ( .A1(state_w[27]), .A2(reg_w_n337), .ZN(reg_w_n320) );
  NAND2_X1 reg_w_U178 ( .A1(round_inst_srout_w[43]), .A2(reg_w_n336), .ZN(
        reg_w_n321) );
  NAND2_X1 reg_w_U177 ( .A1(reg_w_n319), .A2(reg_w_n318), .ZN(reg_w_n158) );
  NAND2_X1 reg_w_U176 ( .A1(state_w[26]), .A2(reg_w_n337), .ZN(reg_w_n318) );
  NAND2_X1 reg_w_U175 ( .A1(round_inst_aout_w[27]), .A2(reg_w_n336), .ZN(
        reg_w_n319) );
  NAND2_X1 reg_w_U174 ( .A1(reg_w_n317), .A2(reg_w_n316), .ZN(reg_w_n157) );
  NAND2_X1 reg_w_U173 ( .A1(state_w[25]), .A2(reg_w_n337), .ZN(reg_w_n316) );
  NAND2_X1 reg_w_U172 ( .A1(round_inst_srout_w[41]), .A2(reg_w_n336), .ZN(
        reg_w_n317) );
  NAND2_X1 reg_w_U171 ( .A1(reg_w_n315), .A2(reg_w_n314), .ZN(reg_w_n156) );
  NAND2_X1 reg_w_U170 ( .A1(state_w[24]), .A2(reg_w_n337), .ZN(reg_w_n314) );
  NAND2_X1 reg_w_U169 ( .A1(round_inst_srout_w[40]), .A2(reg_w_n336), .ZN(
        reg_w_n315) );
  NAND2_X1 reg_w_U168 ( .A1(reg_w_n313), .A2(reg_w_n312), .ZN(reg_w_n155) );
  NAND2_X1 reg_w_U167 ( .A1(state_w[23]), .A2(reg_w_n229), .ZN(reg_w_n312) );
  NAND2_X1 reg_w_U166 ( .A1(round_inst_srout_w[55]), .A2(reg_w_n311), .ZN(
        reg_w_n313) );
  NAND2_X1 reg_w_U165 ( .A1(reg_w_n310), .A2(reg_w_n309), .ZN(reg_w_n154) );
  NAND2_X1 reg_w_U164 ( .A1(state_w[22]), .A2(reg_w_n229), .ZN(reg_w_n309) );
  NAND2_X1 reg_w_U163 ( .A1(round_inst_aout_w[23]), .A2(reg_w_n311), .ZN(
        reg_w_n310) );
  NAND2_X1 reg_w_U162 ( .A1(reg_w_n308), .A2(reg_w_n307), .ZN(reg_w_n153) );
  NAND2_X1 reg_w_U161 ( .A1(state_w[21]), .A2(reg_w_n229), .ZN(reg_w_n307) );
  NAND2_X1 reg_w_U160 ( .A1(round_inst_srout_w[53]), .A2(reg_w_n311), .ZN(
        reg_w_n308) );
  NAND2_X1 reg_w_U159 ( .A1(reg_w_n306), .A2(reg_w_n305), .ZN(reg_w_n152) );
  NAND2_X1 reg_w_U158 ( .A1(state_w[20]), .A2(reg_w_n229), .ZN(reg_w_n305) );
  NAND2_X1 reg_w_U157 ( .A1(round_inst_srout_w[52]), .A2(reg_w_n311), .ZN(
        reg_w_n306) );
  NAND2_X1 reg_w_U156 ( .A1(reg_w_n304), .A2(reg_w_n303), .ZN(reg_w_n151) );
  NAND2_X1 reg_w_U155 ( .A1(state_w[19]), .A2(reg_w_n229), .ZN(reg_w_n303) );
  NAND2_X1 reg_w_U154 ( .A1(round_inst_srout_w[3]), .A2(reg_w_n311), .ZN(
        reg_w_n304) );
  NAND2_X1 reg_w_U153 ( .A1(reg_w_n302), .A2(reg_w_n301), .ZN(reg_w_n150) );
  NAND2_X1 reg_w_U152 ( .A1(state_w[18]), .A2(reg_w_n229), .ZN(reg_w_n301) );
  NAND2_X1 reg_w_U151 ( .A1(round_inst_aout_w[19]), .A2(reg_w_n311), .ZN(
        reg_w_n302) );
  NAND2_X1 reg_w_U150 ( .A1(reg_w_n300), .A2(reg_w_n299), .ZN(reg_w_n149) );
  NAND2_X1 reg_w_U149 ( .A1(state_w[17]), .A2(reg_w_n229), .ZN(reg_w_n299) );
  NAND2_X1 reg_w_U148 ( .A1(round_inst_srout_w[1]), .A2(reg_w_n311), .ZN(
        reg_w_n300) );
  NAND2_X1 reg_w_U147 ( .A1(reg_w_n298), .A2(reg_w_n297), .ZN(reg_w_n148) );
  NAND2_X1 reg_w_U146 ( .A1(state_w[16]), .A2(reg_w_n229), .ZN(reg_w_n297) );
  NAND2_X1 reg_w_U145 ( .A1(round_inst_srout_w[0]), .A2(reg_w_n311), .ZN(
        reg_w_n298) );
  NAND2_X1 reg_w_U144 ( .A1(reg_w_n296), .A2(reg_w_n295), .ZN(reg_w_n147) );
  NAND2_X1 reg_w_U143 ( .A1(state_w[15]), .A2(reg_w_n229), .ZN(reg_w_n295) );
  NAND2_X1 reg_w_U142 ( .A1(round_inst_srout_w[15]), .A2(reg_w_n311), .ZN(
        reg_w_n296) );
  NAND2_X1 reg_w_U141 ( .A1(reg_w_n294), .A2(reg_w_n293), .ZN(reg_w_n146) );
  NAND2_X1 reg_w_U140 ( .A1(state_w[14]), .A2(reg_w_n229), .ZN(reg_w_n293) );
  NAND2_X1 reg_w_U139 ( .A1(round_inst_aout_w[15]), .A2(reg_w_n311), .ZN(
        reg_w_n294) );
  NAND2_X1 reg_w_U138 ( .A1(reg_w_n292), .A2(reg_w_n291), .ZN(reg_w_n145) );
  NAND2_X1 reg_w_U137 ( .A1(state_w[13]), .A2(reg_w_n229), .ZN(reg_w_n291) );
  NAND2_X1 reg_w_U136 ( .A1(round_inst_srout_w[13]), .A2(reg_w_n311), .ZN(
        reg_w_n292) );
  NAND2_X1 reg_w_U135 ( .A1(reg_w_n290), .A2(reg_w_n289), .ZN(reg_w_n144) );
  NAND2_X1 reg_w_U134 ( .A1(state_w[12]), .A2(reg_w_n229), .ZN(reg_w_n289) );
  NAND2_X1 reg_w_U133 ( .A1(round_inst_srout_w[12]), .A2(reg_w_n311), .ZN(
        reg_w_n290) );
  NAND2_X1 reg_w_U132 ( .A1(reg_w_n288), .A2(reg_w_n287), .ZN(reg_w_n143) );
  NAND2_X1 reg_w_U131 ( .A1(state_w[11]), .A2(reg_w_n229), .ZN(reg_w_n287) );
  NAND2_X1 reg_w_U130 ( .A1(round_inst_srout_w[27]), .A2(reg_w_n311), .ZN(
        reg_w_n288) );
  NAND2_X1 reg_w_U129 ( .A1(reg_w_n286), .A2(reg_w_n285), .ZN(reg_w_n142) );
  NAND2_X1 reg_w_U128 ( .A1(state_w[10]), .A2(reg_w_n337), .ZN(reg_w_n285) );
  NAND2_X1 reg_w_U127 ( .A1(round_inst_aout_w[11]), .A2(reg_w_n336), .ZN(
        reg_w_n286) );
  NAND2_X1 reg_w_U126 ( .A1(reg_w_n284), .A2(reg_w_n283), .ZN(reg_w_n141) );
  NAND2_X1 reg_w_U125 ( .A1(state_w[9]), .A2(reg_w_n229), .ZN(reg_w_n283) );
  NAND2_X1 reg_w_U124 ( .A1(round_inst_srout_w[25]), .A2(reg_w_n311), .ZN(
        reg_w_n284) );
  NAND2_X1 reg_w_U123 ( .A1(reg_w_n282), .A2(reg_w_n281), .ZN(reg_w_n140) );
  NAND2_X1 reg_w_U122 ( .A1(state_w[8]), .A2(reg_w_n337), .ZN(reg_w_n281) );
  NAND2_X1 reg_w_U121 ( .A1(round_inst_srout_w[24]), .A2(reg_w_n336), .ZN(
        reg_w_n282) );
  NAND2_X1 reg_w_U120 ( .A1(reg_w_n280), .A2(reg_w_n279), .ZN(reg_w_n139) );
  NAND2_X1 reg_w_U119 ( .A1(state_w[7]), .A2(reg_w_n229), .ZN(reg_w_n279) );
  NAND2_X1 reg_w_U118 ( .A1(round_inst_srout_w[39]), .A2(reg_w_n311), .ZN(
        reg_w_n280) );
  NAND2_X1 reg_w_U117 ( .A1(reg_w_n278), .A2(reg_w_n277), .ZN(reg_w_n136) );
  NAND2_X1 reg_w_U116 ( .A1(state_w[4]), .A2(reg_w_n337), .ZN(reg_w_n277) );
  NAND2_X1 reg_w_U115 ( .A1(round_inst_srout_w[36]), .A2(reg_w_n336), .ZN(
        reg_w_n278) );
  NAND2_X1 reg_w_U114 ( .A1(reg_w_n276), .A2(reg_w_n275), .ZN(reg_w_n135) );
  NAND2_X1 reg_w_U113 ( .A1(state_w[3]), .A2(reg_w_n229), .ZN(reg_w_n275) );
  NAND2_X1 reg_w_U112 ( .A1(round_inst_srout_w[51]), .A2(reg_w_n311), .ZN(
        reg_w_n276) );
  NAND2_X1 reg_w_U111 ( .A1(reg_w_n274), .A2(reg_w_n273), .ZN(reg_w_n134) );
  NAND2_X1 reg_w_U110 ( .A1(state_w[2]), .A2(reg_w_n337), .ZN(reg_w_n273) );
  NAND2_X1 reg_w_U109 ( .A1(round_inst_aout_w[3]), .A2(reg_w_n336), .ZN(
        reg_w_n274) );
  NAND2_X1 reg_w_U108 ( .A1(reg_w_n272), .A2(reg_w_n271), .ZN(reg_w_n133) );
  NAND2_X1 reg_w_U107 ( .A1(state_w[1]), .A2(reg_w_n337), .ZN(reg_w_n271) );
  NAND2_X1 reg_w_U106 ( .A1(round_inst_srout_w[49]), .A2(reg_w_n311), .ZN(
        reg_w_n272) );
  INV_X1 reg_w_U105 ( .A(reg_w_n270), .ZN(reg_w_n311) );
  NAND2_X1 reg_w_U104 ( .A1(reg_w_n269), .A2(reg_w_n268), .ZN(reg_w_n132) );
  NAND2_X1 reg_w_U103 ( .A1(state_w[0]), .A2(reg_w_n337), .ZN(reg_w_n268) );
  NAND2_X1 reg_w_U102 ( .A1(round_inst_srout_w[48]), .A2(reg_w_n336), .ZN(
        reg_w_n269) );
  INV_X1 reg_w_U101 ( .A(reg_w_n270), .ZN(reg_w_n336) );
  NAND2_X1 reg_w_U100 ( .A1(reg_w_n267), .A2(reg_w_n266), .ZN(reg_w_n191) );
  NAND2_X1 reg_w_U99 ( .A1(state_w[59]), .A2(reg_w_n229), .ZN(reg_w_n266) );
  NAND2_X1 reg_w_U98 ( .A1(round_inst_srout_w[11]), .A2(reg_w_n264), .ZN(
        reg_w_n267) );
  NAND2_X1 reg_w_U97 ( .A1(reg_w_n263), .A2(reg_w_n262), .ZN(reg_w_n190) );
  NAND2_X1 reg_w_U96 ( .A1(state_w[58]), .A2(reg_w_n337), .ZN(reg_w_n262) );
  INV_X1 reg_w_U95 ( .A(reg_w_n265), .ZN(reg_w_n337) );
  NAND2_X1 reg_w_U94 ( .A1(round_inst_aout_w[59]), .A2(reg_w_n264), .ZN(
        reg_w_n263) );
  NAND2_X1 reg_w_U93 ( .A1(reg_w_n261), .A2(reg_w_n260), .ZN(reg_w_n189) );
  NAND2_X1 reg_w_U92 ( .A1(state_w[57]), .A2(reg_w_n259), .ZN(reg_w_n260) );
  NAND2_X1 reg_w_U91 ( .A1(round_inst_srout_w[9]), .A2(reg_w_n264), .ZN(
        reg_w_n261) );
  NAND2_X1 reg_w_U90 ( .A1(reg_w_n258), .A2(reg_w_n257), .ZN(reg_w_n188) );
  NAND2_X1 reg_w_U89 ( .A1(state_w[56]), .A2(reg_w_n259), .ZN(reg_w_n257) );
  NAND2_X1 reg_w_U88 ( .A1(round_inst_srout_w[8]), .A2(reg_w_n264), .ZN(
        reg_w_n258) );
  NAND2_X1 reg_w_U87 ( .A1(reg_w_n256), .A2(reg_w_n255), .ZN(reg_w_n187) );
  NAND2_X1 reg_w_U86 ( .A1(state_w[55]), .A2(reg_w_n259), .ZN(reg_w_n255) );
  NAND2_X1 reg_w_U85 ( .A1(round_inst_srout_w[23]), .A2(reg_w_n264), .ZN(
        reg_w_n256) );
  NAND2_X1 reg_w_U84 ( .A1(reg_w_n254), .A2(reg_w_n253), .ZN(reg_w_n186) );
  NAND2_X1 reg_w_U83 ( .A1(state_w[54]), .A2(reg_w_n259), .ZN(reg_w_n253) );
  NAND2_X1 reg_w_U82 ( .A1(round_inst_aout_w[55]), .A2(reg_w_n264), .ZN(
        reg_w_n254) );
  NAND2_X1 reg_w_U81 ( .A1(reg_w_n252), .A2(reg_w_n251), .ZN(reg_w_n185) );
  NAND2_X1 reg_w_U80 ( .A1(state_w[53]), .A2(reg_w_n259), .ZN(reg_w_n251) );
  NAND2_X1 reg_w_U79 ( .A1(round_inst_srout_w[21]), .A2(reg_w_n264), .ZN(
        reg_w_n252) );
  NAND2_X1 reg_w_U78 ( .A1(reg_w_n250), .A2(reg_w_n249), .ZN(reg_w_n184) );
  NAND2_X1 reg_w_U77 ( .A1(state_w[52]), .A2(reg_w_n259), .ZN(reg_w_n249) );
  NAND2_X1 reg_w_U76 ( .A1(round_inst_srout_w[20]), .A2(reg_w_n248), .ZN(
        reg_w_n250) );
  NAND2_X1 reg_w_U75 ( .A1(reg_w_n247), .A2(reg_w_n246), .ZN(reg_w_n183) );
  NAND2_X1 reg_w_U74 ( .A1(state_w[51]), .A2(reg_w_n259), .ZN(reg_w_n246) );
  NAND2_X1 reg_w_U73 ( .A1(round_inst_srout_w[35]), .A2(reg_w_n248), .ZN(
        reg_w_n247) );
  NAND2_X1 reg_w_U72 ( .A1(reg_w_n245), .A2(reg_w_n244), .ZN(reg_w_n182) );
  NAND2_X1 reg_w_U71 ( .A1(state_w[50]), .A2(reg_w_n259), .ZN(reg_w_n244) );
  NAND2_X1 reg_w_U70 ( .A1(round_inst_aout_w[51]), .A2(reg_w_n248), .ZN(
        reg_w_n245) );
  NAND2_X1 reg_w_U69 ( .A1(reg_w_n243), .A2(reg_w_n242), .ZN(reg_w_n181) );
  NAND2_X1 reg_w_U68 ( .A1(state_w[49]), .A2(reg_w_n259), .ZN(reg_w_n242) );
  NAND2_X1 reg_w_U67 ( .A1(round_inst_srout_w[33]), .A2(reg_w_n248), .ZN(
        reg_w_n243) );
  NAND2_X1 reg_w_U66 ( .A1(reg_w_n241), .A2(reg_w_n240), .ZN(reg_w_n180) );
  NAND2_X1 reg_w_U65 ( .A1(state_w[48]), .A2(reg_w_n259), .ZN(reg_w_n240) );
  NAND2_X1 reg_w_U64 ( .A1(round_inst_srout_w[32]), .A2(reg_w_n248), .ZN(
        reg_w_n241) );
  NAND2_X1 reg_w_U63 ( .A1(reg_w_n239), .A2(reg_w_n238), .ZN(reg_w_n179) );
  NAND2_X1 reg_w_U62 ( .A1(state_w[47]), .A2(reg_w_n259), .ZN(reg_w_n238) );
  NAND2_X1 reg_w_U61 ( .A1(round_inst_srout_w[47]), .A2(reg_w_n248), .ZN(
        reg_w_n239) );
  NAND2_X1 reg_w_U60 ( .A1(reg_w_n237), .A2(reg_w_n236), .ZN(reg_w_n178) );
  NAND2_X1 reg_w_U59 ( .A1(state_w[46]), .A2(reg_w_n259), .ZN(reg_w_n236) );
  NAND2_X1 reg_w_U58 ( .A1(round_inst_aout_w[47]), .A2(reg_w_n248), .ZN(
        reg_w_n237) );
  NAND2_X1 reg_w_U57 ( .A1(reg_w_n235), .A2(reg_w_n234), .ZN(reg_w_n177) );
  NAND2_X1 reg_w_U56 ( .A1(state_w[45]), .A2(reg_w_n259), .ZN(reg_w_n234) );
  NAND2_X1 reg_w_U55 ( .A1(round_inst_srout_w[45]), .A2(reg_w_n248), .ZN(
        reg_w_n235) );
  NAND2_X1 reg_w_U54 ( .A1(reg_w_n233), .A2(reg_w_n232), .ZN(reg_w_n176) );
  NAND2_X1 reg_w_U53 ( .A1(state_w[44]), .A2(reg_w_n259), .ZN(reg_w_n232) );
  NAND2_X1 reg_w_U52 ( .A1(round_inst_srout_w[44]), .A2(reg_w_n248), .ZN(
        reg_w_n233) );
  NAND2_X1 reg_w_U51 ( .A1(reg_w_n231), .A2(reg_w_n230), .ZN(reg_w_n175) );
  NAND2_X1 reg_w_U50 ( .A1(state_w[43]), .A2(reg_w_n229), .ZN(reg_w_n230) );
  NAND2_X1 reg_w_U49 ( .A1(round_inst_srout_w[59]), .A2(reg_w_n248), .ZN(
        reg_w_n231) );
  NAND2_X1 reg_w_U48 ( .A1(reg_w_n228), .A2(reg_w_n227), .ZN(reg_w_n174) );
  NAND2_X1 reg_w_U47 ( .A1(state_w[42]), .A2(reg_w_n229), .ZN(reg_w_n227) );
  NAND2_X1 reg_w_U46 ( .A1(round_inst_aout_w[43]), .A2(reg_w_n248), .ZN(
        reg_w_n228) );
  NAND2_X1 reg_w_U45 ( .A1(reg_w_n226), .A2(reg_w_n225), .ZN(reg_w_n173) );
  NAND2_X1 reg_w_U44 ( .A1(state_w[41]), .A2(reg_w_n229), .ZN(reg_w_n225) );
  NAND2_X1 reg_w_U43 ( .A1(round_inst_srout_w[57]), .A2(reg_w_n248), .ZN(
        reg_w_n226) );
  NAND2_X1 reg_w_U42 ( .A1(reg_w_n224), .A2(reg_w_n223), .ZN(reg_w_n172) );
  NAND2_X1 reg_w_U41 ( .A1(state_w[40]), .A2(reg_w_n229), .ZN(reg_w_n223) );
  NAND2_X1 reg_w_U40 ( .A1(round_inst_srout_w[56]), .A2(reg_w_n248), .ZN(
        reg_w_n224) );
  NAND2_X1 reg_w_U39 ( .A1(reg_w_n222), .A2(reg_w_n221), .ZN(reg_w_n171) );
  NAND2_X1 reg_w_U38 ( .A1(state_w[39]), .A2(reg_w_n229), .ZN(reg_w_n221) );
  NAND2_X1 reg_w_U37 ( .A1(round_inst_srout_w[7]), .A2(reg_w_n248), .ZN(
        reg_w_n222) );
  NAND2_X1 reg_w_U36 ( .A1(reg_w_n220), .A2(reg_w_n219), .ZN(reg_w_n170) );
  NAND2_X1 reg_w_U35 ( .A1(state_w[38]), .A2(reg_w_n229), .ZN(reg_w_n219) );
  NAND2_X1 reg_w_U34 ( .A1(round_inst_aout_w[39]), .A2(reg_w_n248), .ZN(
        reg_w_n220) );
  NAND2_X1 reg_w_U33 ( .A1(reg_w_n218), .A2(reg_w_n217), .ZN(reg_w_n169) );
  NAND2_X1 reg_w_U32 ( .A1(state_w[37]), .A2(reg_w_n229), .ZN(reg_w_n217) );
  NAND2_X1 reg_w_U31 ( .A1(round_inst_srout_w[5]), .A2(reg_w_n248), .ZN(
        reg_w_n218) );
  NAND2_X1 reg_w_U30 ( .A1(reg_w_n216), .A2(reg_w_n215), .ZN(reg_w_n168) );
  NAND2_X1 reg_w_U29 ( .A1(state_w[36]), .A2(reg_w_n229), .ZN(reg_w_n215) );
  NAND2_X1 reg_w_U28 ( .A1(round_inst_srout_w[4]), .A2(reg_w_n248), .ZN(
        reg_w_n216) );
  NAND2_X1 reg_w_U27 ( .A1(reg_w_n214), .A2(reg_w_n213), .ZN(reg_w_n195) );
  NAND2_X1 reg_w_U26 ( .A1(state_w[63]), .A2(reg_w_n229), .ZN(reg_w_n213) );
  NAND2_X1 reg_w_U25 ( .A1(round_inst_srout_w[63]), .A2(reg_w_n248), .ZN(
        reg_w_n214) );
  NAND2_X1 reg_w_U24 ( .A1(reg_w_n212), .A2(reg_w_n211), .ZN(reg_w_n194) );
  NAND2_X1 reg_w_U23 ( .A1(state_w[62]), .A2(reg_w_n259), .ZN(reg_w_n211) );
  NAND2_X1 reg_w_U22 ( .A1(round_inst_aout_w[63]), .A2(reg_w_n248), .ZN(
        reg_w_n212) );
  NAND2_X1 reg_w_U21 ( .A1(reg_w_n210), .A2(reg_w_n209), .ZN(reg_w_n193) );
  NAND2_X1 reg_w_U20 ( .A1(state_w[61]), .A2(reg_w_n259), .ZN(reg_w_n209) );
  NAND2_X1 reg_w_U19 ( .A1(round_inst_srout_w[61]), .A2(reg_w_n264), .ZN(
        reg_w_n210) );
  NAND2_X1 reg_w_U18 ( .A1(reg_w_n208), .A2(reg_w_n207), .ZN(reg_w_n192) );
  NAND2_X1 reg_w_U17 ( .A1(state_w[60]), .A2(reg_w_n259), .ZN(reg_w_n207) );
  NAND2_X1 reg_w_U16 ( .A1(round_inst_srout_w[60]), .A2(reg_w_n248), .ZN(
        reg_w_n208) );
  NAND2_X1 reg_w_U15 ( .A1(reg_w_n206), .A2(reg_w_n205), .ZN(reg_w_n138) );
  NAND2_X1 reg_w_U14 ( .A1(state_w[6]), .A2(reg_w_n259), .ZN(reg_w_n205) );
  NAND2_X1 reg_w_U13 ( .A1(round_inst_aout_w[7]), .A2(reg_w_n264), .ZN(
        reg_w_n206) );
  NAND2_X1 reg_w_U12 ( .A1(reg_w_n204), .A2(reg_w_n203), .ZN(reg_w_n137) );
  NAND2_X1 reg_w_U11 ( .A1(reg_w_n248), .A2(round_inst_srout_w[37]), .ZN(
        reg_w_n203) );
  INV_X1 reg_w_U10 ( .A(reg_w_n270), .ZN(reg_w_n248) );
  INV_X1 reg_w_U9 ( .A(reg_w_n264), .ZN(reg_w_n270) );
  NAND2_X1 reg_w_U8 ( .A1(reg_w_n259), .A2(state_w[5]), .ZN(reg_w_n204) );
  INV_X1 reg_w_U7 ( .A(reg_w_n265), .ZN(reg_w_n259) );
  INV_X1 reg_w_U6 ( .A(reg_w_n229), .ZN(reg_w_n265) );
  NOR2_X4 reg_w_U5 ( .A1(rst), .A2(reg_w_n202), .ZN(reg_w_n229) );
  INV_X1 reg_w_U4 ( .A(en_sig), .ZN(reg_w_n202) );
  NOR2_X1 reg_w_U3 ( .A1(rst), .A2(en_sig), .ZN(reg_w_n264) );
  DFF_X1 reg_w_s_current_state_reg_0_ ( .D(reg_w_n132), .CK(clk), .Q(
        round_inst_srout_w[48]) );
  DFF_X1 reg_w_s_current_state_reg_1_ ( .D(reg_w_n133), .CK(clk), .Q(
        round_inst_srout_w[49]) );
  DFF_X1 reg_w_s_current_state_reg_2_ ( .D(reg_w_n134), .CK(clk), .Q(
        round_inst_aout_w[3]) );
  DFF_X1 reg_w_s_current_state_reg_3_ ( .D(reg_w_n135), .CK(clk), .Q(
        round_inst_srout_w[51]) );
  DFF_X1 reg_w_s_current_state_reg_4_ ( .D(reg_w_n136), .CK(clk), .Q(
        round_inst_srout_w[36]) );
  DFF_X1 reg_w_s_current_state_reg_5_ ( .D(reg_w_n137), .CK(clk), .Q(
        round_inst_srout_w[37]) );
  DFF_X1 reg_w_s_current_state_reg_6_ ( .D(reg_w_n138), .CK(clk), .Q(
        round_inst_aout_w[7]) );
  DFF_X1 reg_w_s_current_state_reg_7_ ( .D(reg_w_n139), .CK(clk), .Q(
        round_inst_srout_w[39]) );
  DFF_X1 reg_w_s_current_state_reg_8_ ( .D(reg_w_n140), .CK(clk), .Q(
        round_inst_srout_w[24]) );
  DFF_X1 reg_w_s_current_state_reg_9_ ( .D(reg_w_n141), .CK(clk), .Q(
        round_inst_srout_w[25]) );
  DFF_X1 reg_w_s_current_state_reg_10_ ( .D(reg_w_n142), .CK(clk), .Q(
        round_inst_aout_w[11]) );
  DFF_X1 reg_w_s_current_state_reg_11_ ( .D(reg_w_n143), .CK(clk), .Q(
        round_inst_srout_w[27]) );
  DFF_X1 reg_w_s_current_state_reg_12_ ( .D(reg_w_n144), .CK(clk), .Q(
        round_inst_srout_w[12]) );
  DFF_X1 reg_w_s_current_state_reg_13_ ( .D(reg_w_n145), .CK(clk), .Q(
        round_inst_srout_w[13]) );
  DFF_X1 reg_w_s_current_state_reg_14_ ( .D(reg_w_n146), .CK(clk), .Q(
        round_inst_aout_w[15]) );
  DFF_X1 reg_w_s_current_state_reg_15_ ( .D(reg_w_n147), .CK(clk), .Q(
        round_inst_srout_w[15]) );
  DFF_X1 reg_w_s_current_state_reg_16_ ( .D(reg_w_n148), .CK(clk), .Q(
        round_inst_srout_w[0]) );
  DFF_X1 reg_w_s_current_state_reg_17_ ( .D(reg_w_n149), .CK(clk), .Q(
        round_inst_srout_w[1]) );
  DFF_X1 reg_w_s_current_state_reg_18_ ( .D(reg_w_n150), .CK(clk), .Q(
        round_inst_aout_w[19]) );
  DFF_X1 reg_w_s_current_state_reg_19_ ( .D(reg_w_n151), .CK(clk), .Q(
        round_inst_srout_w[3]) );
  DFF_X1 reg_w_s_current_state_reg_20_ ( .D(reg_w_n152), .CK(clk), .Q(
        round_inst_srout_w[52]) );
  DFF_X1 reg_w_s_current_state_reg_21_ ( .D(reg_w_n153), .CK(clk), .Q(
        round_inst_srout_w[53]) );
  DFF_X1 reg_w_s_current_state_reg_22_ ( .D(reg_w_n154), .CK(clk), .Q(
        round_inst_aout_w[23]) );
  DFF_X1 reg_w_s_current_state_reg_23_ ( .D(reg_w_n155), .CK(clk), .Q(
        round_inst_srout_w[55]) );
  DFF_X1 reg_w_s_current_state_reg_24_ ( .D(reg_w_n156), .CK(clk), .Q(
        round_inst_srout_w[40]) );
  DFF_X1 reg_w_s_current_state_reg_25_ ( .D(reg_w_n157), .CK(clk), .Q(
        round_inst_srout_w[41]) );
  DFF_X1 reg_w_s_current_state_reg_26_ ( .D(reg_w_n158), .CK(clk), .Q(
        round_inst_aout_w[27]) );
  DFF_X1 reg_w_s_current_state_reg_27_ ( .D(reg_w_n159), .CK(clk), .Q(
        round_inst_srout_w[43]) );
  DFF_X1 reg_w_s_current_state_reg_28_ ( .D(reg_w_n160), .CK(clk), .Q(
        round_inst_srout_w[28]) );
  DFF_X1 reg_w_s_current_state_reg_29_ ( .D(reg_w_n161), .CK(clk), .Q(
        round_inst_srout_w[29]) );
  DFF_X1 reg_w_s_current_state_reg_30_ ( .D(reg_w_n162), .CK(clk), .Q(
        round_inst_aout_w[31]) );
  DFF_X1 reg_w_s_current_state_reg_31_ ( .D(reg_w_n163), .CK(clk), .Q(
        round_inst_srout_w[31]) );
  DFF_X1 reg_w_s_current_state_reg_32_ ( .D(reg_w_n164), .CK(clk), .Q(
        round_inst_srout_w[16]) );
  DFF_X1 reg_w_s_current_state_reg_33_ ( .D(reg_w_n165), .CK(clk), .Q(
        round_inst_srout_w[17]) );
  DFF_X1 reg_w_s_current_state_reg_34_ ( .D(reg_w_n166), .CK(clk), .Q(
        round_inst_aout_w[35]) );
  DFF_X1 reg_w_s_current_state_reg_35_ ( .D(reg_w_n167), .CK(clk), .Q(
        round_inst_srout_w[19]) );
  DFF_X1 reg_w_s_current_state_reg_36_ ( .D(reg_w_n168), .CK(clk), .Q(
        round_inst_srout_w[4]) );
  DFF_X1 reg_w_s_current_state_reg_37_ ( .D(reg_w_n169), .CK(clk), .Q(
        round_inst_srout_w[5]) );
  DFF_X1 reg_w_s_current_state_reg_38_ ( .D(reg_w_n170), .CK(clk), .Q(
        round_inst_aout_w[39]) );
  DFF_X1 reg_w_s_current_state_reg_39_ ( .D(reg_w_n171), .CK(clk), .Q(
        round_inst_srout_w[7]) );
  DFF_X1 reg_w_s_current_state_reg_40_ ( .D(reg_w_n172), .CK(clk), .Q(
        round_inst_srout_w[56]) );
  DFF_X1 reg_w_s_current_state_reg_41_ ( .D(reg_w_n173), .CK(clk), .Q(
        round_inst_srout_w[57]) );
  DFF_X1 reg_w_s_current_state_reg_42_ ( .D(reg_w_n174), .CK(clk), .Q(
        round_inst_aout_w[43]) );
  DFF_X1 reg_w_s_current_state_reg_43_ ( .D(reg_w_n175), .CK(clk), .Q(
        round_inst_srout_w[59]) );
  DFF_X1 reg_w_s_current_state_reg_44_ ( .D(reg_w_n176), .CK(clk), .Q(
        round_inst_srout_w[44]) );
  DFF_X1 reg_w_s_current_state_reg_45_ ( .D(reg_w_n177), .CK(clk), .Q(
        round_inst_srout_w[45]) );
  DFF_X1 reg_w_s_current_state_reg_46_ ( .D(reg_w_n178), .CK(clk), .Q(
        round_inst_aout_w[47]) );
  DFF_X1 reg_w_s_current_state_reg_47_ ( .D(reg_w_n179), .CK(clk), .Q(
        round_inst_srout_w[47]) );
  DFF_X1 reg_w_s_current_state_reg_48_ ( .D(reg_w_n180), .CK(clk), .Q(
        round_inst_srout_w[32]) );
  DFF_X1 reg_w_s_current_state_reg_49_ ( .D(reg_w_n181), .CK(clk), .Q(
        round_inst_srout_w[33]) );
  DFF_X1 reg_w_s_current_state_reg_50_ ( .D(reg_w_n182), .CK(clk), .Q(
        round_inst_aout_w[51]) );
  DFF_X1 reg_w_s_current_state_reg_51_ ( .D(reg_w_n183), .CK(clk), .Q(
        round_inst_srout_w[35]) );
  DFF_X1 reg_w_s_current_state_reg_52_ ( .D(reg_w_n184), .CK(clk), .Q(
        round_inst_srout_w[20]) );
  DFF_X1 reg_w_s_current_state_reg_53_ ( .D(reg_w_n185), .CK(clk), .Q(
        round_inst_srout_w[21]) );
  DFF_X1 reg_w_s_current_state_reg_54_ ( .D(reg_w_n186), .CK(clk), .Q(
        round_inst_aout_w[55]) );
  DFF_X1 reg_w_s_current_state_reg_55_ ( .D(reg_w_n187), .CK(clk), .Q(
        round_inst_srout_w[23]) );
  DFF_X1 reg_w_s_current_state_reg_56_ ( .D(reg_w_n188), .CK(clk), .Q(
        round_inst_srout_w[8]) );
  DFF_X1 reg_w_s_current_state_reg_57_ ( .D(reg_w_n189), .CK(clk), .Q(
        round_inst_srout_w[9]) );
  DFF_X1 reg_w_s_current_state_reg_58_ ( .D(reg_w_n190), .CK(clk), .Q(
        round_inst_aout_w[59]) );
  DFF_X1 reg_w_s_current_state_reg_59_ ( .D(reg_w_n191), .CK(clk), .Q(
        round_inst_srout_w[11]) );
  DFF_X1 reg_w_s_current_state_reg_60_ ( .D(reg_w_n192), .CK(clk), .Q(
        round_inst_srout_w[60]) );
  DFF_X1 reg_w_s_current_state_reg_61_ ( .D(reg_w_n193), .CK(clk), .Q(
        round_inst_srout_w[61]) );
  DFF_X1 reg_w_s_current_state_reg_62_ ( .D(reg_w_n194), .CK(clk), .Q(
        round_inst_aout_w[63]) );
  DFF_X1 reg_w_s_current_state_reg_63_ ( .D(reg_w_n195), .CK(clk), .Q(
        round_inst_srout_w[63]) );
  NAND2_X1 reg_x_U205 ( .A1(reg_x_n532), .A2(reg_x_n531), .ZN(reg_x_n231) );
  NAND2_X1 reg_x_U204 ( .A1(state_x[34]), .A2(reg_x_n530), .ZN(reg_x_n531) );
  NAND2_X1 reg_x_U203 ( .A1(round_inst_aout_x[35]), .A2(reg_x_n529), .ZN(
        reg_x_n532) );
  NAND2_X1 reg_x_U202 ( .A1(reg_x_n528), .A2(reg_x_n527), .ZN(reg_x_n232) );
  NAND2_X1 reg_x_U201 ( .A1(state_x[33]), .A2(reg_x_n530), .ZN(reg_x_n527) );
  NAND2_X1 reg_x_U200 ( .A1(round_inst_aout_x[32]), .A2(reg_x_n529), .ZN(
        reg_x_n528) );
  NAND2_X1 reg_x_U199 ( .A1(reg_x_n526), .A2(reg_x_n525), .ZN(reg_x_n233) );
  NAND2_X1 reg_x_U198 ( .A1(state_x[32]), .A2(reg_x_n530), .ZN(reg_x_n525) );
  NAND2_X1 reg_x_U197 ( .A1(round_inst_srout_x[16]), .A2(reg_x_n529), .ZN(
        reg_x_n526) );
  NAND2_X1 reg_x_U196 ( .A1(reg_x_n524), .A2(reg_x_n523), .ZN(reg_x_n235) );
  NAND2_X1 reg_x_U195 ( .A1(state_x[30]), .A2(reg_x_n530), .ZN(reg_x_n523) );
  NAND2_X1 reg_x_U194 ( .A1(round_inst_aout_x[31]), .A2(reg_x_n529), .ZN(
        reg_x_n524) );
  NAND2_X1 reg_x_U193 ( .A1(reg_x_n522), .A2(reg_x_n521), .ZN(reg_x_n236) );
  NAND2_X1 reg_x_U192 ( .A1(state_x[29]), .A2(reg_x_n530), .ZN(reg_x_n521) );
  NAND2_X1 reg_x_U191 ( .A1(round_inst_aout_x[28]), .A2(reg_x_n529), .ZN(
        reg_x_n522) );
  NAND2_X1 reg_x_U190 ( .A1(reg_x_n520), .A2(reg_x_n519), .ZN(reg_x_n237) );
  NAND2_X1 reg_x_U189 ( .A1(state_x[28]), .A2(reg_x_n530), .ZN(reg_x_n519) );
  NAND2_X1 reg_x_U188 ( .A1(round_inst_srout_x[28]), .A2(reg_x_n529), .ZN(
        reg_x_n520) );
  NAND2_X1 reg_x_U187 ( .A1(reg_x_n518), .A2(reg_x_n517), .ZN(reg_x_n238) );
  NAND2_X1 reg_x_U186 ( .A1(state_x[27]), .A2(reg_x_n530), .ZN(reg_x_n517) );
  NAND2_X1 reg_x_U185 ( .A1(round_inst_aout_x[26]), .A2(reg_x_n529), .ZN(
        reg_x_n518) );
  NAND2_X1 reg_x_U184 ( .A1(reg_x_n516), .A2(reg_x_n515), .ZN(reg_x_n239) );
  NAND2_X1 reg_x_U183 ( .A1(state_x[26]), .A2(reg_x_n530), .ZN(reg_x_n515) );
  NAND2_X1 reg_x_U182 ( .A1(round_inst_aout_x[27]), .A2(reg_x_n529), .ZN(
        reg_x_n516) );
  NAND2_X1 reg_x_U181 ( .A1(reg_x_n514), .A2(reg_x_n513), .ZN(reg_x_n240) );
  NAND2_X1 reg_x_U180 ( .A1(state_x[25]), .A2(reg_x_n530), .ZN(reg_x_n513) );
  NAND2_X1 reg_x_U179 ( .A1(round_inst_aout_x[24]), .A2(reg_x_n529), .ZN(
        reg_x_n514) );
  NAND2_X1 reg_x_U178 ( .A1(reg_x_n512), .A2(reg_x_n511), .ZN(reg_x_n241) );
  NAND2_X1 reg_x_U177 ( .A1(state_x[24]), .A2(reg_x_n530), .ZN(reg_x_n511) );
  NAND2_X1 reg_x_U176 ( .A1(round_inst_srout_x[40]), .A2(reg_x_n529), .ZN(
        reg_x_n512) );
  NAND2_X1 reg_x_U175 ( .A1(reg_x_n510), .A2(reg_x_n509), .ZN(reg_x_n242) );
  NAND2_X1 reg_x_U174 ( .A1(state_x[23]), .A2(reg_x_n530), .ZN(reg_x_n509) );
  NAND2_X1 reg_x_U173 ( .A1(round_inst_aout_x[22]), .A2(reg_x_n529), .ZN(
        reg_x_n510) );
  NAND2_X1 reg_x_U172 ( .A1(reg_x_n508), .A2(reg_x_n507), .ZN(reg_x_n243) );
  NAND2_X1 reg_x_U171 ( .A1(state_x[22]), .A2(reg_x_n530), .ZN(reg_x_n507) );
  NAND2_X1 reg_x_U170 ( .A1(round_inst_aout_x[23]), .A2(reg_x_n529), .ZN(
        reg_x_n508) );
  NAND2_X1 reg_x_U169 ( .A1(reg_x_n506), .A2(reg_x_n505), .ZN(reg_x_n244) );
  NAND2_X1 reg_x_U168 ( .A1(state_x[21]), .A2(reg_x_n504), .ZN(reg_x_n505) );
  NAND2_X1 reg_x_U167 ( .A1(round_inst_aout_x[20]), .A2(reg_x_n503), .ZN(
        reg_x_n506) );
  NAND2_X1 reg_x_U166 ( .A1(reg_x_n502), .A2(reg_x_n501), .ZN(reg_x_n245) );
  NAND2_X1 reg_x_U165 ( .A1(state_x[20]), .A2(reg_x_n504), .ZN(reg_x_n501) );
  NAND2_X1 reg_x_U164 ( .A1(round_inst_srout_x[52]), .A2(reg_x_n503), .ZN(
        reg_x_n502) );
  NAND2_X1 reg_x_U163 ( .A1(reg_x_n500), .A2(reg_x_n499), .ZN(reg_x_n247) );
  NAND2_X1 reg_x_U162 ( .A1(state_x[18]), .A2(reg_x_n504), .ZN(reg_x_n499) );
  NAND2_X1 reg_x_U161 ( .A1(round_inst_aout_x[19]), .A2(reg_x_n503), .ZN(
        reg_x_n500) );
  NAND2_X1 reg_x_U160 ( .A1(reg_x_n498), .A2(reg_x_n497), .ZN(reg_x_n248) );
  NAND2_X1 reg_x_U159 ( .A1(state_x[17]), .A2(reg_x_n504), .ZN(reg_x_n497) );
  NAND2_X1 reg_x_U158 ( .A1(round_inst_aout_x[16]), .A2(reg_x_n503), .ZN(
        reg_x_n498) );
  NAND2_X1 reg_x_U157 ( .A1(reg_x_n496), .A2(reg_x_n495), .ZN(reg_x_n249) );
  NAND2_X1 reg_x_U156 ( .A1(state_x[16]), .A2(reg_x_n504), .ZN(reg_x_n495) );
  NAND2_X1 reg_x_U155 ( .A1(round_inst_srout_x[0]), .A2(reg_x_n503), .ZN(
        reg_x_n496) );
  NAND2_X1 reg_x_U154 ( .A1(reg_x_n494), .A2(reg_x_n493), .ZN(reg_x_n251) );
  NAND2_X1 reg_x_U153 ( .A1(state_x[14]), .A2(reg_x_n504), .ZN(reg_x_n493) );
  NAND2_X1 reg_x_U152 ( .A1(round_inst_aout_x[15]), .A2(reg_x_n503), .ZN(
        reg_x_n494) );
  NAND2_X1 reg_x_U151 ( .A1(reg_x_n492), .A2(reg_x_n491), .ZN(reg_x_n252) );
  NAND2_X1 reg_x_U150 ( .A1(state_x[13]), .A2(reg_x_n504), .ZN(reg_x_n491) );
  NAND2_X1 reg_x_U149 ( .A1(round_inst_aout_x[12]), .A2(reg_x_n503), .ZN(
        reg_x_n492) );
  NAND2_X1 reg_x_U148 ( .A1(reg_x_n490), .A2(reg_x_n489), .ZN(reg_x_n253) );
  NAND2_X1 reg_x_U147 ( .A1(state_x[12]), .A2(reg_x_n504), .ZN(reg_x_n489) );
  NAND2_X1 reg_x_U146 ( .A1(round_inst_srout_x[12]), .A2(reg_x_n503), .ZN(
        reg_x_n490) );
  NAND2_X1 reg_x_U145 ( .A1(reg_x_n488), .A2(reg_x_n487), .ZN(reg_x_n254) );
  NAND2_X1 reg_x_U144 ( .A1(state_x[11]), .A2(reg_x_n504), .ZN(reg_x_n487) );
  NAND2_X1 reg_x_U143 ( .A1(round_inst_aout_x[10]), .A2(reg_x_n503), .ZN(
        reg_x_n488) );
  NAND2_X1 reg_x_U142 ( .A1(reg_x_n486), .A2(reg_x_n485), .ZN(reg_x_n255) );
  NAND2_X1 reg_x_U141 ( .A1(state_x[10]), .A2(reg_x_n504), .ZN(reg_x_n485) );
  NAND2_X1 reg_x_U140 ( .A1(round_inst_aout_x[11]), .A2(reg_x_n503), .ZN(
        reg_x_n486) );
  NAND2_X1 reg_x_U139 ( .A1(reg_x_n484), .A2(reg_x_n483), .ZN(reg_x_n256) );
  NAND2_X1 reg_x_U138 ( .A1(state_x[9]), .A2(reg_x_n504), .ZN(reg_x_n483) );
  NAND2_X1 reg_x_U137 ( .A1(round_inst_aout_x[8]), .A2(reg_x_n503), .ZN(
        reg_x_n484) );
  NAND2_X1 reg_x_U136 ( .A1(reg_x_n482), .A2(reg_x_n481), .ZN(reg_x_n258) );
  NAND2_X1 reg_x_U135 ( .A1(state_x[7]), .A2(reg_x_n504), .ZN(reg_x_n481) );
  NAND2_X1 reg_x_U134 ( .A1(round_inst_aout_x[6]), .A2(reg_x_n503), .ZN(
        reg_x_n482) );
  NAND2_X1 reg_x_U133 ( .A1(reg_x_n480), .A2(reg_x_n479), .ZN(reg_x_n259) );
  NAND2_X1 reg_x_U132 ( .A1(state_x[6]), .A2(reg_x_n504), .ZN(reg_x_n479) );
  NAND2_X1 reg_x_U131 ( .A1(round_inst_aout_x[7]), .A2(reg_x_n503), .ZN(
        reg_x_n480) );
  NAND2_X1 reg_x_U130 ( .A1(reg_x_n478), .A2(reg_x_n477), .ZN(reg_x_n262) );
  NAND2_X1 reg_x_U129 ( .A1(state_x[3]), .A2(reg_x_n530), .ZN(reg_x_n477) );
  NAND2_X1 reg_x_U128 ( .A1(round_inst_aout_x[2]), .A2(reg_x_n529), .ZN(
        reg_x_n478) );
  NAND2_X1 reg_x_U127 ( .A1(reg_x_n476), .A2(reg_x_n475), .ZN(reg_x_n263) );
  NAND2_X1 reg_x_U126 ( .A1(state_x[2]), .A2(reg_x_n504), .ZN(reg_x_n475) );
  NAND2_X1 reg_x_U125 ( .A1(round_inst_aout_x[3]), .A2(reg_x_n503), .ZN(
        reg_x_n476) );
  NAND2_X1 reg_x_U124 ( .A1(reg_x_n474), .A2(reg_x_n473), .ZN(reg_x_n264) );
  NAND2_X1 reg_x_U123 ( .A1(state_x[1]), .A2(reg_x_n530), .ZN(reg_x_n473) );
  NAND2_X1 reg_x_U122 ( .A1(round_inst_aout_x[0]), .A2(reg_x_n529), .ZN(
        reg_x_n474) );
  NAND2_X1 reg_x_U121 ( .A1(reg_x_n472), .A2(reg_x_n471), .ZN(reg_x_n265) );
  NAND2_X1 reg_x_U120 ( .A1(state_x[0]), .A2(reg_x_n504), .ZN(reg_x_n471) );
  NAND2_X1 reg_x_U119 ( .A1(round_inst_srout_x[48]), .A2(reg_x_n503), .ZN(
        reg_x_n472) );
  NAND2_X1 reg_x_U118 ( .A1(reg_x_n470), .A2(reg_x_n469), .ZN(reg_x_n206) );
  NAND2_X1 reg_x_U117 ( .A1(state_x[59]), .A2(reg_x_n530), .ZN(reg_x_n469) );
  NAND2_X1 reg_x_U116 ( .A1(round_inst_aout_x[58]), .A2(reg_x_n529), .ZN(
        reg_x_n470) );
  NAND2_X1 reg_x_U115 ( .A1(reg_x_n468), .A2(reg_x_n467), .ZN(reg_x_n207) );
  NAND2_X1 reg_x_U114 ( .A1(state_x[58]), .A2(reg_x_n504), .ZN(reg_x_n467) );
  NAND2_X1 reg_x_U113 ( .A1(round_inst_aout_x[59]), .A2(reg_x_n503), .ZN(
        reg_x_n468) );
  NAND2_X1 reg_x_U112 ( .A1(reg_x_n466), .A2(reg_x_n465), .ZN(reg_x_n208) );
  NAND2_X1 reg_x_U111 ( .A1(state_x[57]), .A2(reg_x_n530), .ZN(reg_x_n465) );
  NAND2_X1 reg_x_U110 ( .A1(round_inst_aout_x[56]), .A2(reg_x_n529), .ZN(
        reg_x_n466) );
  NAND2_X1 reg_x_U109 ( .A1(reg_x_n464), .A2(reg_x_n463), .ZN(reg_x_n209) );
  NAND2_X1 reg_x_U108 ( .A1(state_x[56]), .A2(reg_x_n504), .ZN(reg_x_n463) );
  NAND2_X1 reg_x_U107 ( .A1(round_inst_srout_x[8]), .A2(reg_x_n503), .ZN(
        reg_x_n464) );
  INV_X1 reg_x_U106 ( .A(reg_x_n462), .ZN(reg_x_n503) );
  NAND2_X1 reg_x_U105 ( .A1(reg_x_n461), .A2(reg_x_n460), .ZN(reg_x_n210) );
  NAND2_X1 reg_x_U104 ( .A1(state_x[55]), .A2(reg_x_n530), .ZN(reg_x_n460) );
  NAND2_X1 reg_x_U103 ( .A1(round_inst_aout_x[54]), .A2(reg_x_n529), .ZN(
        reg_x_n461) );
  INV_X1 reg_x_U102 ( .A(reg_x_n462), .ZN(reg_x_n529) );
  NAND2_X1 reg_x_U101 ( .A1(reg_x_n459), .A2(reg_x_n458), .ZN(reg_x_n211) );
  NAND2_X1 reg_x_U100 ( .A1(state_x[54]), .A2(reg_x_n504), .ZN(reg_x_n458) );
  INV_X1 reg_x_U99 ( .A(reg_x_n457), .ZN(reg_x_n504) );
  NAND2_X1 reg_x_U98 ( .A1(round_inst_aout_x[55]), .A2(reg_x_n456), .ZN(
        reg_x_n459) );
  NAND2_X1 reg_x_U97 ( .A1(reg_x_n455), .A2(reg_x_n454), .ZN(reg_x_n212) );
  NAND2_X1 reg_x_U96 ( .A1(state_x[53]), .A2(reg_x_n530), .ZN(reg_x_n454) );
  INV_X1 reg_x_U95 ( .A(reg_x_n457), .ZN(reg_x_n530) );
  NAND2_X1 reg_x_U94 ( .A1(round_inst_aout_x[52]), .A2(reg_x_n456), .ZN(
        reg_x_n455) );
  NAND2_X1 reg_x_U93 ( .A1(reg_x_n453), .A2(reg_x_n452), .ZN(reg_x_n213) );
  NAND2_X1 reg_x_U92 ( .A1(state_x[52]), .A2(reg_x_n451), .ZN(reg_x_n452) );
  NAND2_X1 reg_x_U91 ( .A1(round_inst_srout_x[20]), .A2(reg_x_n456), .ZN(
        reg_x_n453) );
  NAND2_X1 reg_x_U90 ( .A1(reg_x_n450), .A2(reg_x_n449), .ZN(reg_x_n214) );
  NAND2_X1 reg_x_U89 ( .A1(state_x[51]), .A2(reg_x_n451), .ZN(reg_x_n449) );
  NAND2_X1 reg_x_U88 ( .A1(round_inst_aout_x[50]), .A2(reg_x_n456), .ZN(
        reg_x_n450) );
  NAND2_X1 reg_x_U87 ( .A1(reg_x_n448), .A2(reg_x_n447), .ZN(reg_x_n215) );
  NAND2_X1 reg_x_U86 ( .A1(state_x[50]), .A2(reg_x_n451), .ZN(reg_x_n447) );
  NAND2_X1 reg_x_U85 ( .A1(round_inst_aout_x[51]), .A2(reg_x_n456), .ZN(
        reg_x_n448) );
  NAND2_X1 reg_x_U84 ( .A1(reg_x_n446), .A2(reg_x_n445), .ZN(reg_x_n216) );
  NAND2_X1 reg_x_U83 ( .A1(state_x[49]), .A2(reg_x_n451), .ZN(reg_x_n445) );
  NAND2_X1 reg_x_U82 ( .A1(round_inst_aout_x[48]), .A2(reg_x_n456), .ZN(
        reg_x_n446) );
  NAND2_X1 reg_x_U81 ( .A1(reg_x_n444), .A2(reg_x_n443), .ZN(reg_x_n217) );
  NAND2_X1 reg_x_U80 ( .A1(state_x[48]), .A2(reg_x_n451), .ZN(reg_x_n443) );
  NAND2_X1 reg_x_U79 ( .A1(round_inst_srout_x[32]), .A2(reg_x_n456), .ZN(
        reg_x_n444) );
  NAND2_X1 reg_x_U78 ( .A1(reg_x_n442), .A2(reg_x_n441), .ZN(reg_x_n218) );
  NAND2_X1 reg_x_U77 ( .A1(state_x[47]), .A2(reg_x_n451), .ZN(reg_x_n441) );
  NAND2_X1 reg_x_U76 ( .A1(round_inst_aout_x[46]), .A2(reg_x_n440), .ZN(
        reg_x_n442) );
  NAND2_X1 reg_x_U75 ( .A1(reg_x_n439), .A2(reg_x_n438), .ZN(reg_x_n219) );
  NAND2_X1 reg_x_U74 ( .A1(state_x[46]), .A2(reg_x_n451), .ZN(reg_x_n438) );
  NAND2_X1 reg_x_U73 ( .A1(round_inst_aout_x[47]), .A2(reg_x_n440), .ZN(
        reg_x_n439) );
  NAND2_X1 reg_x_U72 ( .A1(reg_x_n437), .A2(reg_x_n436), .ZN(reg_x_n220) );
  NAND2_X1 reg_x_U71 ( .A1(state_x[45]), .A2(reg_x_n451), .ZN(reg_x_n436) );
  NAND2_X1 reg_x_U70 ( .A1(round_inst_aout_x[44]), .A2(reg_x_n440), .ZN(
        reg_x_n437) );
  NAND2_X1 reg_x_U69 ( .A1(reg_x_n435), .A2(reg_x_n434), .ZN(reg_x_n221) );
  NAND2_X1 reg_x_U68 ( .A1(state_x[44]), .A2(reg_x_n451), .ZN(reg_x_n434) );
  NAND2_X1 reg_x_U67 ( .A1(round_inst_srout_x[44]), .A2(reg_x_n440), .ZN(
        reg_x_n435) );
  NAND2_X1 reg_x_U66 ( .A1(reg_x_n433), .A2(reg_x_n432), .ZN(reg_x_n222) );
  NAND2_X1 reg_x_U65 ( .A1(state_x[43]), .A2(reg_x_n451), .ZN(reg_x_n432) );
  NAND2_X1 reg_x_U64 ( .A1(round_inst_aout_x[42]), .A2(reg_x_n440), .ZN(
        reg_x_n433) );
  NAND2_X1 reg_x_U63 ( .A1(reg_x_n431), .A2(reg_x_n430), .ZN(reg_x_n223) );
  NAND2_X1 reg_x_U62 ( .A1(state_x[42]), .A2(reg_x_n451), .ZN(reg_x_n430) );
  NAND2_X1 reg_x_U61 ( .A1(round_inst_aout_x[43]), .A2(reg_x_n440), .ZN(
        reg_x_n431) );
  NAND2_X1 reg_x_U60 ( .A1(reg_x_n429), .A2(reg_x_n428), .ZN(reg_x_n224) );
  NAND2_X1 reg_x_U59 ( .A1(state_x[41]), .A2(reg_x_n451), .ZN(reg_x_n428) );
  NAND2_X1 reg_x_U58 ( .A1(round_inst_aout_x[40]), .A2(reg_x_n440), .ZN(
        reg_x_n429) );
  NAND2_X1 reg_x_U57 ( .A1(reg_x_n427), .A2(reg_x_n426), .ZN(reg_x_n225) );
  NAND2_X1 reg_x_U56 ( .A1(state_x[40]), .A2(reg_x_n451), .ZN(reg_x_n426) );
  NAND2_X1 reg_x_U55 ( .A1(round_inst_srout_x[56]), .A2(reg_x_n440), .ZN(
        reg_x_n427) );
  NAND2_X1 reg_x_U54 ( .A1(reg_x_n425), .A2(reg_x_n424), .ZN(reg_x_n226) );
  NAND2_X1 reg_x_U53 ( .A1(state_x[39]), .A2(reg_x_n451), .ZN(reg_x_n424) );
  NAND2_X1 reg_x_U52 ( .A1(round_inst_aout_x[38]), .A2(reg_x_n440), .ZN(
        reg_x_n425) );
  NAND2_X1 reg_x_U51 ( .A1(reg_x_n423), .A2(reg_x_n422), .ZN(reg_x_n227) );
  NAND2_X1 reg_x_U50 ( .A1(state_x[38]), .A2(reg_x_n421), .ZN(reg_x_n422) );
  NAND2_X1 reg_x_U49 ( .A1(round_inst_aout_x[39]), .A2(reg_x_n440), .ZN(
        reg_x_n423) );
  NAND2_X1 reg_x_U48 ( .A1(reg_x_n420), .A2(reg_x_n419), .ZN(reg_x_n228) );
  NAND2_X1 reg_x_U47 ( .A1(state_x[37]), .A2(reg_x_n421), .ZN(reg_x_n419) );
  NAND2_X1 reg_x_U46 ( .A1(round_inst_aout_x[36]), .A2(reg_x_n440), .ZN(
        reg_x_n420) );
  NAND2_X1 reg_x_U45 ( .A1(reg_x_n418), .A2(reg_x_n417), .ZN(reg_x_n229) );
  NAND2_X1 reg_x_U44 ( .A1(state_x[36]), .A2(reg_x_n421), .ZN(reg_x_n417) );
  NAND2_X1 reg_x_U43 ( .A1(round_inst_srout_x[4]), .A2(reg_x_n440), .ZN(
        reg_x_n418) );
  NAND2_X1 reg_x_U42 ( .A1(reg_x_n416), .A2(reg_x_n415), .ZN(reg_x_n202) );
  NAND2_X1 reg_x_U41 ( .A1(state_x[63]), .A2(reg_x_n421), .ZN(reg_x_n415) );
  NAND2_X1 reg_x_U40 ( .A1(round_inst_aout_x[62]), .A2(reg_x_n440), .ZN(
        reg_x_n416) );
  NAND2_X1 reg_x_U39 ( .A1(reg_x_n414), .A2(reg_x_n413), .ZN(reg_x_n203) );
  NAND2_X1 reg_x_U38 ( .A1(state_x[62]), .A2(reg_x_n421), .ZN(reg_x_n413) );
  NAND2_X1 reg_x_U37 ( .A1(round_inst_aout_x[63]), .A2(reg_x_n440), .ZN(
        reg_x_n414) );
  NAND2_X1 reg_x_U36 ( .A1(reg_x_n412), .A2(reg_x_n411), .ZN(reg_x_n204) );
  NAND2_X1 reg_x_U35 ( .A1(state_x[61]), .A2(reg_x_n421), .ZN(reg_x_n411) );
  NAND2_X1 reg_x_U34 ( .A1(round_inst_aout_x[60]), .A2(reg_x_n440), .ZN(
        reg_x_n412) );
  NAND2_X1 reg_x_U33 ( .A1(reg_x_n410), .A2(reg_x_n409), .ZN(reg_x_n205) );
  NAND2_X1 reg_x_U32 ( .A1(state_x[60]), .A2(reg_x_n421), .ZN(reg_x_n409) );
  NAND2_X1 reg_x_U31 ( .A1(round_inst_srout_x[60]), .A2(reg_x_n440), .ZN(
        reg_x_n410) );
  NAND2_X1 reg_x_U30 ( .A1(reg_x_n408), .A2(reg_x_n407), .ZN(reg_x_n230) );
  NAND2_X1 reg_x_U29 ( .A1(state_x[35]), .A2(reg_x_n421), .ZN(reg_x_n407) );
  NAND2_X1 reg_x_U28 ( .A1(round_inst_aout_x[34]), .A2(reg_x_n440), .ZN(
        reg_x_n408) );
  NAND2_X1 reg_x_U27 ( .A1(reg_x_n406), .A2(reg_x_n405), .ZN(reg_x_n234) );
  NAND2_X1 reg_x_U26 ( .A1(state_x[31]), .A2(reg_x_n421), .ZN(reg_x_n405) );
  NAND2_X1 reg_x_U25 ( .A1(round_inst_aout_x[30]), .A2(reg_x_n440), .ZN(
        reg_x_n406) );
  NAND2_X1 reg_x_U24 ( .A1(reg_x_n404), .A2(reg_x_n403), .ZN(reg_x_n246) );
  NAND2_X1 reg_x_U23 ( .A1(state_x[19]), .A2(reg_x_n451), .ZN(reg_x_n403) );
  NAND2_X1 reg_x_U22 ( .A1(round_inst_aout_x[18]), .A2(reg_x_n440), .ZN(
        reg_x_n404) );
  NAND2_X1 reg_x_U21 ( .A1(reg_x_n402), .A2(reg_x_n401), .ZN(reg_x_n250) );
  NAND2_X1 reg_x_U20 ( .A1(state_x[15]), .A2(reg_x_n451), .ZN(reg_x_n401) );
  NAND2_X1 reg_x_U19 ( .A1(round_inst_aout_x[14]), .A2(reg_x_n456), .ZN(
        reg_x_n402) );
  NAND2_X1 reg_x_U18 ( .A1(reg_x_n400), .A2(reg_x_n399), .ZN(reg_x_n257) );
  NAND2_X1 reg_x_U17 ( .A1(state_x[8]), .A2(reg_x_n451), .ZN(reg_x_n399) );
  NAND2_X1 reg_x_U16 ( .A1(round_inst_srout_x[24]), .A2(reg_x_n440), .ZN(
        reg_x_n400) );
  NAND2_X1 reg_x_U15 ( .A1(reg_x_n398), .A2(reg_x_n397), .ZN(reg_x_n260) );
  NAND2_X1 reg_x_U14 ( .A1(state_x[5]), .A2(reg_x_n451), .ZN(reg_x_n397) );
  NAND2_X1 reg_x_U13 ( .A1(round_inst_aout_x[4]), .A2(reg_x_n456), .ZN(
        reg_x_n398) );
  NAND2_X1 reg_x_U12 ( .A1(reg_x_n396), .A2(reg_x_n395), .ZN(reg_x_n261) );
  NAND2_X1 reg_x_U11 ( .A1(reg_x_n440), .A2(round_inst_srout_x[36]), .ZN(
        reg_x_n395) );
  INV_X1 reg_x_U10 ( .A(reg_x_n462), .ZN(reg_x_n440) );
  INV_X1 reg_x_U9 ( .A(reg_x_n456), .ZN(reg_x_n462) );
  NAND2_X1 reg_x_U8 ( .A1(reg_x_n451), .A2(state_x[4]), .ZN(reg_x_n396) );
  INV_X1 reg_x_U7 ( .A(reg_x_n457), .ZN(reg_x_n451) );
  INV_X1 reg_x_U6 ( .A(reg_x_n421), .ZN(reg_x_n457) );
  INV_X1 reg_x_U5 ( .A(en_sig), .ZN(reg_x_n394) );
  NOR2_X1 reg_x_U4 ( .A1(rst), .A2(reg_x_n394), .ZN(reg_x_n421) );
  NOR2_X1 reg_x_U3 ( .A1(rst), .A2(en_sig), .ZN(reg_x_n456) );
  DFF_X1 reg_x_s_current_state_reg_0_ ( .D(reg_x_n265), .CK(clk), .Q(
        round_inst_srout_x[48]) );
  DFF_X1 reg_x_s_current_state_reg_1_ ( .D(reg_x_n264), .CK(clk), .Q(
        round_inst_aout_x[0]) );
  DFF_X1 reg_x_s_current_state_reg_2_ ( .D(reg_x_n263), .CK(clk), .Q(
        round_inst_aout_x[3]) );
  DFF_X1 reg_x_s_current_state_reg_3_ ( .D(reg_x_n262), .CK(clk), .Q(
        round_inst_aout_x[2]) );
  DFF_X1 reg_x_s_current_state_reg_4_ ( .D(reg_x_n261), .CK(clk), .Q(
        round_inst_srout_x[36]) );
  DFF_X1 reg_x_s_current_state_reg_5_ ( .D(reg_x_n260), .CK(clk), .Q(
        round_inst_aout_x[4]) );
  DFF_X1 reg_x_s_current_state_reg_6_ ( .D(reg_x_n259), .CK(clk), .Q(
        round_inst_aout_x[7]) );
  DFF_X1 reg_x_s_current_state_reg_7_ ( .D(reg_x_n258), .CK(clk), .Q(
        round_inst_aout_x[6]) );
  DFF_X1 reg_x_s_current_state_reg_8_ ( .D(reg_x_n257), .CK(clk), .Q(
        round_inst_srout_x[24]) );
  DFF_X1 reg_x_s_current_state_reg_9_ ( .D(reg_x_n256), .CK(clk), .Q(
        round_inst_aout_x[8]) );
  DFF_X1 reg_x_s_current_state_reg_10_ ( .D(reg_x_n255), .CK(clk), .Q(
        round_inst_aout_x[11]) );
  DFF_X1 reg_x_s_current_state_reg_11_ ( .D(reg_x_n254), .CK(clk), .Q(
        round_inst_aout_x[10]) );
  DFF_X1 reg_x_s_current_state_reg_12_ ( .D(reg_x_n253), .CK(clk), .Q(
        round_inst_srout_x[12]) );
  DFF_X1 reg_x_s_current_state_reg_13_ ( .D(reg_x_n252), .CK(clk), .Q(
        round_inst_aout_x[12]) );
  DFF_X1 reg_x_s_current_state_reg_14_ ( .D(reg_x_n251), .CK(clk), .Q(
        round_inst_aout_x[15]) );
  DFF_X1 reg_x_s_current_state_reg_15_ ( .D(reg_x_n250), .CK(clk), .Q(
        round_inst_aout_x[14]) );
  DFF_X1 reg_x_s_current_state_reg_16_ ( .D(reg_x_n249), .CK(clk), .Q(
        round_inst_srout_x[0]) );
  DFF_X1 reg_x_s_current_state_reg_17_ ( .D(reg_x_n248), .CK(clk), .Q(
        round_inst_aout_x[16]) );
  DFF_X1 reg_x_s_current_state_reg_18_ ( .D(reg_x_n247), .CK(clk), .Q(
        round_inst_aout_x[19]) );
  DFF_X1 reg_x_s_current_state_reg_19_ ( .D(reg_x_n246), .CK(clk), .Q(
        round_inst_aout_x[18]) );
  DFF_X1 reg_x_s_current_state_reg_20_ ( .D(reg_x_n245), .CK(clk), .Q(
        round_inst_srout_x[52]) );
  DFF_X1 reg_x_s_current_state_reg_21_ ( .D(reg_x_n244), .CK(clk), .Q(
        round_inst_aout_x[20]) );
  DFF_X1 reg_x_s_current_state_reg_22_ ( .D(reg_x_n243), .CK(clk), .Q(
        round_inst_aout_x[23]) );
  DFF_X1 reg_x_s_current_state_reg_23_ ( .D(reg_x_n242), .CK(clk), .Q(
        round_inst_aout_x[22]) );
  DFF_X1 reg_x_s_current_state_reg_24_ ( .D(reg_x_n241), .CK(clk), .Q(
        round_inst_srout_x[40]) );
  DFF_X1 reg_x_s_current_state_reg_25_ ( .D(reg_x_n240), .CK(clk), .Q(
        round_inst_aout_x[24]) );
  DFF_X1 reg_x_s_current_state_reg_26_ ( .D(reg_x_n239), .CK(clk), .Q(
        round_inst_aout_x[27]) );
  DFF_X1 reg_x_s_current_state_reg_27_ ( .D(reg_x_n238), .CK(clk), .Q(
        round_inst_aout_x[26]) );
  DFF_X1 reg_x_s_current_state_reg_28_ ( .D(reg_x_n237), .CK(clk), .Q(
        round_inst_srout_x[28]) );
  DFF_X1 reg_x_s_current_state_reg_29_ ( .D(reg_x_n236), .CK(clk), .Q(
        round_inst_aout_x[28]) );
  DFF_X1 reg_x_s_current_state_reg_30_ ( .D(reg_x_n235), .CK(clk), .Q(
        round_inst_aout_x[31]) );
  DFF_X1 reg_x_s_current_state_reg_31_ ( .D(reg_x_n234), .CK(clk), .Q(
        round_inst_aout_x[30]) );
  DFF_X1 reg_x_s_current_state_reg_32_ ( .D(reg_x_n233), .CK(clk), .Q(
        round_inst_srout_x[16]) );
  DFF_X1 reg_x_s_current_state_reg_33_ ( .D(reg_x_n232), .CK(clk), .Q(
        round_inst_aout_x[32]) );
  DFF_X1 reg_x_s_current_state_reg_34_ ( .D(reg_x_n231), .CK(clk), .Q(
        round_inst_aout_x[35]) );
  DFF_X1 reg_x_s_current_state_reg_35_ ( .D(reg_x_n230), .CK(clk), .Q(
        round_inst_aout_x[34]) );
  DFF_X1 reg_x_s_current_state_reg_36_ ( .D(reg_x_n229), .CK(clk), .Q(
        round_inst_srout_x[4]) );
  DFF_X1 reg_x_s_current_state_reg_37_ ( .D(reg_x_n228), .CK(clk), .Q(
        round_inst_aout_x[36]) );
  DFF_X1 reg_x_s_current_state_reg_38_ ( .D(reg_x_n227), .CK(clk), .Q(
        round_inst_aout_x[39]) );
  DFF_X1 reg_x_s_current_state_reg_39_ ( .D(reg_x_n226), .CK(clk), .Q(
        round_inst_aout_x[38]) );
  DFF_X1 reg_x_s_current_state_reg_40_ ( .D(reg_x_n225), .CK(clk), .Q(
        round_inst_srout_x[56]) );
  DFF_X1 reg_x_s_current_state_reg_41_ ( .D(reg_x_n224), .CK(clk), .Q(
        round_inst_aout_x[40]) );
  DFF_X1 reg_x_s_current_state_reg_42_ ( .D(reg_x_n223), .CK(clk), .Q(
        round_inst_aout_x[43]) );
  DFF_X1 reg_x_s_current_state_reg_43_ ( .D(reg_x_n222), .CK(clk), .Q(
        round_inst_aout_x[42]) );
  DFF_X1 reg_x_s_current_state_reg_44_ ( .D(reg_x_n221), .CK(clk), .Q(
        round_inst_srout_x[44]) );
  DFF_X1 reg_x_s_current_state_reg_45_ ( .D(reg_x_n220), .CK(clk), .Q(
        round_inst_aout_x[44]) );
  DFF_X1 reg_x_s_current_state_reg_46_ ( .D(reg_x_n219), .CK(clk), .Q(
        round_inst_aout_x[47]) );
  DFF_X1 reg_x_s_current_state_reg_47_ ( .D(reg_x_n218), .CK(clk), .Q(
        round_inst_aout_x[46]) );
  DFF_X1 reg_x_s_current_state_reg_48_ ( .D(reg_x_n217), .CK(clk), .Q(
        round_inst_srout_x[32]) );
  DFF_X1 reg_x_s_current_state_reg_49_ ( .D(reg_x_n216), .CK(clk), .Q(
        round_inst_aout_x[48]) );
  DFF_X1 reg_x_s_current_state_reg_50_ ( .D(reg_x_n215), .CK(clk), .Q(
        round_inst_aout_x[51]) );
  DFF_X1 reg_x_s_current_state_reg_51_ ( .D(reg_x_n214), .CK(clk), .Q(
        round_inst_aout_x[50]) );
  DFF_X1 reg_x_s_current_state_reg_52_ ( .D(reg_x_n213), .CK(clk), .Q(
        round_inst_srout_x[20]) );
  DFF_X1 reg_x_s_current_state_reg_53_ ( .D(reg_x_n212), .CK(clk), .Q(
        round_inst_aout_x[52]) );
  DFF_X1 reg_x_s_current_state_reg_54_ ( .D(reg_x_n211), .CK(clk), .Q(
        round_inst_aout_x[55]) );
  DFF_X1 reg_x_s_current_state_reg_55_ ( .D(reg_x_n210), .CK(clk), .Q(
        round_inst_aout_x[54]) );
  DFF_X1 reg_x_s_current_state_reg_56_ ( .D(reg_x_n209), .CK(clk), .Q(
        round_inst_srout_x[8]) );
  DFF_X1 reg_x_s_current_state_reg_57_ ( .D(reg_x_n208), .CK(clk), .Q(
        round_inst_aout_x[56]) );
  DFF_X1 reg_x_s_current_state_reg_58_ ( .D(reg_x_n207), .CK(clk), .Q(
        round_inst_aout_x[59]) );
  DFF_X1 reg_x_s_current_state_reg_59_ ( .D(reg_x_n206), .CK(clk), .Q(
        round_inst_aout_x[58]) );
  DFF_X1 reg_x_s_current_state_reg_60_ ( .D(reg_x_n205), .CK(clk), .Q(
        round_inst_srout_x[60]) );
  DFF_X1 reg_x_s_current_state_reg_61_ ( .D(reg_x_n204), .CK(clk), .Q(
        round_inst_aout_x[60]) );
  DFF_X1 reg_x_s_current_state_reg_62_ ( .D(reg_x_n203), .CK(clk), .Q(
        round_inst_aout_x[63]) );
  DFF_X1 reg_x_s_current_state_reg_63_ ( .D(reg_x_n202), .CK(clk), .Q(
        round_inst_aout_x[62]) );
  NAND2_X1 reg_y_U205 ( .A1(reg_y_n532), .A2(reg_y_n531), .ZN(reg_y_n230) );
  NAND2_X1 reg_y_U204 ( .A1(state_y[35]), .A2(reg_y_n530), .ZN(reg_y_n531) );
  NAND2_X1 reg_y_U203 ( .A1(round_inst_aout_y[34]), .A2(reg_y_n529), .ZN(
        reg_y_n532) );
  NAND2_X1 reg_y_U202 ( .A1(reg_y_n528), .A2(reg_y_n527), .ZN(reg_y_n231) );
  NAND2_X1 reg_y_U201 ( .A1(state_y[34]), .A2(reg_y_n530), .ZN(reg_y_n527) );
  NAND2_X1 reg_y_U200 ( .A1(round_inst_aout_y[35]), .A2(reg_y_n529), .ZN(
        reg_y_n528) );
  NAND2_X1 reg_y_U199 ( .A1(reg_y_n526), .A2(reg_y_n525), .ZN(reg_y_n232) );
  NAND2_X1 reg_y_U198 ( .A1(state_y[33]), .A2(reg_y_n530), .ZN(reg_y_n525) );
  NAND2_X1 reg_y_U197 ( .A1(round_inst_aout_y[32]), .A2(reg_y_n529), .ZN(
        reg_y_n526) );
  NAND2_X1 reg_y_U196 ( .A1(reg_y_n524), .A2(reg_y_n523), .ZN(reg_y_n233) );
  NAND2_X1 reg_y_U195 ( .A1(state_y[32]), .A2(reg_y_n530), .ZN(reg_y_n523) );
  NAND2_X1 reg_y_U194 ( .A1(round_inst_srout_y[16]), .A2(reg_y_n529), .ZN(
        reg_y_n524) );
  NAND2_X1 reg_y_U193 ( .A1(reg_y_n522), .A2(reg_y_n521), .ZN(reg_y_n234) );
  NAND2_X1 reg_y_U192 ( .A1(state_y[31]), .A2(reg_y_n530), .ZN(reg_y_n521) );
  NAND2_X1 reg_y_U191 ( .A1(round_inst_aout_y[30]), .A2(reg_y_n529), .ZN(
        reg_y_n522) );
  NAND2_X1 reg_y_U190 ( .A1(reg_y_n520), .A2(reg_y_n519), .ZN(reg_y_n235) );
  NAND2_X1 reg_y_U189 ( .A1(state_y[30]), .A2(reg_y_n530), .ZN(reg_y_n519) );
  NAND2_X1 reg_y_U188 ( .A1(round_inst_aout_y[31]), .A2(reg_y_n529), .ZN(
        reg_y_n520) );
  NAND2_X1 reg_y_U187 ( .A1(reg_y_n518), .A2(reg_y_n517), .ZN(reg_y_n237) );
  NAND2_X1 reg_y_U186 ( .A1(state_y[28]), .A2(reg_y_n530), .ZN(reg_y_n517) );
  NAND2_X1 reg_y_U185 ( .A1(round_inst_srout_y[28]), .A2(reg_y_n529), .ZN(
        reg_y_n518) );
  NAND2_X1 reg_y_U184 ( .A1(reg_y_n516), .A2(reg_y_n515), .ZN(reg_y_n238) );
  NAND2_X1 reg_y_U183 ( .A1(state_y[27]), .A2(reg_y_n530), .ZN(reg_y_n515) );
  NAND2_X1 reg_y_U182 ( .A1(round_inst_aout_y[26]), .A2(reg_y_n529), .ZN(
        reg_y_n516) );
  NAND2_X1 reg_y_U181 ( .A1(reg_y_n514), .A2(reg_y_n513), .ZN(reg_y_n239) );
  NAND2_X1 reg_y_U180 ( .A1(state_y[26]), .A2(reg_y_n530), .ZN(reg_y_n513) );
  NAND2_X1 reg_y_U179 ( .A1(round_inst_aout_y[27]), .A2(reg_y_n529), .ZN(
        reg_y_n514) );
  NAND2_X1 reg_y_U178 ( .A1(reg_y_n512), .A2(reg_y_n511), .ZN(reg_y_n241) );
  NAND2_X1 reg_y_U177 ( .A1(state_y[24]), .A2(reg_y_n530), .ZN(reg_y_n511) );
  NAND2_X1 reg_y_U176 ( .A1(round_inst_srout_y[40]), .A2(reg_y_n529), .ZN(
        reg_y_n512) );
  NAND2_X1 reg_y_U175 ( .A1(reg_y_n510), .A2(reg_y_n509), .ZN(reg_y_n242) );
  NAND2_X1 reg_y_U174 ( .A1(state_y[23]), .A2(reg_y_n530), .ZN(reg_y_n509) );
  NAND2_X1 reg_y_U173 ( .A1(round_inst_aout_y[22]), .A2(reg_y_n529), .ZN(
        reg_y_n510) );
  NAND2_X1 reg_y_U172 ( .A1(reg_y_n508), .A2(reg_y_n507), .ZN(reg_y_n243) );
  NAND2_X1 reg_y_U171 ( .A1(state_y[22]), .A2(reg_y_n530), .ZN(reg_y_n507) );
  NAND2_X1 reg_y_U170 ( .A1(round_inst_aout_y[23]), .A2(reg_y_n529), .ZN(
        reg_y_n508) );
  NAND2_X1 reg_y_U169 ( .A1(reg_y_n506), .A2(reg_y_n505), .ZN(reg_y_n244) );
  NAND2_X1 reg_y_U168 ( .A1(state_y[21]), .A2(reg_y_n504), .ZN(reg_y_n505) );
  NAND2_X1 reg_y_U167 ( .A1(round_inst_aout_y[20]), .A2(reg_y_n503), .ZN(
        reg_y_n506) );
  NAND2_X1 reg_y_U166 ( .A1(reg_y_n502), .A2(reg_y_n501), .ZN(reg_y_n245) );
  NAND2_X1 reg_y_U165 ( .A1(state_y[20]), .A2(reg_y_n504), .ZN(reg_y_n501) );
  NAND2_X1 reg_y_U164 ( .A1(round_inst_srout_y[52]), .A2(reg_y_n503), .ZN(
        reg_y_n502) );
  NAND2_X1 reg_y_U163 ( .A1(reg_y_n500), .A2(reg_y_n499), .ZN(reg_y_n246) );
  NAND2_X1 reg_y_U162 ( .A1(state_y[19]), .A2(reg_y_n504), .ZN(reg_y_n499) );
  NAND2_X1 reg_y_U161 ( .A1(round_inst_aout_y[18]), .A2(reg_y_n503), .ZN(
        reg_y_n500) );
  NAND2_X1 reg_y_U160 ( .A1(reg_y_n498), .A2(reg_y_n497), .ZN(reg_y_n247) );
  NAND2_X1 reg_y_U159 ( .A1(state_y[18]), .A2(reg_y_n504), .ZN(reg_y_n497) );
  NAND2_X1 reg_y_U158 ( .A1(round_inst_aout_y[19]), .A2(reg_y_n503), .ZN(
        reg_y_n498) );
  NAND2_X1 reg_y_U157 ( .A1(reg_y_n496), .A2(reg_y_n495), .ZN(reg_y_n248) );
  NAND2_X1 reg_y_U156 ( .A1(state_y[17]), .A2(reg_y_n504), .ZN(reg_y_n495) );
  NAND2_X1 reg_y_U155 ( .A1(round_inst_aout_y[16]), .A2(reg_y_n503), .ZN(
        reg_y_n496) );
  NAND2_X1 reg_y_U154 ( .A1(reg_y_n494), .A2(reg_y_n493), .ZN(reg_y_n249) );
  NAND2_X1 reg_y_U153 ( .A1(state_y[16]), .A2(reg_y_n504), .ZN(reg_y_n493) );
  NAND2_X1 reg_y_U152 ( .A1(round_inst_srout_y[0]), .A2(reg_y_n503), .ZN(
        reg_y_n494) );
  NAND2_X1 reg_y_U151 ( .A1(reg_y_n492), .A2(reg_y_n491), .ZN(reg_y_n251) );
  NAND2_X1 reg_y_U150 ( .A1(state_y[14]), .A2(reg_y_n504), .ZN(reg_y_n491) );
  NAND2_X1 reg_y_U149 ( .A1(round_inst_aout_y[15]), .A2(reg_y_n503), .ZN(
        reg_y_n492) );
  NAND2_X1 reg_y_U148 ( .A1(reg_y_n490), .A2(reg_y_n489), .ZN(reg_y_n252) );
  NAND2_X1 reg_y_U147 ( .A1(state_y[13]), .A2(reg_y_n504), .ZN(reg_y_n489) );
  NAND2_X1 reg_y_U146 ( .A1(round_inst_aout_y[12]), .A2(reg_y_n503), .ZN(
        reg_y_n490) );
  NAND2_X1 reg_y_U145 ( .A1(reg_y_n488), .A2(reg_y_n487), .ZN(reg_y_n253) );
  NAND2_X1 reg_y_U144 ( .A1(state_y[12]), .A2(reg_y_n504), .ZN(reg_y_n487) );
  NAND2_X1 reg_y_U143 ( .A1(round_inst_srout_y[12]), .A2(reg_y_n503), .ZN(
        reg_y_n488) );
  NAND2_X1 reg_y_U142 ( .A1(reg_y_n486), .A2(reg_y_n485), .ZN(reg_y_n255) );
  NAND2_X1 reg_y_U141 ( .A1(state_y[10]), .A2(reg_y_n504), .ZN(reg_y_n485) );
  NAND2_X1 reg_y_U140 ( .A1(round_inst_aout_y[11]), .A2(reg_y_n503), .ZN(
        reg_y_n486) );
  NAND2_X1 reg_y_U139 ( .A1(reg_y_n484), .A2(reg_y_n483), .ZN(reg_y_n256) );
  NAND2_X1 reg_y_U138 ( .A1(state_y[9]), .A2(reg_y_n504), .ZN(reg_y_n483) );
  NAND2_X1 reg_y_U137 ( .A1(round_inst_aout_y[8]), .A2(reg_y_n503), .ZN(
        reg_y_n484) );
  NAND2_X1 reg_y_U136 ( .A1(reg_y_n482), .A2(reg_y_n481), .ZN(reg_y_n257) );
  NAND2_X1 reg_y_U135 ( .A1(state_y[8]), .A2(reg_y_n504), .ZN(reg_y_n481) );
  NAND2_X1 reg_y_U134 ( .A1(round_inst_srout_y[24]), .A2(reg_y_n503), .ZN(
        reg_y_n482) );
  NAND2_X1 reg_y_U133 ( .A1(reg_y_n480), .A2(reg_y_n479), .ZN(reg_y_n260) );
  NAND2_X1 reg_y_U132 ( .A1(state_y[5]), .A2(reg_y_n504), .ZN(reg_y_n479) );
  NAND2_X1 reg_y_U131 ( .A1(round_inst_aout_y[4]), .A2(reg_y_n503), .ZN(
        reg_y_n480) );
  NAND2_X1 reg_y_U130 ( .A1(reg_y_n478), .A2(reg_y_n477), .ZN(reg_y_n261) );
  NAND2_X1 reg_y_U129 ( .A1(state_y[4]), .A2(reg_y_n530), .ZN(reg_y_n477) );
  NAND2_X1 reg_y_U128 ( .A1(round_inst_srout_y[36]), .A2(reg_y_n529), .ZN(
        reg_y_n478) );
  NAND2_X1 reg_y_U127 ( .A1(reg_y_n476), .A2(reg_y_n475), .ZN(reg_y_n262) );
  NAND2_X1 reg_y_U126 ( .A1(state_y[3]), .A2(reg_y_n504), .ZN(reg_y_n475) );
  NAND2_X1 reg_y_U125 ( .A1(round_inst_aout_y[2]), .A2(reg_y_n503), .ZN(
        reg_y_n476) );
  NAND2_X1 reg_y_U124 ( .A1(reg_y_n474), .A2(reg_y_n473), .ZN(reg_y_n263) );
  NAND2_X1 reg_y_U123 ( .A1(state_y[2]), .A2(reg_y_n530), .ZN(reg_y_n473) );
  NAND2_X1 reg_y_U122 ( .A1(round_inst_aout_y[3]), .A2(reg_y_n529), .ZN(
        reg_y_n474) );
  NAND2_X1 reg_y_U121 ( .A1(reg_y_n472), .A2(reg_y_n471), .ZN(reg_y_n264) );
  NAND2_X1 reg_y_U120 ( .A1(state_y[1]), .A2(reg_y_n504), .ZN(reg_y_n471) );
  NAND2_X1 reg_y_U119 ( .A1(round_inst_aout_y[0]), .A2(reg_y_n503), .ZN(
        reg_y_n472) );
  NAND2_X1 reg_y_U118 ( .A1(reg_y_n470), .A2(reg_y_n469), .ZN(reg_y_n265) );
  NAND2_X1 reg_y_U117 ( .A1(state_y[0]), .A2(reg_y_n530), .ZN(reg_y_n469) );
  NAND2_X1 reg_y_U116 ( .A1(round_inst_srout_y[48]), .A2(reg_y_n529), .ZN(
        reg_y_n470) );
  NAND2_X1 reg_y_U115 ( .A1(reg_y_n468), .A2(reg_y_n467), .ZN(reg_y_n206) );
  NAND2_X1 reg_y_U114 ( .A1(state_y[59]), .A2(reg_y_n504), .ZN(reg_y_n467) );
  NAND2_X1 reg_y_U113 ( .A1(round_inst_aout_y[58]), .A2(reg_y_n503), .ZN(
        reg_y_n468) );
  NAND2_X1 reg_y_U112 ( .A1(reg_y_n466), .A2(reg_y_n465), .ZN(reg_y_n207) );
  NAND2_X1 reg_y_U111 ( .A1(state_y[58]), .A2(reg_y_n530), .ZN(reg_y_n465) );
  NAND2_X1 reg_y_U110 ( .A1(round_inst_aout_y[59]), .A2(reg_y_n529), .ZN(
        reg_y_n466) );
  NAND2_X1 reg_y_U109 ( .A1(reg_y_n464), .A2(reg_y_n463), .ZN(reg_y_n208) );
  NAND2_X1 reg_y_U108 ( .A1(state_y[57]), .A2(reg_y_n504), .ZN(reg_y_n463) );
  NAND2_X1 reg_y_U107 ( .A1(round_inst_aout_y[56]), .A2(reg_y_n503), .ZN(
        reg_y_n464) );
  INV_X1 reg_y_U106 ( .A(reg_y_n462), .ZN(reg_y_n503) );
  NAND2_X1 reg_y_U105 ( .A1(reg_y_n461), .A2(reg_y_n460), .ZN(reg_y_n209) );
  NAND2_X1 reg_y_U104 ( .A1(state_y[56]), .A2(reg_y_n530), .ZN(reg_y_n460) );
  NAND2_X1 reg_y_U103 ( .A1(round_inst_srout_y[8]), .A2(reg_y_n529), .ZN(
        reg_y_n461) );
  INV_X1 reg_y_U102 ( .A(reg_y_n462), .ZN(reg_y_n529) );
  NAND2_X1 reg_y_U101 ( .A1(reg_y_n459), .A2(reg_y_n458), .ZN(reg_y_n210) );
  NAND2_X1 reg_y_U100 ( .A1(state_y[55]), .A2(reg_y_n504), .ZN(reg_y_n458) );
  INV_X1 reg_y_U99 ( .A(reg_y_n457), .ZN(reg_y_n504) );
  NAND2_X1 reg_y_U98 ( .A1(round_inst_aout_y[54]), .A2(reg_y_n456), .ZN(
        reg_y_n459) );
  NAND2_X1 reg_y_U97 ( .A1(reg_y_n455), .A2(reg_y_n454), .ZN(reg_y_n211) );
  NAND2_X1 reg_y_U96 ( .A1(state_y[54]), .A2(reg_y_n530), .ZN(reg_y_n454) );
  INV_X1 reg_y_U95 ( .A(reg_y_n457), .ZN(reg_y_n530) );
  NAND2_X1 reg_y_U94 ( .A1(round_inst_aout_y[55]), .A2(reg_y_n456), .ZN(
        reg_y_n455) );
  NAND2_X1 reg_y_U93 ( .A1(reg_y_n453), .A2(reg_y_n452), .ZN(reg_y_n212) );
  NAND2_X1 reg_y_U92 ( .A1(state_y[53]), .A2(reg_y_n451), .ZN(reg_y_n452) );
  NAND2_X1 reg_y_U91 ( .A1(round_inst_aout_y[52]), .A2(reg_y_n456), .ZN(
        reg_y_n453) );
  NAND2_X1 reg_y_U90 ( .A1(reg_y_n450), .A2(reg_y_n449), .ZN(reg_y_n213) );
  NAND2_X1 reg_y_U89 ( .A1(state_y[52]), .A2(reg_y_n451), .ZN(reg_y_n449) );
  NAND2_X1 reg_y_U88 ( .A1(round_inst_srout_y[20]), .A2(reg_y_n456), .ZN(
        reg_y_n450) );
  NAND2_X1 reg_y_U87 ( .A1(reg_y_n448), .A2(reg_y_n447), .ZN(reg_y_n214) );
  NAND2_X1 reg_y_U86 ( .A1(state_y[51]), .A2(reg_y_n451), .ZN(reg_y_n447) );
  NAND2_X1 reg_y_U85 ( .A1(round_inst_aout_y[50]), .A2(reg_y_n456), .ZN(
        reg_y_n448) );
  NAND2_X1 reg_y_U84 ( .A1(reg_y_n446), .A2(reg_y_n445), .ZN(reg_y_n215) );
  NAND2_X1 reg_y_U83 ( .A1(state_y[50]), .A2(reg_y_n451), .ZN(reg_y_n445) );
  NAND2_X1 reg_y_U82 ( .A1(round_inst_aout_y[51]), .A2(reg_y_n456), .ZN(
        reg_y_n446) );
  NAND2_X1 reg_y_U81 ( .A1(reg_y_n444), .A2(reg_y_n443), .ZN(reg_y_n216) );
  NAND2_X1 reg_y_U80 ( .A1(state_y[49]), .A2(reg_y_n451), .ZN(reg_y_n443) );
  NAND2_X1 reg_y_U79 ( .A1(round_inst_aout_y[48]), .A2(reg_y_n456), .ZN(
        reg_y_n444) );
  NAND2_X1 reg_y_U78 ( .A1(reg_y_n442), .A2(reg_y_n441), .ZN(reg_y_n217) );
  NAND2_X1 reg_y_U77 ( .A1(state_y[48]), .A2(reg_y_n451), .ZN(reg_y_n441) );
  NAND2_X1 reg_y_U76 ( .A1(round_inst_srout_y[32]), .A2(reg_y_n440), .ZN(
        reg_y_n442) );
  NAND2_X1 reg_y_U75 ( .A1(reg_y_n439), .A2(reg_y_n438), .ZN(reg_y_n218) );
  NAND2_X1 reg_y_U74 ( .A1(state_y[47]), .A2(reg_y_n451), .ZN(reg_y_n438) );
  NAND2_X1 reg_y_U73 ( .A1(round_inst_aout_y[46]), .A2(reg_y_n440), .ZN(
        reg_y_n439) );
  NAND2_X1 reg_y_U72 ( .A1(reg_y_n437), .A2(reg_y_n436), .ZN(reg_y_n219) );
  NAND2_X1 reg_y_U71 ( .A1(state_y[46]), .A2(reg_y_n451), .ZN(reg_y_n436) );
  NAND2_X1 reg_y_U70 ( .A1(round_inst_aout_y[47]), .A2(reg_y_n440), .ZN(
        reg_y_n437) );
  NAND2_X1 reg_y_U69 ( .A1(reg_y_n435), .A2(reg_y_n434), .ZN(reg_y_n220) );
  NAND2_X1 reg_y_U68 ( .A1(state_y[45]), .A2(reg_y_n451), .ZN(reg_y_n434) );
  NAND2_X1 reg_y_U67 ( .A1(round_inst_aout_y[44]), .A2(reg_y_n440), .ZN(
        reg_y_n435) );
  NAND2_X1 reg_y_U66 ( .A1(reg_y_n433), .A2(reg_y_n432), .ZN(reg_y_n221) );
  NAND2_X1 reg_y_U65 ( .A1(state_y[44]), .A2(reg_y_n451), .ZN(reg_y_n432) );
  NAND2_X1 reg_y_U64 ( .A1(round_inst_srout_y[44]), .A2(reg_y_n440), .ZN(
        reg_y_n433) );
  NAND2_X1 reg_y_U63 ( .A1(reg_y_n431), .A2(reg_y_n430), .ZN(reg_y_n222) );
  NAND2_X1 reg_y_U62 ( .A1(state_y[43]), .A2(reg_y_n451), .ZN(reg_y_n430) );
  NAND2_X1 reg_y_U61 ( .A1(round_inst_aout_y[42]), .A2(reg_y_n440), .ZN(
        reg_y_n431) );
  NAND2_X1 reg_y_U60 ( .A1(reg_y_n429), .A2(reg_y_n428), .ZN(reg_y_n223) );
  NAND2_X1 reg_y_U59 ( .A1(state_y[42]), .A2(reg_y_n451), .ZN(reg_y_n428) );
  NAND2_X1 reg_y_U58 ( .A1(round_inst_aout_y[43]), .A2(reg_y_n440), .ZN(
        reg_y_n429) );
  NAND2_X1 reg_y_U57 ( .A1(reg_y_n427), .A2(reg_y_n426), .ZN(reg_y_n224) );
  NAND2_X1 reg_y_U56 ( .A1(state_y[41]), .A2(reg_y_n451), .ZN(reg_y_n426) );
  NAND2_X1 reg_y_U55 ( .A1(round_inst_aout_y[40]), .A2(reg_y_n440), .ZN(
        reg_y_n427) );
  NAND2_X1 reg_y_U54 ( .A1(reg_y_n425), .A2(reg_y_n424), .ZN(reg_y_n225) );
  NAND2_X1 reg_y_U53 ( .A1(state_y[40]), .A2(reg_y_n451), .ZN(reg_y_n424) );
  NAND2_X1 reg_y_U52 ( .A1(round_inst_srout_y[56]), .A2(reg_y_n440), .ZN(
        reg_y_n425) );
  NAND2_X1 reg_y_U51 ( .A1(reg_y_n423), .A2(reg_y_n422), .ZN(reg_y_n226) );
  NAND2_X1 reg_y_U50 ( .A1(state_y[39]), .A2(reg_y_n421), .ZN(reg_y_n422) );
  NAND2_X1 reg_y_U49 ( .A1(round_inst_aout_y[38]), .A2(reg_y_n440), .ZN(
        reg_y_n423) );
  NAND2_X1 reg_y_U48 ( .A1(reg_y_n420), .A2(reg_y_n419), .ZN(reg_y_n227) );
  NAND2_X1 reg_y_U47 ( .A1(state_y[38]), .A2(reg_y_n421), .ZN(reg_y_n419) );
  NAND2_X1 reg_y_U46 ( .A1(round_inst_aout_y[39]), .A2(reg_y_n440), .ZN(
        reg_y_n420) );
  NAND2_X1 reg_y_U45 ( .A1(reg_y_n418), .A2(reg_y_n417), .ZN(reg_y_n228) );
  NAND2_X1 reg_y_U44 ( .A1(state_y[37]), .A2(reg_y_n421), .ZN(reg_y_n417) );
  NAND2_X1 reg_y_U43 ( .A1(round_inst_aout_y[36]), .A2(reg_y_n440), .ZN(
        reg_y_n418) );
  NAND2_X1 reg_y_U42 ( .A1(reg_y_n416), .A2(reg_y_n415), .ZN(reg_y_n229) );
  NAND2_X1 reg_y_U41 ( .A1(state_y[36]), .A2(reg_y_n421), .ZN(reg_y_n415) );
  NAND2_X1 reg_y_U40 ( .A1(round_inst_srout_y[4]), .A2(reg_y_n440), .ZN(
        reg_y_n416) );
  NAND2_X1 reg_y_U39 ( .A1(reg_y_n414), .A2(reg_y_n413), .ZN(reg_y_n202) );
  NAND2_X1 reg_y_U38 ( .A1(state_y[63]), .A2(reg_y_n421), .ZN(reg_y_n413) );
  NAND2_X1 reg_y_U37 ( .A1(round_inst_aout_y[62]), .A2(reg_y_n440), .ZN(
        reg_y_n414) );
  NAND2_X1 reg_y_U36 ( .A1(reg_y_n412), .A2(reg_y_n411), .ZN(reg_y_n203) );
  NAND2_X1 reg_y_U35 ( .A1(state_y[62]), .A2(reg_y_n421), .ZN(reg_y_n411) );
  NAND2_X1 reg_y_U34 ( .A1(round_inst_aout_y[63]), .A2(reg_y_n440), .ZN(
        reg_y_n412) );
  NAND2_X1 reg_y_U33 ( .A1(reg_y_n410), .A2(reg_y_n409), .ZN(reg_y_n204) );
  NAND2_X1 reg_y_U32 ( .A1(state_y[61]), .A2(reg_y_n421), .ZN(reg_y_n409) );
  NAND2_X1 reg_y_U31 ( .A1(round_inst_aout_y[60]), .A2(reg_y_n440), .ZN(
        reg_y_n410) );
  NAND2_X1 reg_y_U30 ( .A1(reg_y_n408), .A2(reg_y_n407), .ZN(reg_y_n205) );
  NAND2_X1 reg_y_U29 ( .A1(state_y[60]), .A2(reg_y_n421), .ZN(reg_y_n407) );
  NAND2_X1 reg_y_U28 ( .A1(round_inst_srout_y[60]), .A2(reg_y_n440), .ZN(
        reg_y_n408) );
  NAND2_X1 reg_y_U27 ( .A1(reg_y_n406), .A2(reg_y_n405), .ZN(reg_y_n236) );
  NAND2_X1 reg_y_U26 ( .A1(state_y[29]), .A2(reg_y_n421), .ZN(reg_y_n405) );
  NAND2_X1 reg_y_U25 ( .A1(round_inst_aout_y[28]), .A2(reg_y_n440), .ZN(
        reg_y_n406) );
  NAND2_X1 reg_y_U24 ( .A1(reg_y_n404), .A2(reg_y_n403), .ZN(reg_y_n240) );
  NAND2_X1 reg_y_U23 ( .A1(state_y[25]), .A2(reg_y_n451), .ZN(reg_y_n403) );
  NAND2_X1 reg_y_U22 ( .A1(round_inst_aout_y[24]), .A2(reg_y_n440), .ZN(
        reg_y_n404) );
  NAND2_X1 reg_y_U21 ( .A1(reg_y_n402), .A2(reg_y_n401), .ZN(reg_y_n250) );
  NAND2_X1 reg_y_U20 ( .A1(state_y[15]), .A2(reg_y_n451), .ZN(reg_y_n401) );
  NAND2_X1 reg_y_U19 ( .A1(round_inst_aout_y[14]), .A2(reg_y_n456), .ZN(
        reg_y_n402) );
  NAND2_X1 reg_y_U18 ( .A1(reg_y_n400), .A2(reg_y_n399), .ZN(reg_y_n254) );
  NAND2_X1 reg_y_U17 ( .A1(state_y[11]), .A2(reg_y_n451), .ZN(reg_y_n399) );
  NAND2_X1 reg_y_U16 ( .A1(round_inst_aout_y[10]), .A2(reg_y_n440), .ZN(
        reg_y_n400) );
  NAND2_X1 reg_y_U15 ( .A1(reg_y_n398), .A2(reg_y_n397), .ZN(reg_y_n258) );
  NAND2_X1 reg_y_U14 ( .A1(state_y[7]), .A2(reg_y_n451), .ZN(reg_y_n397) );
  NAND2_X1 reg_y_U13 ( .A1(round_inst_aout_y[6]), .A2(reg_y_n456), .ZN(
        reg_y_n398) );
  NAND2_X1 reg_y_U12 ( .A1(reg_y_n396), .A2(reg_y_n395), .ZN(reg_y_n259) );
  NAND2_X1 reg_y_U11 ( .A1(reg_y_n440), .A2(round_inst_aout_y[7]), .ZN(
        reg_y_n395) );
  INV_X1 reg_y_U10 ( .A(reg_y_n462), .ZN(reg_y_n440) );
  INV_X1 reg_y_U9 ( .A(reg_y_n456), .ZN(reg_y_n462) );
  NAND2_X1 reg_y_U8 ( .A1(reg_y_n451), .A2(state_y[6]), .ZN(reg_y_n396) );
  INV_X1 reg_y_U7 ( .A(reg_y_n457), .ZN(reg_y_n451) );
  INV_X1 reg_y_U6 ( .A(reg_y_n421), .ZN(reg_y_n457) );
  INV_X1 reg_y_U5 ( .A(en_sig), .ZN(reg_y_n394) );
  NOR2_X1 reg_y_U4 ( .A1(rst), .A2(reg_y_n394), .ZN(reg_y_n421) );
  NOR2_X1 reg_y_U3 ( .A1(rst), .A2(en_sig), .ZN(reg_y_n456) );
  DFF_X1 reg_y_s_current_state_reg_0_ ( .D(reg_y_n265), .CK(clk), .Q(
        round_inst_srout_y[48]) );
  DFF_X1 reg_y_s_current_state_reg_1_ ( .D(reg_y_n264), .CK(clk), .Q(
        round_inst_aout_y[0]) );
  DFF_X1 reg_y_s_current_state_reg_2_ ( .D(reg_y_n263), .CK(clk), .Q(
        round_inst_aout_y[3]) );
  DFF_X1 reg_y_s_current_state_reg_3_ ( .D(reg_y_n262), .CK(clk), .Q(
        round_inst_aout_y[2]) );
  DFF_X1 reg_y_s_current_state_reg_4_ ( .D(reg_y_n261), .CK(clk), .Q(
        round_inst_srout_y[36]) );
  DFF_X1 reg_y_s_current_state_reg_5_ ( .D(reg_y_n260), .CK(clk), .Q(
        round_inst_aout_y[4]) );
  DFF_X1 reg_y_s_current_state_reg_6_ ( .D(reg_y_n259), .CK(clk), .Q(
        round_inst_aout_y[7]) );
  DFF_X1 reg_y_s_current_state_reg_7_ ( .D(reg_y_n258), .CK(clk), .Q(
        round_inst_aout_y[6]) );
  DFF_X1 reg_y_s_current_state_reg_8_ ( .D(reg_y_n257), .CK(clk), .Q(
        round_inst_srout_y[24]) );
  DFF_X1 reg_y_s_current_state_reg_9_ ( .D(reg_y_n256), .CK(clk), .Q(
        round_inst_aout_y[8]) );
  DFF_X1 reg_y_s_current_state_reg_10_ ( .D(reg_y_n255), .CK(clk), .Q(
        round_inst_aout_y[11]) );
  DFF_X1 reg_y_s_current_state_reg_11_ ( .D(reg_y_n254), .CK(clk), .Q(
        round_inst_aout_y[10]) );
  DFF_X1 reg_y_s_current_state_reg_12_ ( .D(reg_y_n253), .CK(clk), .Q(
        round_inst_srout_y[12]) );
  DFF_X1 reg_y_s_current_state_reg_13_ ( .D(reg_y_n252), .CK(clk), .Q(
        round_inst_aout_y[12]) );
  DFF_X1 reg_y_s_current_state_reg_14_ ( .D(reg_y_n251), .CK(clk), .Q(
        round_inst_aout_y[15]) );
  DFF_X1 reg_y_s_current_state_reg_15_ ( .D(reg_y_n250), .CK(clk), .Q(
        round_inst_aout_y[14]) );
  DFF_X1 reg_y_s_current_state_reg_16_ ( .D(reg_y_n249), .CK(clk), .Q(
        round_inst_srout_y[0]) );
  DFF_X1 reg_y_s_current_state_reg_17_ ( .D(reg_y_n248), .CK(clk), .Q(
        round_inst_aout_y[16]) );
  DFF_X1 reg_y_s_current_state_reg_18_ ( .D(reg_y_n247), .CK(clk), .Q(
        round_inst_aout_y[19]) );
  DFF_X1 reg_y_s_current_state_reg_19_ ( .D(reg_y_n246), .CK(clk), .Q(
        round_inst_aout_y[18]) );
  DFF_X1 reg_y_s_current_state_reg_20_ ( .D(reg_y_n245), .CK(clk), .Q(
        round_inst_srout_y[52]) );
  DFF_X1 reg_y_s_current_state_reg_21_ ( .D(reg_y_n244), .CK(clk), .Q(
        round_inst_aout_y[20]) );
  DFF_X1 reg_y_s_current_state_reg_22_ ( .D(reg_y_n243), .CK(clk), .Q(
        round_inst_aout_y[23]) );
  DFF_X1 reg_y_s_current_state_reg_23_ ( .D(reg_y_n242), .CK(clk), .Q(
        round_inst_aout_y[22]) );
  DFF_X1 reg_y_s_current_state_reg_24_ ( .D(reg_y_n241), .CK(clk), .Q(
        round_inst_srout_y[40]) );
  DFF_X1 reg_y_s_current_state_reg_25_ ( .D(reg_y_n240), .CK(clk), .Q(
        round_inst_aout_y[24]) );
  DFF_X1 reg_y_s_current_state_reg_26_ ( .D(reg_y_n239), .CK(clk), .Q(
        round_inst_aout_y[27]) );
  DFF_X1 reg_y_s_current_state_reg_27_ ( .D(reg_y_n238), .CK(clk), .Q(
        round_inst_aout_y[26]) );
  DFF_X1 reg_y_s_current_state_reg_28_ ( .D(reg_y_n237), .CK(clk), .Q(
        round_inst_srout_y[28]) );
  DFF_X1 reg_y_s_current_state_reg_29_ ( .D(reg_y_n236), .CK(clk), .Q(
        round_inst_aout_y[28]) );
  DFF_X1 reg_y_s_current_state_reg_30_ ( .D(reg_y_n235), .CK(clk), .Q(
        round_inst_aout_y[31]) );
  DFF_X1 reg_y_s_current_state_reg_31_ ( .D(reg_y_n234), .CK(clk), .Q(
        round_inst_aout_y[30]) );
  DFF_X1 reg_y_s_current_state_reg_32_ ( .D(reg_y_n233), .CK(clk), .Q(
        round_inst_srout_y[16]) );
  DFF_X1 reg_y_s_current_state_reg_33_ ( .D(reg_y_n232), .CK(clk), .Q(
        round_inst_aout_y[32]) );
  DFF_X1 reg_y_s_current_state_reg_34_ ( .D(reg_y_n231), .CK(clk), .Q(
        round_inst_aout_y[35]) );
  DFF_X1 reg_y_s_current_state_reg_35_ ( .D(reg_y_n230), .CK(clk), .Q(
        round_inst_aout_y[34]) );
  DFF_X1 reg_y_s_current_state_reg_36_ ( .D(reg_y_n229), .CK(clk), .Q(
        round_inst_srout_y[4]) );
  DFF_X1 reg_y_s_current_state_reg_37_ ( .D(reg_y_n228), .CK(clk), .Q(
        round_inst_aout_y[36]) );
  DFF_X1 reg_y_s_current_state_reg_38_ ( .D(reg_y_n227), .CK(clk), .Q(
        round_inst_aout_y[39]) );
  DFF_X1 reg_y_s_current_state_reg_39_ ( .D(reg_y_n226), .CK(clk), .Q(
        round_inst_aout_y[38]) );
  DFF_X1 reg_y_s_current_state_reg_40_ ( .D(reg_y_n225), .CK(clk), .Q(
        round_inst_srout_y[56]) );
  DFF_X1 reg_y_s_current_state_reg_41_ ( .D(reg_y_n224), .CK(clk), .Q(
        round_inst_aout_y[40]) );
  DFF_X1 reg_y_s_current_state_reg_42_ ( .D(reg_y_n223), .CK(clk), .Q(
        round_inst_aout_y[43]) );
  DFF_X1 reg_y_s_current_state_reg_43_ ( .D(reg_y_n222), .CK(clk), .Q(
        round_inst_aout_y[42]) );
  DFF_X1 reg_y_s_current_state_reg_44_ ( .D(reg_y_n221), .CK(clk), .Q(
        round_inst_srout_y[44]) );
  DFF_X1 reg_y_s_current_state_reg_45_ ( .D(reg_y_n220), .CK(clk), .Q(
        round_inst_aout_y[44]) );
  DFF_X1 reg_y_s_current_state_reg_46_ ( .D(reg_y_n219), .CK(clk), .Q(
        round_inst_aout_y[47]) );
  DFF_X1 reg_y_s_current_state_reg_47_ ( .D(reg_y_n218), .CK(clk), .Q(
        round_inst_aout_y[46]) );
  DFF_X1 reg_y_s_current_state_reg_48_ ( .D(reg_y_n217), .CK(clk), .Q(
        round_inst_srout_y[32]) );
  DFF_X1 reg_y_s_current_state_reg_49_ ( .D(reg_y_n216), .CK(clk), .Q(
        round_inst_aout_y[48]) );
  DFF_X1 reg_y_s_current_state_reg_50_ ( .D(reg_y_n215), .CK(clk), .Q(
        round_inst_aout_y[51]) );
  DFF_X1 reg_y_s_current_state_reg_51_ ( .D(reg_y_n214), .CK(clk), .Q(
        round_inst_aout_y[50]) );
  DFF_X1 reg_y_s_current_state_reg_52_ ( .D(reg_y_n213), .CK(clk), .Q(
        round_inst_srout_y[20]) );
  DFF_X1 reg_y_s_current_state_reg_53_ ( .D(reg_y_n212), .CK(clk), .Q(
        round_inst_aout_y[52]) );
  DFF_X1 reg_y_s_current_state_reg_54_ ( .D(reg_y_n211), .CK(clk), .Q(
        round_inst_aout_y[55]) );
  DFF_X1 reg_y_s_current_state_reg_55_ ( .D(reg_y_n210), .CK(clk), .Q(
        round_inst_aout_y[54]) );
  DFF_X1 reg_y_s_current_state_reg_56_ ( .D(reg_y_n209), .CK(clk), .Q(
        round_inst_srout_y[8]) );
  DFF_X1 reg_y_s_current_state_reg_57_ ( .D(reg_y_n208), .CK(clk), .Q(
        round_inst_aout_y[56]) );
  DFF_X1 reg_y_s_current_state_reg_58_ ( .D(reg_y_n207), .CK(clk), .Q(
        round_inst_aout_y[59]) );
  DFF_X1 reg_y_s_current_state_reg_59_ ( .D(reg_y_n206), .CK(clk), .Q(
        round_inst_aout_y[58]) );
  DFF_X1 reg_y_s_current_state_reg_60_ ( .D(reg_y_n205), .CK(clk), .Q(
        round_inst_srout_y[60]) );
  DFF_X1 reg_y_s_current_state_reg_61_ ( .D(reg_y_n204), .CK(clk), .Q(
        round_inst_aout_y[60]) );
  DFF_X1 reg_y_s_current_state_reg_62_ ( .D(reg_y_n203), .CK(clk), .Q(
        round_inst_aout_y[63]) );
  DFF_X1 reg_y_s_current_state_reg_63_ ( .D(reg_y_n202), .CK(clk), .Q(
        round_inst_aout_y[62]) );
  NAND2_X1 reg_z_U205 ( .A1(reg_z_n532), .A2(reg_z_n531), .ZN(reg_z_n231) );
  NAND2_X1 reg_z_U204 ( .A1(state_z[34]), .A2(reg_z_n530), .ZN(reg_z_n531) );
  NAND2_X1 reg_z_U203 ( .A1(round_inst_aout_z[35]), .A2(reg_z_n529), .ZN(
        reg_z_n532) );
  NAND2_X1 reg_z_U202 ( .A1(reg_z_n528), .A2(reg_z_n527), .ZN(reg_z_n232) );
  NAND2_X1 reg_z_U201 ( .A1(state_z[33]), .A2(reg_z_n530), .ZN(reg_z_n527) );
  NAND2_X1 reg_z_U200 ( .A1(round_inst_aout_z[32]), .A2(reg_z_n529), .ZN(
        reg_z_n528) );
  NAND2_X1 reg_z_U199 ( .A1(reg_z_n526), .A2(reg_z_n525), .ZN(reg_z_n235) );
  NAND2_X1 reg_z_U198 ( .A1(state_z[30]), .A2(reg_z_n530), .ZN(reg_z_n525) );
  NAND2_X1 reg_z_U197 ( .A1(round_inst_aout_z[31]), .A2(reg_z_n529), .ZN(
        reg_z_n526) );
  NAND2_X1 reg_z_U196 ( .A1(reg_z_n524), .A2(reg_z_n523), .ZN(reg_z_n236) );
  NAND2_X1 reg_z_U195 ( .A1(state_z[29]), .A2(reg_z_n530), .ZN(reg_z_n523) );
  NAND2_X1 reg_z_U194 ( .A1(round_inst_aout_z[28]), .A2(reg_z_n529), .ZN(
        reg_z_n524) );
  NAND2_X1 reg_z_U193 ( .A1(reg_z_n522), .A2(reg_z_n521), .ZN(reg_z_n237) );
  NAND2_X1 reg_z_U192 ( .A1(state_z[28]), .A2(reg_z_n530), .ZN(reg_z_n521) );
  NAND2_X1 reg_z_U191 ( .A1(round_inst_srout_z[28]), .A2(reg_z_n529), .ZN(
        reg_z_n522) );
  NAND2_X1 reg_z_U190 ( .A1(reg_z_n520), .A2(reg_z_n519), .ZN(reg_z_n238) );
  NAND2_X1 reg_z_U189 ( .A1(state_z[27]), .A2(reg_z_n530), .ZN(reg_z_n519) );
  NAND2_X1 reg_z_U188 ( .A1(round_inst_aout_z[26]), .A2(reg_z_n529), .ZN(
        reg_z_n520) );
  NAND2_X1 reg_z_U187 ( .A1(reg_z_n518), .A2(reg_z_n517), .ZN(reg_z_n239) );
  NAND2_X1 reg_z_U186 ( .A1(state_z[26]), .A2(reg_z_n530), .ZN(reg_z_n517) );
  NAND2_X1 reg_z_U185 ( .A1(round_inst_aout_z[27]), .A2(reg_z_n529), .ZN(
        reg_z_n518) );
  NAND2_X1 reg_z_U184 ( .A1(reg_z_n516), .A2(reg_z_n515), .ZN(reg_z_n240) );
  NAND2_X1 reg_z_U183 ( .A1(state_z[25]), .A2(reg_z_n530), .ZN(reg_z_n515) );
  NAND2_X1 reg_z_U182 ( .A1(round_inst_aout_z[24]), .A2(reg_z_n529), .ZN(
        reg_z_n516) );
  NAND2_X1 reg_z_U181 ( .A1(reg_z_n514), .A2(reg_z_n513), .ZN(reg_z_n241) );
  NAND2_X1 reg_z_U180 ( .A1(state_z[24]), .A2(reg_z_n530), .ZN(reg_z_n513) );
  NAND2_X1 reg_z_U179 ( .A1(round_inst_srout_z[40]), .A2(reg_z_n529), .ZN(
        reg_z_n514) );
  NAND2_X1 reg_z_U178 ( .A1(reg_z_n512), .A2(reg_z_n511), .ZN(reg_z_n242) );
  NAND2_X1 reg_z_U177 ( .A1(state_z[23]), .A2(reg_z_n530), .ZN(reg_z_n511) );
  NAND2_X1 reg_z_U176 ( .A1(round_inst_aout_z[22]), .A2(reg_z_n529), .ZN(
        reg_z_n512) );
  NAND2_X1 reg_z_U175 ( .A1(reg_z_n510), .A2(reg_z_n509), .ZN(reg_z_n244) );
  NAND2_X1 reg_z_U174 ( .A1(state_z[21]), .A2(reg_z_n530), .ZN(reg_z_n509) );
  NAND2_X1 reg_z_U173 ( .A1(round_inst_aout_z[20]), .A2(reg_z_n529), .ZN(
        reg_z_n510) );
  NAND2_X1 reg_z_U172 ( .A1(reg_z_n508), .A2(reg_z_n507), .ZN(reg_z_n246) );
  NAND2_X1 reg_z_U171 ( .A1(state_z[19]), .A2(reg_z_n530), .ZN(reg_z_n507) );
  NAND2_X1 reg_z_U170 ( .A1(round_inst_aout_z[18]), .A2(reg_z_n529), .ZN(
        reg_z_n508) );
  NAND2_X1 reg_z_U169 ( .A1(reg_z_n506), .A2(reg_z_n505), .ZN(reg_z_n247) );
  NAND2_X1 reg_z_U168 ( .A1(state_z[18]), .A2(reg_z_n504), .ZN(reg_z_n505) );
  NAND2_X1 reg_z_U167 ( .A1(round_inst_aout_z[19]), .A2(reg_z_n503), .ZN(
        reg_z_n506) );
  NAND2_X1 reg_z_U166 ( .A1(reg_z_n502), .A2(reg_z_n501), .ZN(reg_z_n248) );
  NAND2_X1 reg_z_U165 ( .A1(state_z[17]), .A2(reg_z_n504), .ZN(reg_z_n501) );
  NAND2_X1 reg_z_U164 ( .A1(round_inst_aout_z[16]), .A2(reg_z_n503), .ZN(
        reg_z_n502) );
  NAND2_X1 reg_z_U163 ( .A1(reg_z_n500), .A2(reg_z_n499), .ZN(reg_z_n250) );
  NAND2_X1 reg_z_U162 ( .A1(state_z[15]), .A2(reg_z_n504), .ZN(reg_z_n499) );
  NAND2_X1 reg_z_U161 ( .A1(round_inst_aout_z[14]), .A2(reg_z_n503), .ZN(
        reg_z_n500) );
  NAND2_X1 reg_z_U160 ( .A1(reg_z_n498), .A2(reg_z_n497), .ZN(reg_z_n251) );
  NAND2_X1 reg_z_U159 ( .A1(state_z[14]), .A2(reg_z_n504), .ZN(reg_z_n497) );
  NAND2_X1 reg_z_U158 ( .A1(round_inst_aout_z[15]), .A2(reg_z_n503), .ZN(
        reg_z_n498) );
  NAND2_X1 reg_z_U157 ( .A1(reg_z_n496), .A2(reg_z_n495), .ZN(reg_z_n252) );
  NAND2_X1 reg_z_U156 ( .A1(state_z[13]), .A2(reg_z_n504), .ZN(reg_z_n495) );
  NAND2_X1 reg_z_U155 ( .A1(round_inst_aout_z[12]), .A2(reg_z_n503), .ZN(
        reg_z_n496) );
  NAND2_X1 reg_z_U154 ( .A1(reg_z_n494), .A2(reg_z_n493), .ZN(reg_z_n253) );
  NAND2_X1 reg_z_U153 ( .A1(state_z[12]), .A2(reg_z_n504), .ZN(reg_z_n493) );
  NAND2_X1 reg_z_U152 ( .A1(round_inst_srout_z[12]), .A2(reg_z_n503), .ZN(
        reg_z_n494) );
  NAND2_X1 reg_z_U151 ( .A1(reg_z_n492), .A2(reg_z_n491), .ZN(reg_z_n254) );
  NAND2_X1 reg_z_U150 ( .A1(state_z[11]), .A2(reg_z_n504), .ZN(reg_z_n491) );
  NAND2_X1 reg_z_U149 ( .A1(round_inst_aout_z[10]), .A2(reg_z_n503), .ZN(
        reg_z_n492) );
  NAND2_X1 reg_z_U148 ( .A1(reg_z_n490), .A2(reg_z_n489), .ZN(reg_z_n255) );
  NAND2_X1 reg_z_U147 ( .A1(state_z[10]), .A2(reg_z_n504), .ZN(reg_z_n489) );
  NAND2_X1 reg_z_U146 ( .A1(round_inst_aout_z[11]), .A2(reg_z_n503), .ZN(
        reg_z_n490) );
  NAND2_X1 reg_z_U145 ( .A1(reg_z_n488), .A2(reg_z_n487), .ZN(reg_z_n256) );
  NAND2_X1 reg_z_U144 ( .A1(state_z[9]), .A2(reg_z_n504), .ZN(reg_z_n487) );
  NAND2_X1 reg_z_U143 ( .A1(round_inst_aout_z[8]), .A2(reg_z_n503), .ZN(
        reg_z_n488) );
  NAND2_X1 reg_z_U142 ( .A1(reg_z_n486), .A2(reg_z_n485), .ZN(reg_z_n257) );
  NAND2_X1 reg_z_U141 ( .A1(state_z[8]), .A2(reg_z_n504), .ZN(reg_z_n485) );
  NAND2_X1 reg_z_U140 ( .A1(round_inst_srout_z[24]), .A2(reg_z_n503), .ZN(
        reg_z_n486) );
  NAND2_X1 reg_z_U139 ( .A1(reg_z_n484), .A2(reg_z_n483), .ZN(reg_z_n258) );
  NAND2_X1 reg_z_U138 ( .A1(state_z[7]), .A2(reg_z_n504), .ZN(reg_z_n483) );
  NAND2_X1 reg_z_U137 ( .A1(round_inst_aout_z[6]), .A2(reg_z_n503), .ZN(
        reg_z_n484) );
  NAND2_X1 reg_z_U136 ( .A1(reg_z_n482), .A2(reg_z_n481), .ZN(reg_z_n259) );
  NAND2_X1 reg_z_U135 ( .A1(state_z[6]), .A2(reg_z_n504), .ZN(reg_z_n481) );
  NAND2_X1 reg_z_U134 ( .A1(round_inst_aout_z[7]), .A2(reg_z_n503), .ZN(
        reg_z_n482) );
  NAND2_X1 reg_z_U133 ( .A1(reg_z_n480), .A2(reg_z_n479), .ZN(reg_z_n260) );
  NAND2_X1 reg_z_U132 ( .A1(state_z[5]), .A2(reg_z_n504), .ZN(reg_z_n479) );
  NAND2_X1 reg_z_U131 ( .A1(round_inst_aout_z[4]), .A2(reg_z_n503), .ZN(
        reg_z_n480) );
  NAND2_X1 reg_z_U130 ( .A1(reg_z_n478), .A2(reg_z_n477), .ZN(reg_z_n261) );
  NAND2_X1 reg_z_U129 ( .A1(state_z[4]), .A2(reg_z_n530), .ZN(reg_z_n477) );
  NAND2_X1 reg_z_U128 ( .A1(round_inst_srout_z[36]), .A2(reg_z_n529), .ZN(
        reg_z_n478) );
  NAND2_X1 reg_z_U127 ( .A1(reg_z_n476), .A2(reg_z_n475), .ZN(reg_z_n262) );
  NAND2_X1 reg_z_U126 ( .A1(state_z[3]), .A2(reg_z_n504), .ZN(reg_z_n475) );
  NAND2_X1 reg_z_U125 ( .A1(round_inst_aout_z[2]), .A2(reg_z_n503), .ZN(
        reg_z_n476) );
  NAND2_X1 reg_z_U124 ( .A1(reg_z_n474), .A2(reg_z_n473), .ZN(reg_z_n263) );
  NAND2_X1 reg_z_U123 ( .A1(state_z[2]), .A2(reg_z_n530), .ZN(reg_z_n473) );
  NAND2_X1 reg_z_U122 ( .A1(round_inst_aout_z[3]), .A2(reg_z_n529), .ZN(
        reg_z_n474) );
  NAND2_X1 reg_z_U121 ( .A1(reg_z_n472), .A2(reg_z_n471), .ZN(reg_z_n265) );
  NAND2_X1 reg_z_U120 ( .A1(state_z[0]), .A2(reg_z_n504), .ZN(reg_z_n471) );
  NAND2_X1 reg_z_U119 ( .A1(round_inst_srout_z[48]), .A2(reg_z_n503), .ZN(
        reg_z_n472) );
  NAND2_X1 reg_z_U118 ( .A1(reg_z_n470), .A2(reg_z_n469), .ZN(reg_z_n206) );
  NAND2_X1 reg_z_U117 ( .A1(state_z[59]), .A2(reg_z_n530), .ZN(reg_z_n469) );
  NAND2_X1 reg_z_U116 ( .A1(round_inst_aout_z[58]), .A2(reg_z_n529), .ZN(
        reg_z_n470) );
  NAND2_X1 reg_z_U115 ( .A1(reg_z_n468), .A2(reg_z_n467), .ZN(reg_z_n207) );
  NAND2_X1 reg_z_U114 ( .A1(state_z[58]), .A2(reg_z_n504), .ZN(reg_z_n467) );
  NAND2_X1 reg_z_U113 ( .A1(round_inst_aout_z[59]), .A2(reg_z_n503), .ZN(
        reg_z_n468) );
  NAND2_X1 reg_z_U112 ( .A1(reg_z_n466), .A2(reg_z_n465), .ZN(reg_z_n208) );
  NAND2_X1 reg_z_U111 ( .A1(state_z[57]), .A2(reg_z_n530), .ZN(reg_z_n465) );
  NAND2_X1 reg_z_U110 ( .A1(round_inst_aout_z[56]), .A2(reg_z_n529), .ZN(
        reg_z_n466) );
  NAND2_X1 reg_z_U109 ( .A1(reg_z_n464), .A2(reg_z_n463), .ZN(reg_z_n209) );
  NAND2_X1 reg_z_U108 ( .A1(state_z[56]), .A2(reg_z_n504), .ZN(reg_z_n463) );
  NAND2_X1 reg_z_U107 ( .A1(round_inst_srout_z[8]), .A2(reg_z_n503), .ZN(
        reg_z_n464) );
  INV_X1 reg_z_U106 ( .A(reg_z_n462), .ZN(reg_z_n503) );
  NAND2_X1 reg_z_U105 ( .A1(reg_z_n461), .A2(reg_z_n460), .ZN(reg_z_n210) );
  NAND2_X1 reg_z_U104 ( .A1(state_z[55]), .A2(reg_z_n530), .ZN(reg_z_n460) );
  NAND2_X1 reg_z_U103 ( .A1(round_inst_aout_z[54]), .A2(reg_z_n529), .ZN(
        reg_z_n461) );
  INV_X1 reg_z_U102 ( .A(reg_z_n462), .ZN(reg_z_n529) );
  NAND2_X1 reg_z_U101 ( .A1(reg_z_n459), .A2(reg_z_n458), .ZN(reg_z_n211) );
  NAND2_X1 reg_z_U100 ( .A1(state_z[54]), .A2(reg_z_n504), .ZN(reg_z_n458) );
  INV_X1 reg_z_U99 ( .A(reg_z_n457), .ZN(reg_z_n504) );
  NAND2_X1 reg_z_U98 ( .A1(round_inst_aout_z[55]), .A2(reg_z_n456), .ZN(
        reg_z_n459) );
  NAND2_X1 reg_z_U97 ( .A1(reg_z_n455), .A2(reg_z_n454), .ZN(reg_z_n212) );
  NAND2_X1 reg_z_U96 ( .A1(state_z[53]), .A2(reg_z_n530), .ZN(reg_z_n454) );
  INV_X1 reg_z_U95 ( .A(reg_z_n457), .ZN(reg_z_n530) );
  NAND2_X1 reg_z_U94 ( .A1(round_inst_aout_z[52]), .A2(reg_z_n456), .ZN(
        reg_z_n455) );
  NAND2_X1 reg_z_U93 ( .A1(reg_z_n453), .A2(reg_z_n452), .ZN(reg_z_n213) );
  NAND2_X1 reg_z_U92 ( .A1(state_z[52]), .A2(reg_z_n451), .ZN(reg_z_n452) );
  NAND2_X1 reg_z_U91 ( .A1(round_inst_srout_z[20]), .A2(reg_z_n456), .ZN(
        reg_z_n453) );
  NAND2_X1 reg_z_U90 ( .A1(reg_z_n450), .A2(reg_z_n449), .ZN(reg_z_n214) );
  NAND2_X1 reg_z_U89 ( .A1(state_z[51]), .A2(reg_z_n451), .ZN(reg_z_n449) );
  NAND2_X1 reg_z_U88 ( .A1(round_inst_aout_z[50]), .A2(reg_z_n456), .ZN(
        reg_z_n450) );
  NAND2_X1 reg_z_U87 ( .A1(reg_z_n448), .A2(reg_z_n447), .ZN(reg_z_n215) );
  NAND2_X1 reg_z_U86 ( .A1(state_z[50]), .A2(reg_z_n451), .ZN(reg_z_n447) );
  NAND2_X1 reg_z_U85 ( .A1(round_inst_aout_z[51]), .A2(reg_z_n456), .ZN(
        reg_z_n448) );
  NAND2_X1 reg_z_U84 ( .A1(reg_z_n446), .A2(reg_z_n445), .ZN(reg_z_n216) );
  NAND2_X1 reg_z_U83 ( .A1(state_z[49]), .A2(reg_z_n451), .ZN(reg_z_n445) );
  NAND2_X1 reg_z_U82 ( .A1(round_inst_aout_z[48]), .A2(reg_z_n456), .ZN(
        reg_z_n446) );
  NAND2_X1 reg_z_U81 ( .A1(reg_z_n444), .A2(reg_z_n443), .ZN(reg_z_n217) );
  NAND2_X1 reg_z_U80 ( .A1(state_z[48]), .A2(reg_z_n451), .ZN(reg_z_n443) );
  NAND2_X1 reg_z_U79 ( .A1(round_inst_srout_z[32]), .A2(reg_z_n456), .ZN(
        reg_z_n444) );
  NAND2_X1 reg_z_U78 ( .A1(reg_z_n442), .A2(reg_z_n441), .ZN(reg_z_n218) );
  NAND2_X1 reg_z_U77 ( .A1(state_z[47]), .A2(reg_z_n451), .ZN(reg_z_n441) );
  NAND2_X1 reg_z_U76 ( .A1(round_inst_aout_z[46]), .A2(reg_z_n440), .ZN(
        reg_z_n442) );
  NAND2_X1 reg_z_U75 ( .A1(reg_z_n439), .A2(reg_z_n438), .ZN(reg_z_n219) );
  NAND2_X1 reg_z_U74 ( .A1(state_z[46]), .A2(reg_z_n451), .ZN(reg_z_n438) );
  NAND2_X1 reg_z_U73 ( .A1(round_inst_aout_z[47]), .A2(reg_z_n440), .ZN(
        reg_z_n439) );
  NAND2_X1 reg_z_U72 ( .A1(reg_z_n437), .A2(reg_z_n436), .ZN(reg_z_n220) );
  NAND2_X1 reg_z_U71 ( .A1(state_z[45]), .A2(reg_z_n451), .ZN(reg_z_n436) );
  NAND2_X1 reg_z_U70 ( .A1(round_inst_aout_z[44]), .A2(reg_z_n440), .ZN(
        reg_z_n437) );
  NAND2_X1 reg_z_U69 ( .A1(reg_z_n435), .A2(reg_z_n434), .ZN(reg_z_n221) );
  NAND2_X1 reg_z_U68 ( .A1(state_z[44]), .A2(reg_z_n451), .ZN(reg_z_n434) );
  NAND2_X1 reg_z_U67 ( .A1(round_inst_srout_z[44]), .A2(reg_z_n440), .ZN(
        reg_z_n435) );
  NAND2_X1 reg_z_U66 ( .A1(reg_z_n433), .A2(reg_z_n432), .ZN(reg_z_n222) );
  NAND2_X1 reg_z_U65 ( .A1(state_z[43]), .A2(reg_z_n451), .ZN(reg_z_n432) );
  NAND2_X1 reg_z_U64 ( .A1(round_inst_aout_z[42]), .A2(reg_z_n440), .ZN(
        reg_z_n433) );
  NAND2_X1 reg_z_U63 ( .A1(reg_z_n431), .A2(reg_z_n430), .ZN(reg_z_n223) );
  NAND2_X1 reg_z_U62 ( .A1(state_z[42]), .A2(reg_z_n451), .ZN(reg_z_n430) );
  NAND2_X1 reg_z_U61 ( .A1(round_inst_aout_z[43]), .A2(reg_z_n440), .ZN(
        reg_z_n431) );
  NAND2_X1 reg_z_U60 ( .A1(reg_z_n429), .A2(reg_z_n428), .ZN(reg_z_n224) );
  NAND2_X1 reg_z_U59 ( .A1(state_z[41]), .A2(reg_z_n451), .ZN(reg_z_n428) );
  NAND2_X1 reg_z_U58 ( .A1(round_inst_aout_z[40]), .A2(reg_z_n440), .ZN(
        reg_z_n429) );
  NAND2_X1 reg_z_U57 ( .A1(reg_z_n427), .A2(reg_z_n426), .ZN(reg_z_n225) );
  NAND2_X1 reg_z_U56 ( .A1(state_z[40]), .A2(reg_z_n451), .ZN(reg_z_n426) );
  NAND2_X1 reg_z_U55 ( .A1(round_inst_srout_z[56]), .A2(reg_z_n440), .ZN(
        reg_z_n427) );
  NAND2_X1 reg_z_U54 ( .A1(reg_z_n425), .A2(reg_z_n424), .ZN(reg_z_n226) );
  NAND2_X1 reg_z_U53 ( .A1(state_z[39]), .A2(reg_z_n451), .ZN(reg_z_n424) );
  NAND2_X1 reg_z_U52 ( .A1(round_inst_aout_z[38]), .A2(reg_z_n440), .ZN(
        reg_z_n425) );
  NAND2_X1 reg_z_U51 ( .A1(reg_z_n423), .A2(reg_z_n422), .ZN(reg_z_n227) );
  NAND2_X1 reg_z_U50 ( .A1(state_z[38]), .A2(reg_z_n421), .ZN(reg_z_n422) );
  NAND2_X1 reg_z_U49 ( .A1(round_inst_aout_z[39]), .A2(reg_z_n440), .ZN(
        reg_z_n423) );
  NAND2_X1 reg_z_U48 ( .A1(reg_z_n420), .A2(reg_z_n419), .ZN(reg_z_n228) );
  NAND2_X1 reg_z_U47 ( .A1(state_z[37]), .A2(reg_z_n421), .ZN(reg_z_n419) );
  NAND2_X1 reg_z_U46 ( .A1(round_inst_aout_z[36]), .A2(reg_z_n440), .ZN(
        reg_z_n420) );
  NAND2_X1 reg_z_U45 ( .A1(reg_z_n418), .A2(reg_z_n417), .ZN(reg_z_n229) );
  NAND2_X1 reg_z_U44 ( .A1(state_z[36]), .A2(reg_z_n421), .ZN(reg_z_n417) );
  NAND2_X1 reg_z_U43 ( .A1(round_inst_srout_z[4]), .A2(reg_z_n440), .ZN(
        reg_z_n418) );
  NAND2_X1 reg_z_U42 ( .A1(reg_z_n416), .A2(reg_z_n415), .ZN(reg_z_n202) );
  NAND2_X1 reg_z_U41 ( .A1(state_z[63]), .A2(reg_z_n421), .ZN(reg_z_n415) );
  NAND2_X1 reg_z_U40 ( .A1(round_inst_aout_z[62]), .A2(reg_z_n440), .ZN(
        reg_z_n416) );
  NAND2_X1 reg_z_U39 ( .A1(reg_z_n414), .A2(reg_z_n413), .ZN(reg_z_n203) );
  NAND2_X1 reg_z_U38 ( .A1(state_z[62]), .A2(reg_z_n421), .ZN(reg_z_n413) );
  NAND2_X1 reg_z_U37 ( .A1(round_inst_aout_z[63]), .A2(reg_z_n440), .ZN(
        reg_z_n414) );
  NAND2_X1 reg_z_U36 ( .A1(reg_z_n412), .A2(reg_z_n411), .ZN(reg_z_n204) );
  NAND2_X1 reg_z_U35 ( .A1(state_z[61]), .A2(reg_z_n421), .ZN(reg_z_n411) );
  NAND2_X1 reg_z_U34 ( .A1(round_inst_aout_z[60]), .A2(reg_z_n440), .ZN(
        reg_z_n412) );
  NAND2_X1 reg_z_U33 ( .A1(reg_z_n410), .A2(reg_z_n409), .ZN(reg_z_n205) );
  NAND2_X1 reg_z_U32 ( .A1(state_z[60]), .A2(reg_z_n421), .ZN(reg_z_n409) );
  NAND2_X1 reg_z_U31 ( .A1(round_inst_srout_z[60]), .A2(reg_z_n440), .ZN(
        reg_z_n410) );
  NAND2_X1 reg_z_U30 ( .A1(reg_z_n408), .A2(reg_z_n407), .ZN(reg_z_n230) );
  NAND2_X1 reg_z_U29 ( .A1(state_z[35]), .A2(reg_z_n421), .ZN(reg_z_n407) );
  NAND2_X1 reg_z_U28 ( .A1(round_inst_aout_z[34]), .A2(reg_z_n440), .ZN(
        reg_z_n408) );
  NAND2_X1 reg_z_U27 ( .A1(reg_z_n406), .A2(reg_z_n405), .ZN(reg_z_n233) );
  NAND2_X1 reg_z_U26 ( .A1(state_z[32]), .A2(reg_z_n421), .ZN(reg_z_n405) );
  NAND2_X1 reg_z_U25 ( .A1(round_inst_srout_z[16]), .A2(reg_z_n440), .ZN(
        reg_z_n406) );
  NAND2_X1 reg_z_U24 ( .A1(reg_z_n404), .A2(reg_z_n403), .ZN(reg_z_n234) );
  NAND2_X1 reg_z_U23 ( .A1(state_z[31]), .A2(reg_z_n451), .ZN(reg_z_n403) );
  NAND2_X1 reg_z_U22 ( .A1(round_inst_aout_z[30]), .A2(reg_z_n440), .ZN(
        reg_z_n404) );
  NAND2_X1 reg_z_U21 ( .A1(reg_z_n402), .A2(reg_z_n401), .ZN(reg_z_n243) );
  NAND2_X1 reg_z_U20 ( .A1(state_z[22]), .A2(reg_z_n451), .ZN(reg_z_n401) );
  NAND2_X1 reg_z_U19 ( .A1(round_inst_aout_z[23]), .A2(reg_z_n456), .ZN(
        reg_z_n402) );
  NAND2_X1 reg_z_U18 ( .A1(reg_z_n400), .A2(reg_z_n399), .ZN(reg_z_n245) );
  NAND2_X1 reg_z_U17 ( .A1(state_z[20]), .A2(reg_z_n451), .ZN(reg_z_n399) );
  NAND2_X1 reg_z_U16 ( .A1(round_inst_srout_z[52]), .A2(reg_z_n440), .ZN(
        reg_z_n400) );
  NAND2_X1 reg_z_U15 ( .A1(reg_z_n398), .A2(reg_z_n397), .ZN(reg_z_n249) );
  NAND2_X1 reg_z_U14 ( .A1(state_z[16]), .A2(reg_z_n451), .ZN(reg_z_n397) );
  NAND2_X1 reg_z_U13 ( .A1(round_inst_srout_z[0]), .A2(reg_z_n456), .ZN(
        reg_z_n398) );
  NAND2_X1 reg_z_U12 ( .A1(reg_z_n396), .A2(reg_z_n395), .ZN(reg_z_n264) );
  NAND2_X1 reg_z_U11 ( .A1(reg_z_n440), .A2(round_inst_aout_z[0]), .ZN(
        reg_z_n395) );
  INV_X1 reg_z_U10 ( .A(reg_z_n462), .ZN(reg_z_n440) );
  INV_X1 reg_z_U9 ( .A(reg_z_n456), .ZN(reg_z_n462) );
  NAND2_X1 reg_z_U8 ( .A1(reg_z_n451), .A2(state_z[1]), .ZN(reg_z_n396) );
  INV_X1 reg_z_U7 ( .A(reg_z_n457), .ZN(reg_z_n451) );
  INV_X1 reg_z_U6 ( .A(reg_z_n421), .ZN(reg_z_n457) );
  INV_X1 reg_z_U5 ( .A(en_sig), .ZN(reg_z_n394) );
  NOR2_X1 reg_z_U4 ( .A1(rst), .A2(reg_z_n394), .ZN(reg_z_n421) );
  NOR2_X1 reg_z_U3 ( .A1(rst), .A2(en_sig), .ZN(reg_z_n456) );
  DFF_X1 reg_z_s_current_state_reg_0_ ( .D(reg_z_n265), .CK(clk), .Q(
        round_inst_srout_z[48]) );
  DFF_X1 reg_z_s_current_state_reg_1_ ( .D(reg_z_n264), .CK(clk), .Q(
        round_inst_aout_z[0]) );
  DFF_X1 reg_z_s_current_state_reg_2_ ( .D(reg_z_n263), .CK(clk), .Q(
        round_inst_aout_z[3]) );
  DFF_X1 reg_z_s_current_state_reg_3_ ( .D(reg_z_n262), .CK(clk), .Q(
        round_inst_aout_z[2]) );
  DFF_X1 reg_z_s_current_state_reg_4_ ( .D(reg_z_n261), .CK(clk), .Q(
        round_inst_srout_z[36]) );
  DFF_X1 reg_z_s_current_state_reg_5_ ( .D(reg_z_n260), .CK(clk), .Q(
        round_inst_aout_z[4]) );
  DFF_X1 reg_z_s_current_state_reg_6_ ( .D(reg_z_n259), .CK(clk), .Q(
        round_inst_aout_z[7]) );
  DFF_X1 reg_z_s_current_state_reg_7_ ( .D(reg_z_n258), .CK(clk), .Q(
        round_inst_aout_z[6]) );
  DFF_X1 reg_z_s_current_state_reg_8_ ( .D(reg_z_n257), .CK(clk), .Q(
        round_inst_srout_z[24]) );
  DFF_X1 reg_z_s_current_state_reg_9_ ( .D(reg_z_n256), .CK(clk), .Q(
        round_inst_aout_z[8]) );
  DFF_X1 reg_z_s_current_state_reg_10_ ( .D(reg_z_n255), .CK(clk), .Q(
        round_inst_aout_z[11]) );
  DFF_X1 reg_z_s_current_state_reg_11_ ( .D(reg_z_n254), .CK(clk), .Q(
        round_inst_aout_z[10]) );
  DFF_X1 reg_z_s_current_state_reg_12_ ( .D(reg_z_n253), .CK(clk), .Q(
        round_inst_srout_z[12]) );
  DFF_X1 reg_z_s_current_state_reg_13_ ( .D(reg_z_n252), .CK(clk), .Q(
        round_inst_aout_z[12]) );
  DFF_X1 reg_z_s_current_state_reg_14_ ( .D(reg_z_n251), .CK(clk), .Q(
        round_inst_aout_z[15]) );
  DFF_X1 reg_z_s_current_state_reg_15_ ( .D(reg_z_n250), .CK(clk), .Q(
        round_inst_aout_z[14]) );
  DFF_X1 reg_z_s_current_state_reg_16_ ( .D(reg_z_n249), .CK(clk), .Q(
        round_inst_srout_z[0]) );
  DFF_X1 reg_z_s_current_state_reg_17_ ( .D(reg_z_n248), .CK(clk), .Q(
        round_inst_aout_z[16]) );
  DFF_X1 reg_z_s_current_state_reg_18_ ( .D(reg_z_n247), .CK(clk), .Q(
        round_inst_aout_z[19]) );
  DFF_X1 reg_z_s_current_state_reg_19_ ( .D(reg_z_n246), .CK(clk), .Q(
        round_inst_aout_z[18]) );
  DFF_X1 reg_z_s_current_state_reg_20_ ( .D(reg_z_n245), .CK(clk), .Q(
        round_inst_srout_z[52]) );
  DFF_X1 reg_z_s_current_state_reg_21_ ( .D(reg_z_n244), .CK(clk), .Q(
        round_inst_aout_z[20]) );
  DFF_X1 reg_z_s_current_state_reg_22_ ( .D(reg_z_n243), .CK(clk), .Q(
        round_inst_aout_z[23]) );
  DFF_X1 reg_z_s_current_state_reg_23_ ( .D(reg_z_n242), .CK(clk), .Q(
        round_inst_aout_z[22]) );
  DFF_X1 reg_z_s_current_state_reg_24_ ( .D(reg_z_n241), .CK(clk), .Q(
        round_inst_srout_z[40]) );
  DFF_X1 reg_z_s_current_state_reg_25_ ( .D(reg_z_n240), .CK(clk), .Q(
        round_inst_aout_z[24]) );
  DFF_X1 reg_z_s_current_state_reg_26_ ( .D(reg_z_n239), .CK(clk), .Q(
        round_inst_aout_z[27]) );
  DFF_X1 reg_z_s_current_state_reg_27_ ( .D(reg_z_n238), .CK(clk), .Q(
        round_inst_aout_z[26]) );
  DFF_X1 reg_z_s_current_state_reg_28_ ( .D(reg_z_n237), .CK(clk), .Q(
        round_inst_srout_z[28]) );
  DFF_X1 reg_z_s_current_state_reg_29_ ( .D(reg_z_n236), .CK(clk), .Q(
        round_inst_aout_z[28]) );
  DFF_X1 reg_z_s_current_state_reg_30_ ( .D(reg_z_n235), .CK(clk), .Q(
        round_inst_aout_z[31]) );
  DFF_X1 reg_z_s_current_state_reg_31_ ( .D(reg_z_n234), .CK(clk), .Q(
        round_inst_aout_z[30]) );
  DFF_X1 reg_z_s_current_state_reg_32_ ( .D(reg_z_n233), .CK(clk), .Q(
        round_inst_srout_z[16]) );
  DFF_X1 reg_z_s_current_state_reg_33_ ( .D(reg_z_n232), .CK(clk), .Q(
        round_inst_aout_z[32]) );
  DFF_X1 reg_z_s_current_state_reg_34_ ( .D(reg_z_n231), .CK(clk), .Q(
        round_inst_aout_z[35]) );
  DFF_X1 reg_z_s_current_state_reg_35_ ( .D(reg_z_n230), .CK(clk), .Q(
        round_inst_aout_z[34]) );
  DFF_X1 reg_z_s_current_state_reg_36_ ( .D(reg_z_n229), .CK(clk), .Q(
        round_inst_srout_z[4]) );
  DFF_X1 reg_z_s_current_state_reg_37_ ( .D(reg_z_n228), .CK(clk), .Q(
        round_inst_aout_z[36]) );
  DFF_X1 reg_z_s_current_state_reg_38_ ( .D(reg_z_n227), .CK(clk), .Q(
        round_inst_aout_z[39]) );
  DFF_X1 reg_z_s_current_state_reg_39_ ( .D(reg_z_n226), .CK(clk), .Q(
        round_inst_aout_z[38]) );
  DFF_X1 reg_z_s_current_state_reg_40_ ( .D(reg_z_n225), .CK(clk), .Q(
        round_inst_srout_z[56]) );
  DFF_X1 reg_z_s_current_state_reg_41_ ( .D(reg_z_n224), .CK(clk), .Q(
        round_inst_aout_z[40]) );
  DFF_X1 reg_z_s_current_state_reg_42_ ( .D(reg_z_n223), .CK(clk), .Q(
        round_inst_aout_z[43]) );
  DFF_X1 reg_z_s_current_state_reg_43_ ( .D(reg_z_n222), .CK(clk), .Q(
        round_inst_aout_z[42]) );
  DFF_X1 reg_z_s_current_state_reg_44_ ( .D(reg_z_n221), .CK(clk), .Q(
        round_inst_srout_z[44]) );
  DFF_X1 reg_z_s_current_state_reg_45_ ( .D(reg_z_n220), .CK(clk), .Q(
        round_inst_aout_z[44]) );
  DFF_X1 reg_z_s_current_state_reg_46_ ( .D(reg_z_n219), .CK(clk), .Q(
        round_inst_aout_z[47]) );
  DFF_X1 reg_z_s_current_state_reg_47_ ( .D(reg_z_n218), .CK(clk), .Q(
        round_inst_aout_z[46]) );
  DFF_X1 reg_z_s_current_state_reg_48_ ( .D(reg_z_n217), .CK(clk), .Q(
        round_inst_srout_z[32]) );
  DFF_X1 reg_z_s_current_state_reg_49_ ( .D(reg_z_n216), .CK(clk), .Q(
        round_inst_aout_z[48]) );
  DFF_X1 reg_z_s_current_state_reg_50_ ( .D(reg_z_n215), .CK(clk), .Q(
        round_inst_aout_z[51]) );
  DFF_X1 reg_z_s_current_state_reg_51_ ( .D(reg_z_n214), .CK(clk), .Q(
        round_inst_aout_z[50]) );
  DFF_X1 reg_z_s_current_state_reg_52_ ( .D(reg_z_n213), .CK(clk), .Q(
        round_inst_srout_z[20]) );
  DFF_X1 reg_z_s_current_state_reg_53_ ( .D(reg_z_n212), .CK(clk), .Q(
        round_inst_aout_z[52]) );
  DFF_X1 reg_z_s_current_state_reg_54_ ( .D(reg_z_n211), .CK(clk), .Q(
        round_inst_aout_z[55]) );
  DFF_X1 reg_z_s_current_state_reg_55_ ( .D(reg_z_n210), .CK(clk), .Q(
        round_inst_aout_z[54]) );
  DFF_X1 reg_z_s_current_state_reg_56_ ( .D(reg_z_n209), .CK(clk), .Q(
        round_inst_srout_z[8]) );
  DFF_X1 reg_z_s_current_state_reg_57_ ( .D(reg_z_n208), .CK(clk), .Q(
        round_inst_aout_z[56]) );
  DFF_X1 reg_z_s_current_state_reg_58_ ( .D(reg_z_n207), .CK(clk), .Q(
        round_inst_aout_z[59]) );
  DFF_X1 reg_z_s_current_state_reg_59_ ( .D(reg_z_n206), .CK(clk), .Q(
        round_inst_aout_z[58]) );
  DFF_X1 reg_z_s_current_state_reg_60_ ( .D(reg_z_n205), .CK(clk), .Q(
        round_inst_srout_z[60]) );
  DFF_X1 reg_z_s_current_state_reg_61_ ( .D(reg_z_n204), .CK(clk), .Q(
        round_inst_aout_z[60]) );
  DFF_X1 reg_z_s_current_state_reg_62_ ( .D(reg_z_n203), .CK(clk), .Q(
        round_inst_aout_z[63]) );
  DFF_X1 reg_z_s_current_state_reg_63_ ( .D(reg_z_n202), .CK(clk), .Q(
        round_inst_aout_z[62]) );
  NAND2_X1 reg_b_U17 ( .A1(reg_b_n16), .A2(reg_b_n11), .ZN(reg_b_n15) );
  NAND2_X1 reg_b_U16 ( .A1(bin[3]), .A2(reg_b_n10), .ZN(reg_b_n11) );
  NAND2_X1 reg_b_U15 ( .A1(state_b[3]), .A2(reg_b_n9), .ZN(reg_b_n16) );
  NAND2_X1 reg_b_U14 ( .A1(reg_b_n8), .A2(reg_b_n7), .ZN(reg_b_n14) );
  NAND2_X1 reg_b_U13 ( .A1(bin[2]), .A2(reg_b_n10), .ZN(reg_b_n7) );
  NAND2_X1 reg_b_U12 ( .A1(state_b[2]), .A2(reg_b_n9), .ZN(reg_b_n8) );
  NAND2_X1 reg_b_U11 ( .A1(reg_b_n6), .A2(reg_b_n5), .ZN(reg_b_n13) );
  NAND2_X1 reg_b_U10 ( .A1(bin[1]), .A2(reg_b_n10), .ZN(reg_b_n5) );
  NAND2_X1 reg_b_U9 ( .A1(state_b[1]), .A2(reg_b_n9), .ZN(reg_b_n6) );
  NAND2_X1 reg_b_U8 ( .A1(reg_b_n4), .A2(reg_b_n3), .ZN(reg_b_n12) );
  NAND2_X1 reg_b_U7 ( .A1(reg_b_n9), .A2(state_b[0]), .ZN(reg_b_n3) );
  NOR2_X1 reg_b_U6 ( .A1(rst), .A2(reg_b_n2), .ZN(reg_b_n9) );
  INV_X1 reg_b_U5 ( .A(en_sig), .ZN(reg_b_n2) );
  NAND2_X1 reg_b_U4 ( .A1(reg_b_n10), .A2(bin[0]), .ZN(reg_b_n4) );
  NOR2_X1 reg_b_U3 ( .A1(en_sig), .A2(rst), .ZN(reg_b_n10) );
  DFF_X1 reg_b_s_current_state_reg_0_ ( .D(reg_b_n12), .CK(clk), .Q(bin[0]) );
  DFF_X1 reg_b_s_current_state_reg_1_ ( .D(reg_b_n13), .CK(clk), .Q(bin[1]) );
  DFF_X1 reg_b_s_current_state_reg_2_ ( .D(reg_b_n14), .CK(clk), .Q(bin[2]) );
  DFF_X1 reg_b_s_current_state_reg_3_ ( .D(reg_b_n15), .CK(clk), .Q(bin[3]) );
  NAND2_X1 reg_c_U17 ( .A1(reg_c_n40), .A2(reg_c_n39), .ZN(reg_c_n17) );
  NAND2_X1 reg_c_U16 ( .A1(cin[2]), .A2(reg_c_n38), .ZN(reg_c_n39) );
  NAND2_X1 reg_c_U15 ( .A1(state_c[2]), .A2(reg_c_n37), .ZN(reg_c_n40) );
  NAND2_X1 reg_c_U14 ( .A1(reg_c_n36), .A2(reg_c_n35), .ZN(reg_c_n18) );
  NAND2_X1 reg_c_U13 ( .A1(cin[1]), .A2(reg_c_n38), .ZN(reg_c_n35) );
  NAND2_X1 reg_c_U12 ( .A1(state_c[1]), .A2(reg_c_n37), .ZN(reg_c_n36) );
  NAND2_X1 reg_c_U11 ( .A1(reg_c_n34), .A2(reg_c_n33), .ZN(reg_c_n19) );
  NAND2_X1 reg_c_U10 ( .A1(cin[0]), .A2(reg_c_n38), .ZN(reg_c_n33) );
  NAND2_X1 reg_c_U9 ( .A1(state_c[0]), .A2(reg_c_n37), .ZN(reg_c_n34) );
  NAND2_X1 reg_c_U8 ( .A1(reg_c_n32), .A2(reg_c_n31), .ZN(reg_c_n16) );
  NAND2_X1 reg_c_U7 ( .A1(reg_c_n37), .A2(state_c[3]), .ZN(reg_c_n31) );
  NOR2_X1 reg_c_U6 ( .A1(rst), .A2(reg_c_n30), .ZN(reg_c_n37) );
  INV_X1 reg_c_U5 ( .A(en_sig), .ZN(reg_c_n30) );
  NAND2_X1 reg_c_U4 ( .A1(reg_c_n38), .A2(cin[3]), .ZN(reg_c_n32) );
  NOR2_X1 reg_c_U3 ( .A1(en_sig), .A2(rst), .ZN(reg_c_n38) );
  DFF_X1 reg_c_s_current_state_reg_0_ ( .D(reg_c_n19), .CK(clk), .Q(cin[0]) );
  DFF_X1 reg_c_s_current_state_reg_1_ ( .D(reg_c_n18), .CK(clk), .Q(cin[1]) );
  DFF_X1 reg_c_s_current_state_reg_2_ ( .D(reg_c_n17), .CK(clk), .Q(cin[2]) );
  DFF_X1 reg_c_s_current_state_reg_3_ ( .D(reg_c_n16), .CK(clk), .Q(cin[3]) );
  NAND2_X1 reg_d_U17 ( .A1(reg_d_n40), .A2(reg_d_n39), .ZN(reg_d_n16) );
  NAND2_X1 reg_d_U16 ( .A1(din[3]), .A2(reg_d_n38), .ZN(reg_d_n39) );
  NAND2_X1 reg_d_U15 ( .A1(state_d[3]), .A2(reg_d_n37), .ZN(reg_d_n40) );
  NAND2_X1 reg_d_U14 ( .A1(reg_d_n36), .A2(reg_d_n35), .ZN(reg_d_n17) );
  NAND2_X1 reg_d_U13 ( .A1(din[2]), .A2(reg_d_n38), .ZN(reg_d_n35) );
  NAND2_X1 reg_d_U12 ( .A1(state_d[2]), .A2(reg_d_n37), .ZN(reg_d_n36) );
  NAND2_X1 reg_d_U11 ( .A1(reg_d_n34), .A2(reg_d_n33), .ZN(reg_d_n18) );
  NAND2_X1 reg_d_U10 ( .A1(din[1]), .A2(reg_d_n38), .ZN(reg_d_n33) );
  NAND2_X1 reg_d_U9 ( .A1(state_d[1]), .A2(reg_d_n37), .ZN(reg_d_n34) );
  NAND2_X1 reg_d_U8 ( .A1(reg_d_n32), .A2(reg_d_n31), .ZN(reg_d_n19) );
  NAND2_X1 reg_d_U7 ( .A1(reg_d_n37), .A2(state_d[0]), .ZN(reg_d_n31) );
  NOR2_X1 reg_d_U6 ( .A1(rst), .A2(reg_d_n30), .ZN(reg_d_n37) );
  INV_X1 reg_d_U5 ( .A(en_sig), .ZN(reg_d_n30) );
  NAND2_X1 reg_d_U4 ( .A1(reg_d_n38), .A2(din[0]), .ZN(reg_d_n32) );
  NOR2_X1 reg_d_U3 ( .A1(en_sig), .A2(rst), .ZN(reg_d_n38) );
  DFF_X1 reg_d_s_current_state_reg_0_ ( .D(reg_d_n19), .CK(clk), .Q(din[0]) );
  DFF_X1 reg_d_s_current_state_reg_1_ ( .D(reg_d_n18), .CK(clk), .Q(din[1]) );
  DFF_X1 reg_d_s_current_state_reg_2_ ( .D(reg_d_n17), .CK(clk), .Q(din[2]) );
  DFF_X1 reg_d_s_current_state_reg_3_ ( .D(reg_d_n16), .CK(clk), .Q(din[3]) );
  NAND2_X1 cntrl_inst_U183 ( .A1(cntrl_inst_n218), .A2(cntrl_inst_n217), .ZN(
        cntrl_inst_n102) );
  NAND3_X1 cntrl_inst_U182 ( .A1(cntrl_inst_n206), .A2(cntrl_inst_counter[0]), 
        .A3(cntrl_inst_n216), .ZN(cntrl_inst_n218) );
  MUX2_X1 cntrl_inst_U181 ( .A(cntrl_inst_n215), .B(cntrl_inst_n214), .S(
        cntrl_inst_n219), .Z(cntrl_inst_n98) );
  NOR2_X1 cntrl_inst_U180 ( .A1(cntrl_inst_n216), .A2(cntrl_inst_n221), .ZN(
        cntrl_inst_n214) );
  NAND2_X1 cntrl_inst_U179 ( .A1(cntrl_inst_n217), .A2(cntrl_inst_n213), .ZN(
        cntrl_inst_n215) );
  NAND2_X1 cntrl_inst_U178 ( .A1(cntrl_inst_n206), .A2(cntrl_inst_n216), .ZN(
        cntrl_inst_n213) );
  NAND2_X1 cntrl_inst_U177 ( .A1(cntrl_inst_n212), .A2(cntrl_inst_n221), .ZN(
        cntrl_inst_n217) );
  INV_X1 cntrl_inst_U176 ( .A(cntrl_inst_n216), .ZN(cntrl_inst_n212) );
  MUX2_X1 cntrl_inst_U175 ( .A(cntrl_inst_n211), .B(cntrl_inst_n210), .S(
        cntrl_inst_n220), .Z(cntrl_inst_n99) );
  MUX2_X1 cntrl_inst_U174 ( .A(cntrl_inst_n209), .B(cntrl_inst_n206), .S(
        cntrl_inst_n216), .Z(cntrl_inst_n211) );
  NAND2_X1 cntrl_inst_U173 ( .A1(cntrl_inst_counter[0]), .A2(
        cntrl_inst_counter[1]), .ZN(cntrl_inst_n209) );
  NAND2_X1 cntrl_inst_U172 ( .A1(cntrl_inst_n208), .A2(cntrl_inst_n207), .ZN(
        cntrl_inst_n100) );
  NAND2_X1 cntrl_inst_U171 ( .A1(cntrl_inst_n206), .A2(cntrl_inst_n222), .ZN(
        cntrl_inst_n207) );
  NAND2_X1 cntrl_inst_U170 ( .A1(cntrl_inst_counter[2]), .A2(cntrl_inst_n210), 
        .ZN(cntrl_inst_n208) );
  NOR3_X1 cntrl_inst_U169 ( .A1(cntrl_inst_n219), .A2(cntrl_inst_n221), .A3(
        cntrl_inst_n216), .ZN(cntrl_inst_n210) );
  NAND3_X1 cntrl_inst_U168 ( .A1(cntrl_inst_n206), .A2(cntrl_inst_n205), .A3(
        en), .ZN(cntrl_inst_n216) );
  OR3_X1 cntrl_inst_U167 ( .A1(cntrl_inst_n204), .A2(cntrl_inst_n220), .A3(
        inv_sig), .ZN(cntrl_inst_n205) );
  NOR2_X1 cntrl_inst_U166 ( .A1(cntrl_inst_counter[1]), .A2(
        cntrl_inst_counter[0]), .ZN(cntrl_inst_n204) );
  INV_X1 cntrl_inst_U165 ( .A(rst), .ZN(cntrl_inst_n206) );
  XOR2_X1 cntrl_inst_U164 ( .A(k[56]), .B(cntrl_inst_n203), .Z(rc_56_) );
  XOR2_X1 cntrl_inst_U163 ( .A(k[44]), .B(cntrl_inst_n202), .Z(rc_44_) );
  XNOR2_X1 cntrl_inst_U162 ( .A(cntrl_inst_n201), .B(k[28]), .ZN(rc_28_) );
  XOR2_X1 cntrl_inst_U161 ( .A(k[9]), .B(cntrl_inst_n203), .Z(rc_9_) );
  NAND3_X1 cntrl_inst_U160 ( .A1(cntrl_inst_n200), .A2(cntrl_inst_n199), .A3(
        cntrl_inst_n198), .ZN(cntrl_inst_n203) );
  XOR2_X1 cntrl_inst_U159 ( .A(k[17]), .B(cntrl_inst_n202), .Z(rc_17_) );
  XNOR2_X1 cntrl_inst_U158 ( .A(cntrl_inst_n201), .B(k[5]), .ZN(rc_5_) );
  XOR2_X1 cntrl_inst_U157 ( .A(k[58]), .B(cntrl_inst_n197), .Z(rc_58_) );
  XNOR2_X1 cntrl_inst_U156 ( .A(cntrl_inst_n196), .B(k[26]), .ZN(rc_26_) );
  XNOR2_X1 cntrl_inst_U155 ( .A(cntrl_inst_n201), .B(k[38]), .ZN(rc_38_) );
  XNOR2_X1 cntrl_inst_U154 ( .A(cntrl_inst_n196), .B(k[10]), .ZN(rc_10_) );
  XNOR2_X1 cntrl_inst_U153 ( .A(cntrl_inst_n196), .B(k[46]), .ZN(rc_46_) );
  XNOR2_X1 cntrl_inst_U152 ( .A(cntrl_inst_n196), .B(k[11]), .ZN(rc_11_) );
  XNOR2_X1 cntrl_inst_U151 ( .A(cntrl_inst_n196), .B(k[59]), .ZN(rc_59_) );
  XOR2_X1 cntrl_inst_U150 ( .A(k[23]), .B(cntrl_inst_n197), .Z(rc_23_) );
  NAND2_X1 cntrl_inst_U149 ( .A1(cntrl_inst_n195), .A2(cntrl_inst_n201), .ZN(
        cntrl_inst_n197) );
  NOR2_X1 cntrl_inst_U148 ( .A1(cntrl_inst_n194), .A2(cntrl_inst_n193), .ZN(
        cntrl_inst_n201) );
  XOR2_X1 cntrl_inst_U147 ( .A(k[0]), .B(cntrl_inst_n192), .Z(rc_0_) );
  XNOR2_X1 cntrl_inst_U146 ( .A(cntrl_inst_n191), .B(k[12]), .ZN(rc_12_) );
  XNOR2_X1 cntrl_inst_U145 ( .A(k[13]), .B(cntrl_inst_n190), .ZN(rc_13_) );
  NOR2_X1 cntrl_inst_U144 ( .A1(cntrl_inst_n189), .A2(cntrl_inst_n202), .ZN(
        cntrl_inst_n190) );
  NAND2_X1 cntrl_inst_U143 ( .A1(cntrl_inst_n195), .A2(cntrl_inst_n188), .ZN(
        cntrl_inst_n202) );
  XNOR2_X1 cntrl_inst_U142 ( .A(k[14]), .B(cntrl_inst_n187), .ZN(rc_14_) );
  NOR3_X1 cntrl_inst_U141 ( .A1(cntrl_inst_n186), .A2(cntrl_inst_n185), .A3(
        cntrl_inst_n184), .ZN(cntrl_inst_n187) );
  XOR2_X1 cntrl_inst_U140 ( .A(k[16]), .B(cntrl_inst_n183), .Z(rc_16_) );
  XOR2_X1 cntrl_inst_U139 ( .A(k[18]), .B(cntrl_inst_n182), .Z(rc_18_) );
  XNOR2_X1 cntrl_inst_U138 ( .A(k[19]), .B(cntrl_inst_n181), .ZN(rc_19_) );
  NOR3_X1 cntrl_inst_U137 ( .A1(cntrl_inst_n180), .A2(cntrl_inst_n179), .A3(
        cntrl_inst_n178), .ZN(cntrl_inst_n181) );
  NAND2_X1 cntrl_inst_U136 ( .A1(cntrl_inst_n177), .A2(cntrl_inst_n198), .ZN(
        cntrl_inst_n178) );
  XOR2_X1 cntrl_inst_U135 ( .A(k[1]), .B(cntrl_inst_n194), .Z(rc_1_) );
  NAND2_X1 cntrl_inst_U134 ( .A1(cntrl_inst_n199), .A2(cntrl_inst_n198), .ZN(
        cntrl_inst_n194) );
  XNOR2_X1 cntrl_inst_U133 ( .A(cntrl_inst_n191), .B(k[20]), .ZN(rc_20_) );
  XNOR2_X1 cntrl_inst_U132 ( .A(cntrl_inst_n176), .B(k[21]), .ZN(rc_21_) );
  NOR2_X1 cntrl_inst_U131 ( .A1(cntrl_inst_n175), .A2(cntrl_inst_n185), .ZN(
        cntrl_inst_n176) );
  XNOR2_X1 cntrl_inst_U130 ( .A(k[22]), .B(cntrl_inst_n174), .ZN(rc_22_) );
  NOR3_X1 cntrl_inst_U129 ( .A1(cntrl_inst_n173), .A2(cntrl_inst_n172), .A3(
        cntrl_inst_n184), .ZN(cntrl_inst_n174) );
  NAND2_X1 cntrl_inst_U128 ( .A1(cntrl_inst_n171), .A2(cntrl_inst_n170), .ZN(
        cntrl_inst_n184) );
  NAND2_X1 cntrl_inst_U127 ( .A1(cntrl_inst_n169), .A2(cntrl_inst_n168), .ZN(
        cntrl_inst_n170) );
  XOR2_X1 cntrl_inst_U126 ( .A(k[24]), .B(cntrl_inst_n167), .Z(rc_24_) );
  NAND2_X1 cntrl_inst_U125 ( .A1(cntrl_inst_n198), .A2(cntrl_inst_n166), .ZN(
        cntrl_inst_n167) );
  NOR2_X1 cntrl_inst_U124 ( .A1(cntrl_inst_n165), .A2(cntrl_inst_n164), .ZN(
        cntrl_inst_n166) );
  XOR2_X1 cntrl_inst_U123 ( .A(cntrl_inst_n189), .B(k[25]), .Z(rc_25_) );
  XOR2_X1 cntrl_inst_U122 ( .A(k[27]), .B(cntrl_inst_n163), .Z(rc_27_) );
  NAND2_X1 cntrl_inst_U121 ( .A1(cntrl_inst_n162), .A2(cntrl_inst_n161), .ZN(
        cntrl_inst_n163) );
  XOR2_X1 cntrl_inst_U120 ( .A(k[29]), .B(cntrl_inst_n160), .Z(rc_29_) );
  NAND2_X1 cntrl_inst_U119 ( .A1(cntrl_inst_n159), .A2(cntrl_inst_n158), .ZN(
        cntrl_inst_n160) );
  XNOR2_X1 cntrl_inst_U118 ( .A(cntrl_inst_n157), .B(k[2]), .ZN(rc_2_) );
  XOR2_X1 cntrl_inst_U117 ( .A(k[30]), .B(cntrl_inst_n156), .Z(rc_30_) );
  XOR2_X1 cntrl_inst_U116 ( .A(k[31]), .B(cntrl_inst_n156), .Z(rc_31_) );
  XOR2_X1 cntrl_inst_U115 ( .A(k[32]), .B(cntrl_inst_n155), .Z(rc_32_) );
  NAND3_X1 cntrl_inst_U114 ( .A1(cntrl_inst_n154), .A2(cntrl_inst_n153), .A3(
        cntrl_inst_n152), .ZN(cntrl_inst_n155) );
  XNOR2_X1 cntrl_inst_U113 ( .A(cntrl_inst_n151), .B(k[33]), .ZN(rc_33_) );
  XNOR2_X1 cntrl_inst_U112 ( .A(cntrl_inst_n157), .B(k[34]), .ZN(rc_34_) );
  NOR2_X1 cntrl_inst_U111 ( .A1(cntrl_inst_n175), .A2(cntrl_inst_n172), .ZN(
        cntrl_inst_n157) );
  XOR2_X1 cntrl_inst_U110 ( .A(k[35]), .B(cntrl_inst_n150), .Z(rc_35_) );
  XOR2_X1 cntrl_inst_U109 ( .A(k[36]), .B(cntrl_inst_n156), .Z(rc_36_) );
  NAND2_X1 cntrl_inst_U108 ( .A1(cntrl_inst_n161), .A2(cntrl_inst_n152), .ZN(
        cntrl_inst_n156) );
  XNOR2_X1 cntrl_inst_U107 ( .A(cntrl_inst_n191), .B(k[37]), .ZN(rc_37_) );
  NOR3_X1 cntrl_inst_U106 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n165), .A3(
        cntrl_inst_n164), .ZN(cntrl_inst_n191) );
  XNOR2_X1 cntrl_inst_U105 ( .A(k[39]), .B(cntrl_inst_n148), .ZN(rc_39_) );
  NOR3_X1 cntrl_inst_U104 ( .A1(cntrl_inst_n180), .A2(cntrl_inst_n179), .A3(
        cntrl_inst_n172), .ZN(cntrl_inst_n148) );
  XNOR2_X1 cntrl_inst_U103 ( .A(cntrl_inst_n147), .B(k[3]), .ZN(rc_3_) );
  XNOR2_X1 cntrl_inst_U102 ( .A(cntrl_inst_n146), .B(k[40]), .ZN(rc_40_) );
  XOR2_X1 cntrl_inst_U101 ( .A(k[41]), .B(cntrl_inst_n150), .Z(rc_41_) );
  NAND2_X1 cntrl_inst_U100 ( .A1(cntrl_inst_n200), .A2(cntrl_inst_n196), .ZN(
        cntrl_inst_n150) );
  NOR2_X1 cntrl_inst_U99 ( .A1(cntrl_inst_n180), .A2(cntrl_inst_n165), .ZN(
        cntrl_inst_n196) );
  XOR2_X1 cntrl_inst_U98 ( .A(cntrl_inst_n193), .B(k[42]), .Z(rc_42_) );
  XOR2_X1 cntrl_inst_U97 ( .A(k[43]), .B(cntrl_inst_n145), .Z(rc_43_) );
  NAND2_X1 cntrl_inst_U96 ( .A1(cntrl_inst_n198), .A2(cntrl_inst_n144), .ZN(
        cntrl_inst_n145) );
  XOR2_X1 cntrl_inst_U95 ( .A(k[45]), .B(cntrl_inst_n143), .Z(rc_45_) );
  NAND2_X1 cntrl_inst_U94 ( .A1(cntrl_inst_n153), .A2(cntrl_inst_n158), .ZN(
        cntrl_inst_n143) );
  XOR2_X1 cntrl_inst_U93 ( .A(k[47]), .B(cntrl_inst_n142), .Z(rc_47_) );
  NAND2_X1 cntrl_inst_U92 ( .A1(cntrl_inst_n200), .A2(cntrl_inst_n188), .ZN(
        cntrl_inst_n142) );
  INV_X1 cntrl_inst_U91 ( .A(cntrl_inst_n189), .ZN(cntrl_inst_n200) );
  XOR2_X1 cntrl_inst_U90 ( .A(k[48]), .B(cntrl_inst_n141), .Z(rc_48_) );
  NAND2_X1 cntrl_inst_U89 ( .A1(cntrl_inst_n140), .A2(cntrl_inst_n139), .ZN(
        cntrl_inst_n141) );
  NAND2_X1 cntrl_inst_U88 ( .A1(cntrl_inst_n138), .A2(cntrl_inst_n169), .ZN(
        cntrl_inst_n140) );
  XNOR2_X1 cntrl_inst_U87 ( .A(cntrl_inst_n188), .B(k[49]), .ZN(rc_49_) );
  NOR2_X1 cntrl_inst_U86 ( .A1(cntrl_inst_n137), .A2(cntrl_inst_n136), .ZN(
        cntrl_inst_n188) );
  INV_X1 cntrl_inst_U85 ( .A(cntrl_inst_n135), .ZN(cntrl_inst_n137) );
  XNOR2_X1 cntrl_inst_U84 ( .A(k[4]), .B(cntrl_inst_n134), .ZN(rc_4_) );
  NOR3_X1 cntrl_inst_U83 ( .A1(cntrl_inst_n133), .A2(cntrl_inst_n165), .A3(
        cntrl_inst_n179), .ZN(cntrl_inst_n134) );
  XNOR2_X1 cntrl_inst_U82 ( .A(cntrl_inst_n147), .B(k[50]), .ZN(rc_50_) );
  NOR3_X1 cntrl_inst_U81 ( .A1(cntrl_inst_n180), .A2(cntrl_inst_n179), .A3(
        cntrl_inst_n185), .ZN(cntrl_inst_n147) );
  XOR2_X1 cntrl_inst_U80 ( .A(k[51]), .B(cntrl_inst_n132), .Z(rc_51_) );
  NAND2_X1 cntrl_inst_U79 ( .A1(cntrl_inst_n144), .A2(cntrl_inst_n199), .ZN(
        cntrl_inst_n132) );
  INV_X1 cntrl_inst_U78 ( .A(cntrl_inst_n149), .ZN(cntrl_inst_n199) );
  NOR2_X1 cntrl_inst_U77 ( .A1(cntrl_inst_n131), .A2(cntrl_inst_n164), .ZN(
        cntrl_inst_n144) );
  NAND2_X1 cntrl_inst_U76 ( .A1(cntrl_inst_n130), .A2(cntrl_inst_n177), .ZN(
        cntrl_inst_n164) );
  XNOR2_X1 cntrl_inst_U75 ( .A(cntrl_inst_n129), .B(k[52]), .ZN(rc_52_) );
  XOR2_X1 cntrl_inst_U74 ( .A(k[53]), .B(cntrl_inst_n192), .Z(rc_53_) );
  NAND2_X1 cntrl_inst_U73 ( .A1(cntrl_inst_n161), .A2(cntrl_inst_n128), .ZN(
        cntrl_inst_n192) );
  XOR2_X1 cntrl_inst_U72 ( .A(cntrl_inst_n193), .B(k[54]), .Z(rc_54_) );
  XOR2_X1 cntrl_inst_U71 ( .A(k[55]), .B(cntrl_inst_n127), .Z(rc_55_) );
  NAND2_X1 cntrl_inst_U70 ( .A1(cntrl_inst_n153), .A2(cntrl_inst_n159), .ZN(
        cntrl_inst_n127) );
  XNOR2_X1 cntrl_inst_U69 ( .A(cntrl_inst_n129), .B(k[57]), .ZN(rc_57_) );
  XNOR2_X1 cntrl_inst_U68 ( .A(cntrl_inst_n129), .B(k[60]), .ZN(rc_60_) );
  NOR2_X1 cntrl_inst_U67 ( .A1(cntrl_inst_n189), .A2(cntrl_inst_n193), .ZN(
        cntrl_inst_n129) );
  INV_X1 cntrl_inst_U66 ( .A(cntrl_inst_n126), .ZN(cntrl_inst_n193) );
  XOR2_X1 cntrl_inst_U65 ( .A(k[61]), .B(cntrl_inst_n183), .Z(rc_61_) );
  NAND2_X1 cntrl_inst_U64 ( .A1(cntrl_inst_n195), .A2(cntrl_inst_n126), .ZN(
        cntrl_inst_n183) );
  NOR2_X1 cntrl_inst_U63 ( .A1(cntrl_inst_n186), .A2(cntrl_inst_n173), .ZN(
        cntrl_inst_n126) );
  INV_X1 cntrl_inst_U62 ( .A(cntrl_inst_n125), .ZN(cntrl_inst_n186) );
  NOR2_X1 cntrl_inst_U61 ( .A1(cntrl_inst_n124), .A2(cntrl_inst_n123), .ZN(
        cntrl_inst_n195) );
  XNOR2_X1 cntrl_inst_U60 ( .A(cntrl_inst_n146), .B(k[62]), .ZN(rc_62_) );
  NOR3_X1 cntrl_inst_U59 ( .A1(cntrl_inst_n165), .A2(cntrl_inst_n179), .A3(
        cntrl_inst_n172), .ZN(cntrl_inst_n146) );
  INV_X1 cntrl_inst_U58 ( .A(cntrl_inst_n128), .ZN(cntrl_inst_n172) );
  NOR2_X1 cntrl_inst_U57 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n123), .ZN(
        cntrl_inst_n128) );
  NOR2_X1 cntrl_inst_U56 ( .A1(cntrl_inst_n122), .A2(cntrl_inst_n152), .ZN(
        cntrl_inst_n123) );
  INV_X1 cntrl_inst_U55 ( .A(cntrl_inst_n185), .ZN(cntrl_inst_n152) );
  NOR2_X1 cntrl_inst_U54 ( .A1(cntrl_inst_n162), .A2(cntrl_inst_n122), .ZN(
        cntrl_inst_n149) );
  XOR2_X1 cntrl_inst_U53 ( .A(k[63]), .B(cntrl_inst_n121), .Z(rc_63_) );
  NAND4_X1 cntrl_inst_U52 ( .A1(cntrl_inst_n154), .A2(cntrl_inst_n177), .A3(
        cntrl_inst_n153), .A4(cntrl_inst_n198), .ZN(cntrl_inst_n121) );
  XNOR2_X1 cntrl_inst_U51 ( .A(cntrl_inst_n151), .B(k[6]), .ZN(rc_6_) );
  NOR2_X1 cntrl_inst_U50 ( .A1(cntrl_inst_n133), .A2(cntrl_inst_n175), .ZN(
        cntrl_inst_n151) );
  NAND2_X1 cntrl_inst_U49 ( .A1(cntrl_inst_n130), .A2(cntrl_inst_n154), .ZN(
        cntrl_inst_n175) );
  NOR2_X1 cntrl_inst_U48 ( .A1(cntrl_inst_n136), .A2(cntrl_inst_n173), .ZN(
        cntrl_inst_n154) );
  NOR2_X1 cntrl_inst_U47 ( .A1(cntrl_inst_n158), .A2(cntrl_inst_n120), .ZN(
        cntrl_inst_n173) );
  INV_X1 cntrl_inst_U46 ( .A(cntrl_inst_n119), .ZN(cntrl_inst_n120) );
  AND2_X1 cntrl_inst_U45 ( .A1(cntrl_inst_n118), .A2(cntrl_inst_n165), .ZN(
        cntrl_inst_n136) );
  NOR2_X1 cntrl_inst_U44 ( .A1(cntrl_inst_n117), .A2(cntrl_inst_n116), .ZN(
        cntrl_inst_n130) );
  NOR2_X1 cntrl_inst_U43 ( .A1(cntrl_inst_n138), .A2(cntrl_inst_n153), .ZN(
        cntrl_inst_n116) );
  XOR2_X1 cntrl_inst_U42 ( .A(k[7]), .B(cntrl_inst_n182), .Z(rc_7_) );
  NAND3_X1 cntrl_inst_U41 ( .A1(cntrl_inst_n161), .A2(cntrl_inst_n177), .A3(
        cntrl_inst_n198), .ZN(cntrl_inst_n182) );
  NAND2_X1 cntrl_inst_U40 ( .A1(cntrl_inst_n122), .A2(cntrl_inst_n185), .ZN(
        cntrl_inst_n198) );
  INV_X1 cntrl_inst_U39 ( .A(cntrl_inst_n124), .ZN(cntrl_inst_n177) );
  NOR2_X1 cntrl_inst_U38 ( .A1(cntrl_inst_n118), .A2(cntrl_inst_n162), .ZN(
        cntrl_inst_n124) );
  INV_X1 cntrl_inst_U37 ( .A(cntrl_inst_n133), .ZN(cntrl_inst_n162) );
  NOR2_X1 cntrl_inst_U36 ( .A1(cntrl_inst_n179), .A2(cntrl_inst_n131), .ZN(
        cntrl_inst_n161) );
  NAND2_X1 cntrl_inst_U35 ( .A1(cntrl_inst_n135), .A2(cntrl_inst_n125), .ZN(
        cntrl_inst_n131) );
  NAND2_X1 cntrl_inst_U34 ( .A1(cntrl_inst_n122), .A2(cntrl_inst_n165), .ZN(
        cntrl_inst_n125) );
  NOR2_X1 cntrl_inst_U33 ( .A1(cntrl_inst_n168), .A2(cntrl_inst_n159), .ZN(
        cntrl_inst_n165) );
  NAND2_X1 cntrl_inst_U32 ( .A1(cntrl_inst_n122), .A2(cntrl_inst_n180), .ZN(
        cntrl_inst_n135) );
  NOR2_X1 cntrl_inst_U31 ( .A1(cntrl_inst_n138), .A2(cntrl_inst_n158), .ZN(
        cntrl_inst_n180) );
  XNOR2_X1 cntrl_inst_U30 ( .A(k[8]), .B(cntrl_inst_n115), .ZN(rc_8_) );
  NOR3_X1 cntrl_inst_U29 ( .A1(cntrl_inst_n133), .A2(cntrl_inst_n185), .A3(
        cntrl_inst_n189), .ZN(cntrl_inst_n115) );
  NAND2_X1 cntrl_inst_U28 ( .A1(cntrl_inst_n171), .A2(cntrl_inst_n114), .ZN(
        cntrl_inst_n189) );
  NAND2_X1 cntrl_inst_U27 ( .A1(cntrl_inst_n138), .A2(cntrl_inst_n179), .ZN(
        cntrl_inst_n114) );
  INV_X1 cntrl_inst_U26 ( .A(cntrl_inst_n153), .ZN(cntrl_inst_n179) );
  NAND2_X1 cntrl_inst_U25 ( .A1(cntrl_inst_n113), .A2(cntrl_inst_n169), .ZN(
        cntrl_inst_n153) );
  NOR2_X1 cntrl_inst_U24 ( .A1(cntrl_inst_n112), .A2(cntrl_inst_n118), .ZN(
        cntrl_inst_n169) );
  INV_X1 cntrl_inst_U23 ( .A(cntrl_inst_n117), .ZN(cntrl_inst_n171) );
  NOR2_X1 cntrl_inst_U22 ( .A1(cntrl_inst_n113), .A2(cntrl_inst_n139), .ZN(
        cntrl_inst_n117) );
  NAND2_X1 cntrl_inst_U21 ( .A1(cntrl_inst_n112), .A2(cntrl_inst_n119), .ZN(
        cntrl_inst_n139) );
  NOR2_X1 cntrl_inst_U20 ( .A1(cntrl_inst_n122), .A2(cntrl_inst_n138), .ZN(
        cntrl_inst_n119) );
  INV_X1 cntrl_inst_U19 ( .A(cntrl_inst_n118), .ZN(cntrl_inst_n122) );
  XOR2_X1 cntrl_inst_U18 ( .A(cntrl_inst_n219), .B(enc), .Z(cntrl_inst_n118)
         );
  NOR2_X1 cntrl_inst_U17 ( .A1(cntrl_inst_n138), .A2(cntrl_inst_n159), .ZN(
        cntrl_inst_n185) );
  NAND2_X1 cntrl_inst_U16 ( .A1(cntrl_inst_n112), .A2(cntrl_inst_n113), .ZN(
        cntrl_inst_n159) );
  INV_X1 cntrl_inst_U15 ( .A(cntrl_inst_n168), .ZN(cntrl_inst_n138) );
  NOR2_X1 cntrl_inst_U14 ( .A1(cntrl_inst_n168), .A2(cntrl_inst_n158), .ZN(
        cntrl_inst_n133) );
  OR2_X1 cntrl_inst_U13 ( .A1(cntrl_inst_n112), .A2(cntrl_inst_n113), .ZN(
        cntrl_inst_n158) );
  XNOR2_X1 cntrl_inst_U12 ( .A(enc), .B(cntrl_inst_n222), .ZN(cntrl_inst_n113)
         );
  XNOR2_X1 cntrl_inst_U11 ( .A(enc), .B(cntrl_inst_n220), .ZN(cntrl_inst_n112)
         );
  XOR2_X1 cntrl_inst_U10 ( .A(enc), .B(cntrl_inst_n221), .Z(cntrl_inst_n168)
         );
  INV_X1 cntrl_inst_U9 ( .A(cntrl_inst_n110), .ZN(done) );
  INV_X1 cntrl_inst_U8 ( .A(cntrl_inst_n108), .ZN(start_sig) );
  OR3_X1 cntrl_inst_U7 ( .A1(inv_sig), .A2(cntrl_inst_n220), .A3(
        cntrl_inst_n109), .ZN(cntrl_inst_n110) );
  NAND2_X1 cntrl_inst_U6 ( .A1(cntrl_inst_counter[0]), .A2(cntrl_inst_n219), 
        .ZN(cntrl_inst_n109) );
  NOR2_X2 cntrl_inst_U5 ( .A1(done), .A2(cntrl_inst_n111), .ZN(en_sig) );
  INV_X1 cntrl_inst_U4 ( .A(en), .ZN(cntrl_inst_n111) );
  OR4_X1 cntrl_inst_U3 ( .A1(cntrl_inst_counter[2]), .A2(cntrl_inst_n222), 
        .A3(cntrl_inst_n111), .A4(cntrl_inst_n109), .ZN(cntrl_inst_n108) );
  DFF_X1 cntrl_inst_counter_reg_3_ ( .D(cntrl_inst_n100), .CK(clk), .Q(
        cntrl_inst_n222), .QN(inv_sig) );
  DFF_X1 cntrl_inst_counter_reg_2_ ( .D(cntrl_inst_n99), .CK(clk), .Q(
        cntrl_inst_counter[2]), .QN(cntrl_inst_n220) );
  DFF_X1 cntrl_inst_counter_reg_1_ ( .D(cntrl_inst_n98), .CK(clk), .Q(
        cntrl_inst_counter[1]), .QN(cntrl_inst_n219) );
  DFF_X1 cntrl_inst_counter_reg_0_ ( .D(cntrl_inst_n102), .CK(clk), .Q(
        cntrl_inst_counter[0]), .QN(cntrl_inst_n221) );
  XOR2_X1 round_inst_U194 ( .A(rc_0_), .B(round_inst_xin_w[0]), .Z(
        round_inst_srout2_w[16]) );
  XOR2_X1 round_inst_U193 ( .A(rc_10_), .B(round_inst_xin_w[10]), .Z(
        round_inst_srout2_w[58]) );
  XOR2_X1 round_inst_U192 ( .A(rc_11_), .B(round_inst_xin_w[11]), .Z(
        round_inst_srout2_w[59]) );
  XOR2_X1 round_inst_U191 ( .A(rc_12_), .B(round_inst_xin_w[12]), .Z(
        round_inst_srout2_w[12]) );
  XOR2_X1 round_inst_U190 ( .A(rc_13_), .B(round_inst_xin_w[13]), .Z(
        round_inst_srout2_w[13]) );
  XOR2_X1 round_inst_U189 ( .A(rc_14_), .B(round_inst_xin_w[14]), .Z(
        round_inst_srout2_w[14]) );
  XOR2_X1 round_inst_U188 ( .A(k[15]), .B(round_inst_xin_w[15]), .Z(
        round_inst_srout2_w[15]) );
  XOR2_X1 round_inst_U187 ( .A(rc_16_), .B(round_inst_xin_w[16]), .Z(
        round_inst_srout2_w[32]) );
  XOR2_X1 round_inst_U186 ( .A(rc_17_), .B(round_inst_xin_w[17]), .Z(
        round_inst_srout2_w[33]) );
  XOR2_X1 round_inst_U185 ( .A(rc_18_), .B(round_inst_xin_w[18]), .Z(
        round_inst_srout2_w[34]) );
  XOR2_X1 round_inst_U184 ( .A(rc_19_), .B(round_inst_xin_w[19]), .Z(
        round_inst_srout2_w[35]) );
  XOR2_X1 round_inst_U183 ( .A(rc_1_), .B(round_inst_xin_w[1]), .Z(
        round_inst_srout2_w[17]) );
  XOR2_X1 round_inst_U182 ( .A(rc_20_), .B(round_inst_xin_w[20]), .Z(
        round_inst_srout2_w[52]) );
  XOR2_X1 round_inst_U181 ( .A(rc_21_), .B(round_inst_xin_w[21]), .Z(
        round_inst_srout2_w[53]) );
  XOR2_X1 round_inst_U180 ( .A(rc_22_), .B(round_inst_xin_w[22]), .Z(
        round_inst_srout2_w[54]) );
  XOR2_X1 round_inst_U179 ( .A(rc_23_), .B(round_inst_xin_w[23]), .Z(
        round_inst_srout2_w[55]) );
  XOR2_X1 round_inst_U178 ( .A(rc_24_), .B(round_inst_xin_w[24]), .Z(
        round_inst_srout2_w[8]) );
  XOR2_X1 round_inst_U177 ( .A(rc_25_), .B(round_inst_xin_w[25]), .Z(
        round_inst_srout2_w[9]) );
  XOR2_X1 round_inst_U176 ( .A(rc_26_), .B(round_inst_xin_w[26]), .Z(
        round_inst_srout2_w[10]) );
  XOR2_X1 round_inst_U175 ( .A(rc_27_), .B(round_inst_xin_w[27]), .Z(
        round_inst_srout2_w[11]) );
  XOR2_X1 round_inst_U174 ( .A(rc_28_), .B(round_inst_xin_w[28]), .Z(
        round_inst_srout2_w[28]) );
  XOR2_X1 round_inst_U173 ( .A(rc_29_), .B(round_inst_xin_w[29]), .Z(
        round_inst_srout2_w[29]) );
  XOR2_X1 round_inst_U172 ( .A(rc_2_), .B(round_inst_xin_w[2]), .Z(
        round_inst_srout2_w[18]) );
  XOR2_X1 round_inst_U171 ( .A(rc_30_), .B(round_inst_xin_w[30]), .Z(
        round_inst_srout2_w[30]) );
  XOR2_X1 round_inst_U170 ( .A(rc_31_), .B(round_inst_xin_w[31]), .Z(
        round_inst_srout2_w[31]) );
  XOR2_X1 round_inst_U169 ( .A(rc_32_), .B(round_inst_xin_w[32]), .Z(
        round_inst_srout2_w[48]) );
  XOR2_X1 round_inst_U168 ( .A(rc_33_), .B(round_inst_xin_w[33]), .Z(
        round_inst_srout2_w[49]) );
  XOR2_X1 round_inst_U167 ( .A(rc_34_), .B(round_inst_xin_w[34]), .Z(
        round_inst_srout2_w[50]) );
  XOR2_X1 round_inst_U166 ( .A(rc_35_), .B(round_inst_xin_w[35]), .Z(
        round_inst_srout2_w[51]) );
  XOR2_X1 round_inst_U165 ( .A(rc_36_), .B(round_inst_xin_w[36]), .Z(
        round_inst_srout2_w[4]) );
  XOR2_X1 round_inst_U164 ( .A(rc_37_), .B(round_inst_xin_w[37]), .Z(
        round_inst_srout2_w[5]) );
  XOR2_X1 round_inst_U163 ( .A(rc_38_), .B(round_inst_xin_w[38]), .Z(
        round_inst_srout2_w[6]) );
  XOR2_X1 round_inst_U162 ( .A(rc_39_), .B(round_inst_xin_w[39]), .Z(
        round_inst_srout2_w[7]) );
  XOR2_X1 round_inst_U161 ( .A(rc_3_), .B(round_inst_xin_w[3]), .Z(
        round_inst_srout2_w[19]) );
  XOR2_X1 round_inst_U160 ( .A(rc_40_), .B(round_inst_xin_w[40]), .Z(
        round_inst_srout2_w[24]) );
  XOR2_X1 round_inst_U159 ( .A(rc_41_), .B(round_inst_xin_w[41]), .Z(
        round_inst_srout2_w[25]) );
  XOR2_X1 round_inst_U158 ( .A(rc_42_), .B(round_inst_xin_w[42]), .Z(
        round_inst_srout2_w[26]) );
  XOR2_X1 round_inst_U157 ( .A(rc_43_), .B(round_inst_xin_w[43]), .Z(
        round_inst_srout2_w[27]) );
  XOR2_X1 round_inst_U156 ( .A(rc_44_), .B(round_inst_xin_w[44]), .Z(
        round_inst_srout2_w[44]) );
  XOR2_X1 round_inst_U155 ( .A(rc_45_), .B(round_inst_xin_w[45]), .Z(
        round_inst_srout2_w[45]) );
  XOR2_X1 round_inst_U154 ( .A(rc_46_), .B(round_inst_xin_w[46]), .Z(
        round_inst_srout2_w[46]) );
  XOR2_X1 round_inst_U153 ( .A(rc_47_), .B(round_inst_xin_w[47]), .Z(
        round_inst_srout2_w[47]) );
  XOR2_X1 round_inst_U152 ( .A(rc_48_), .B(round_inst_xin_w[48]), .Z(
        round_inst_srout2_w[0]) );
  XOR2_X1 round_inst_U151 ( .A(rc_49_), .B(round_inst_xin_w[49]), .Z(
        round_inst_srout2_w[1]) );
  XOR2_X1 round_inst_U150 ( .A(rc_4_), .B(round_inst_xin_w[4]), .Z(
        round_inst_srout2_w[36]) );
  XOR2_X1 round_inst_U149 ( .A(rc_50_), .B(round_inst_xin_w[50]), .Z(
        round_inst_srout2_w[2]) );
  XOR2_X1 round_inst_U148 ( .A(rc_51_), .B(round_inst_xin_w[51]), .Z(
        round_inst_srout2_w[3]) );
  XOR2_X1 round_inst_U147 ( .A(rc_52_), .B(round_inst_xin_w[52]), .Z(
        round_inst_srout2_w[20]) );
  XOR2_X1 round_inst_U146 ( .A(rc_53_), .B(round_inst_xin_w[53]), .Z(
        round_inst_srout2_w[21]) );
  XOR2_X1 round_inst_U145 ( .A(rc_54_), .B(round_inst_xin_w[54]), .Z(
        round_inst_srout2_w[22]) );
  XOR2_X1 round_inst_U144 ( .A(rc_55_), .B(round_inst_xin_w[55]), .Z(
        round_inst_srout2_w[23]) );
  XOR2_X1 round_inst_U143 ( .A(rc_56_), .B(round_inst_xin_w[56]), .Z(
        round_inst_srout2_w[40]) );
  XOR2_X1 round_inst_U142 ( .A(rc_57_), .B(round_inst_xin_w[57]), .Z(
        round_inst_srout2_w[41]) );
  XOR2_X1 round_inst_U141 ( .A(rc_58_), .B(round_inst_xin_w[58]), .Z(
        round_inst_srout2_w[42]) );
  XOR2_X1 round_inst_U140 ( .A(rc_59_), .B(round_inst_xin_w[59]), .Z(
        round_inst_srout2_w[43]) );
  XOR2_X1 round_inst_U139 ( .A(rc_5_), .B(round_inst_xin_w[5]), .Z(
        round_inst_srout2_w[37]) );
  XOR2_X1 round_inst_U138 ( .A(rc_60_), .B(round_inst_xin_w[60]), .Z(
        round_inst_srout2_w[60]) );
  XOR2_X1 round_inst_U137 ( .A(rc_61_), .B(round_inst_xin_w[61]), .Z(
        round_inst_srout2_w[61]) );
  XOR2_X1 round_inst_U136 ( .A(rc_62_), .B(round_inst_xin_w[62]), .Z(
        round_inst_srout2_w[62]) );
  XOR2_X1 round_inst_U135 ( .A(rc_63_), .B(round_inst_xin_w[63]), .Z(
        round_inst_srout2_w[63]) );
  XOR2_X1 round_inst_U134 ( .A(rc_6_), .B(round_inst_xin_w[6]), .Z(
        round_inst_srout2_w[38]) );
  XOR2_X1 round_inst_U133 ( .A(rc_7_), .B(round_inst_xin_w[7]), .Z(
        round_inst_srout2_w[39]) );
  XOR2_X1 round_inst_U132 ( .A(rc_8_), .B(round_inst_xin_w[8]), .Z(
        round_inst_srout2_w[56]) );
  XOR2_X1 round_inst_U131 ( .A(rc_9_), .B(round_inst_xin_w[9]), .Z(
        round_inst_srout2_w[57]) );
  XOR2_X1 round_inst_U130 ( .A(rc_0_), .B(round_inst_srout_w[0]), .Z(
        round_inst_xout_w[0]) );
  XOR2_X1 round_inst_U129 ( .A(rc_10_), .B(round_inst_aout_w[59]), .Z(
        round_inst_xout_w[10]) );
  XOR2_X1 round_inst_U128 ( .A(rc_11_), .B(round_inst_srout_w[11]), .Z(
        round_inst_xout_w[11]) );
  XOR2_X1 round_inst_U127 ( .A(rc_12_), .B(round_inst_srout_w[12]), .Z(
        round_inst_xout_w[12]) );
  XOR2_X1 round_inst_U126 ( .A(rc_13_), .B(round_inst_srout_w[13]), .Z(
        round_inst_xout_w[13]) );
  XOR2_X1 round_inst_U125 ( .A(rc_14_), .B(round_inst_aout_w[15]), .Z(
        round_inst_xout_w[14]) );
  XOR2_X1 round_inst_U124 ( .A(k[15]), .B(round_inst_srout_w[15]), .Z(
        round_inst_xout_w[15]) );
  XOR2_X1 round_inst_U123 ( .A(rc_16_), .B(round_inst_srout_w[16]), .Z(
        round_inst_xout_w[16]) );
  XOR2_X1 round_inst_U122 ( .A(rc_17_), .B(round_inst_srout_w[17]), .Z(
        round_inst_xout_w[17]) );
  XOR2_X1 round_inst_U121 ( .A(rc_18_), .B(round_inst_aout_w[35]), .Z(
        round_inst_xout_w[18]) );
  XOR2_X1 round_inst_U120 ( .A(rc_19_), .B(round_inst_srout_w[19]), .Z(
        round_inst_xout_w[19]) );
  XOR2_X1 round_inst_U119 ( .A(rc_1_), .B(round_inst_srout_w[1]), .Z(
        round_inst_xout_w[1]) );
  XOR2_X1 round_inst_U118 ( .A(rc_20_), .B(round_inst_srout_w[20]), .Z(
        round_inst_xout_w[20]) );
  XOR2_X1 round_inst_U117 ( .A(rc_21_), .B(round_inst_srout_w[21]), .Z(
        round_inst_xout_w[21]) );
  XOR2_X1 round_inst_U116 ( .A(rc_22_), .B(round_inst_aout_w[55]), .Z(
        round_inst_xout_w[22]) );
  XOR2_X1 round_inst_U115 ( .A(rc_23_), .B(round_inst_srout_w[23]), .Z(
        round_inst_xout_w[23]) );
  XOR2_X1 round_inst_U114 ( .A(rc_24_), .B(round_inst_srout_w[24]), .Z(
        round_inst_xout_w[24]) );
  XOR2_X1 round_inst_U113 ( .A(rc_25_), .B(round_inst_srout_w[25]), .Z(
        round_inst_xout_w[25]) );
  XOR2_X1 round_inst_U112 ( .A(rc_26_), .B(round_inst_aout_w[11]), .Z(
        round_inst_xout_w[26]) );
  XOR2_X1 round_inst_U111 ( .A(rc_27_), .B(round_inst_srout_w[27]), .Z(
        round_inst_xout_w[27]) );
  XOR2_X1 round_inst_U110 ( .A(rc_28_), .B(round_inst_srout_w[28]), .Z(
        round_inst_xout_w[28]) );
  XOR2_X1 round_inst_U109 ( .A(rc_29_), .B(round_inst_srout_w[29]), .Z(
        round_inst_xout_w[29]) );
  XOR2_X1 round_inst_U108 ( .A(rc_2_), .B(round_inst_aout_w[19]), .Z(
        round_inst_xout_w[2]) );
  XOR2_X1 round_inst_U107 ( .A(rc_30_), .B(round_inst_aout_w[31]), .Z(
        round_inst_xout_w[30]) );
  XOR2_X1 round_inst_U106 ( .A(rc_31_), .B(round_inst_srout_w[31]), .Z(
        round_inst_xout_w[31]) );
  XOR2_X1 round_inst_U105 ( .A(rc_32_), .B(round_inst_srout_w[32]), .Z(
        round_inst_xout_w[32]) );
  XOR2_X1 round_inst_U104 ( .A(rc_33_), .B(round_inst_srout_w[33]), .Z(
        round_inst_xout_w[33]) );
  XOR2_X1 round_inst_U103 ( .A(rc_34_), .B(round_inst_aout_w[51]), .Z(
        round_inst_xout_w[34]) );
  XOR2_X1 round_inst_U102 ( .A(rc_35_), .B(round_inst_srout_w[35]), .Z(
        round_inst_xout_w[35]) );
  XOR2_X1 round_inst_U101 ( .A(rc_36_), .B(round_inst_srout_w[36]), .Z(
        round_inst_xout_w[36]) );
  XOR2_X1 round_inst_U100 ( .A(rc_37_), .B(round_inst_srout_w[37]), .Z(
        round_inst_xout_w[37]) );
  XOR2_X1 round_inst_U99 ( .A(rc_38_), .B(round_inst_aout_w[7]), .Z(
        round_inst_xout_w[38]) );
  XOR2_X1 round_inst_U98 ( .A(rc_39_), .B(round_inst_srout_w[39]), .Z(
        round_inst_xout_w[39]) );
  XOR2_X1 round_inst_U97 ( .A(rc_3_), .B(round_inst_srout_w[3]), .Z(
        round_inst_xout_w[3]) );
  XOR2_X1 round_inst_U96 ( .A(rc_40_), .B(round_inst_srout_w[40]), .Z(
        round_inst_xout_w[40]) );
  XOR2_X1 round_inst_U95 ( .A(rc_41_), .B(round_inst_srout_w[41]), .Z(
        round_inst_xout_w[41]) );
  XOR2_X1 round_inst_U94 ( .A(rc_42_), .B(round_inst_aout_w[27]), .Z(
        round_inst_xout_w[42]) );
  XOR2_X1 round_inst_U93 ( .A(rc_43_), .B(round_inst_srout_w[43]), .Z(
        round_inst_xout_w[43]) );
  XOR2_X1 round_inst_U92 ( .A(rc_44_), .B(round_inst_srout_w[44]), .Z(
        round_inst_xout_w[44]) );
  XOR2_X1 round_inst_U91 ( .A(rc_45_), .B(round_inst_srout_w[45]), .Z(
        round_inst_xout_w[45]) );
  XOR2_X1 round_inst_U90 ( .A(rc_46_), .B(round_inst_aout_w[47]), .Z(
        round_inst_xout_w[46]) );
  XOR2_X1 round_inst_U89 ( .A(rc_47_), .B(round_inst_srout_w[47]), .Z(
        round_inst_xout_w[47]) );
  XOR2_X1 round_inst_U88 ( .A(rc_48_), .B(round_inst_srout_w[48]), .Z(
        round_inst_xout_w[48]) );
  XOR2_X1 round_inst_U87 ( .A(rc_49_), .B(round_inst_srout_w[49]), .Z(
        round_inst_xout_w[49]) );
  XOR2_X1 round_inst_U86 ( .A(rc_4_), .B(round_inst_srout_w[4]), .Z(
        round_inst_xout_w[4]) );
  XOR2_X1 round_inst_U85 ( .A(rc_50_), .B(round_inst_aout_w[3]), .Z(
        round_inst_xout_w[50]) );
  XOR2_X1 round_inst_U84 ( .A(rc_51_), .B(round_inst_srout_w[51]), .Z(
        round_inst_xout_w[51]) );
  XOR2_X1 round_inst_U83 ( .A(rc_52_), .B(round_inst_srout_w[52]), .Z(
        round_inst_xout_w[52]) );
  XOR2_X1 round_inst_U82 ( .A(rc_53_), .B(round_inst_srout_w[53]), .Z(
        round_inst_xout_w[53]) );
  XOR2_X1 round_inst_U81 ( .A(rc_54_), .B(round_inst_aout_w[23]), .Z(
        round_inst_xout_w[54]) );
  XOR2_X1 round_inst_U80 ( .A(rc_55_), .B(round_inst_srout_w[55]), .Z(
        round_inst_xout_w[55]) );
  XOR2_X1 round_inst_U79 ( .A(rc_56_), .B(round_inst_srout_w[56]), .Z(
        round_inst_xout_w[56]) );
  XOR2_X1 round_inst_U78 ( .A(rc_57_), .B(round_inst_srout_w[57]), .Z(
        round_inst_xout_w[57]) );
  XOR2_X1 round_inst_U77 ( .A(rc_58_), .B(round_inst_aout_w[43]), .Z(
        round_inst_xout_w[58]) );
  XOR2_X1 round_inst_U76 ( .A(rc_59_), .B(round_inst_srout_w[59]), .Z(
        round_inst_xout_w[59]) );
  XOR2_X1 round_inst_U75 ( .A(rc_5_), .B(round_inst_srout_w[5]), .Z(
        round_inst_xout_w[5]) );
  XOR2_X1 round_inst_U74 ( .A(rc_60_), .B(round_inst_srout_w[60]), .Z(
        round_inst_xout_w[60]) );
  XOR2_X1 round_inst_U73 ( .A(rc_61_), .B(round_inst_srout_w[61]), .Z(
        round_inst_xout_w[61]) );
  XOR2_X1 round_inst_U72 ( .A(rc_62_), .B(round_inst_aout_w[63]), .Z(
        round_inst_xout_w[62]) );
  XOR2_X1 round_inst_U71 ( .A(rc_63_), .B(round_inst_srout_w[63]), .Z(
        round_inst_xout_w[63]) );
  XOR2_X1 round_inst_U70 ( .A(rc_6_), .B(round_inst_aout_w[39]), .Z(
        round_inst_xout_w[6]) );
  XOR2_X1 round_inst_U69 ( .A(rc_7_), .B(round_inst_srout_w[7]), .Z(
        round_inst_xout_w[7]) );
  XOR2_X1 round_inst_U68 ( .A(rc_8_), .B(round_inst_srout_w[8]), .Z(
        round_inst_xout_w[8]) );
  XOR2_X1 round_inst_U67 ( .A(rc_9_), .B(round_inst_srout_w[9]), .Z(
        round_inst_xout_w[9]) );
  INV_X1 round_inst_U66 ( .A(round_inst_sin_x[17]), .ZN(round_inst_n38) );
  INV_X1 round_inst_U65 ( .A(round_inst_sin_y[18]), .ZN(round_inst_n37) );
  INV_X1 round_inst_U64 ( .A(round_inst_sin_y[16]), .ZN(round_inst_n36) );
  INV_X1 round_inst_U63 ( .A(round_inst_sin_y[32]), .ZN(round_inst_n35) );
  INV_X1 round_inst_U62 ( .A(round_inst_sin_x[33]), .ZN(round_inst_n34) );
  INV_X1 round_inst_U61 ( .A(round_inst_sin_y[34]), .ZN(round_inst_n33) );
  INV_X1 round_inst_U60 ( .A(round_inst_sin_y[54]), .ZN(round_inst_n32) );
  INV_X1 round_inst_U59 ( .A(round_inst_sin_x[54]), .ZN(round_inst_n31) );
  INV_X1 round_inst_U58 ( .A(round_inst_sin_x[57]), .ZN(round_inst_n30) );
  INV_X1 round_inst_U57 ( .A(round_inst_sin_y[58]), .ZN(round_inst_n29) );
  INV_X1 round_inst_U56 ( .A(round_inst_sin_y[56]), .ZN(round_inst_n28) );
  INV_X1 round_inst_U55 ( .A(round_inst_sin_y[6]), .ZN(round_inst_n27) );
  INV_X1 round_inst_U54 ( .A(round_inst_sin_y[38]), .ZN(round_inst_n26) );
  INV_X1 round_inst_U53 ( .A(round_inst_sin_y[36]), .ZN(round_inst_n25) );
  INV_X1 round_inst_U52 ( .A(round_inst_sin_x[21]), .ZN(round_inst_n24) );
  INV_X1 round_inst_U51 ( .A(round_inst_sin_y[22]), .ZN(round_inst_n23) );
  INV_X1 round_inst_U50 ( .A(round_inst_sin_y[20]), .ZN(round_inst_n22) );
  INV_X1 round_inst_U49 ( .A(round_inst_sin_y[28]), .ZN(round_inst_n21) );
  INV_X1 round_inst_U48 ( .A(round_inst_sin_x[29]), .ZN(round_inst_n20) );
  INV_X1 round_inst_U47 ( .A(round_inst_sin_y[30]), .ZN(round_inst_n19) );
  INV_X1 round_inst_U46 ( .A(round_inst_sin_y[26]), .ZN(round_inst_n18) );
  INV_X1 round_inst_U45 ( .A(round_inst_sin_x[25]), .ZN(round_inst_n17) );
  INV_X1 round_inst_U44 ( .A(round_inst_sin_y[24]), .ZN(round_inst_n16) );
  INV_X1 round_inst_U43 ( .A(round_inst_sin_y[3]), .ZN(round_inst_n15) );
  INV_X1 round_inst_U42 ( .A(round_inst_sin_w[1]), .ZN(round_inst_n14) );
  INV_X1 round_inst_U41 ( .A(round_inst_sin_x[49]), .ZN(round_inst_n13) );
  INV_X1 round_inst_U40 ( .A(round_inst_sin_y[50]), .ZN(round_inst_n12) );
  INV_X1 round_inst_U39 ( .A(round_inst_sin_y[48]), .ZN(round_inst_n11) );
  INV_X1 round_inst_U38 ( .A(round_inst_sin_y[10]), .ZN(round_inst_n10) );
  INV_X1 round_inst_U37 ( .A(round_inst_sin_y[8]), .ZN(round_inst_n9) );
  INV_X1 round_inst_U36 ( .A(round_inst_sin_x[9]), .ZN(round_inst_n8) );
  INV_X1 round_inst_U35 ( .A(round_inst_sin_z[7]), .ZN(round_inst_n7) );
  INV_X1 round_inst_U34 ( .A(round_inst_n72), .ZN(round_inst_n6) );
  INV_X2 round_inst_U33 ( .A(round_inst_n26), .ZN(round_inst_n55) );
  INV_X2 round_inst_U32 ( .A(round_inst_n8), .ZN(round_inst_n61) );
  INV_X2 round_inst_U31 ( .A(round_inst_n24), .ZN(round_inst_n63) );
  INV_X2 round_inst_U30 ( .A(round_inst_n17), .ZN(round_inst_n64) );
  INV_X2 round_inst_U29 ( .A(round_inst_n20), .ZN(round_inst_n65) );
  INV_X2 round_inst_U28 ( .A(round_inst_n34), .ZN(round_inst_n66) );
  INV_X2 round_inst_U27 ( .A(round_inst_n30), .ZN(round_inst_n69) );
  INV_X2 round_inst_U26 ( .A(round_inst_n12), .ZN(round_inst_n57) );
  INV_X2 round_inst_U25 ( .A(round_inst_n37), .ZN(round_inst_n45) );
  INV_X2 round_inst_U24 ( .A(round_inst_n27), .ZN(round_inst_n41) );
  INV_X2 round_inst_U23 ( .A(round_inst_n15), .ZN(round_inst_n40) );
  INV_X2 round_inst_U22 ( .A(round_inst_n13), .ZN(round_inst_n67) );
  INV_X2 round_inst_U21 ( .A(round_inst_n38), .ZN(round_inst_n62) );
  INV_X2 round_inst_U20 ( .A(round_inst_n10), .ZN(round_inst_n43) );
  INV_X2 round_inst_U19 ( .A(round_inst_n19), .ZN(round_inst_n51) );
  INV_X2 round_inst_U18 ( .A(round_inst_n18), .ZN(round_inst_n49) );
  INV_X2 round_inst_U17 ( .A(round_inst_n33), .ZN(round_inst_n53) );
  INV_X2 round_inst_U16 ( .A(round_inst_n29), .ZN(round_inst_n60) );
  INV_X2 round_inst_U15 ( .A(round_inst_n23), .ZN(round_inst_n47) );
  INV_X2 round_inst_U14 ( .A(round_inst_n32), .ZN(round_inst_n58) );
  INV_X2 round_inst_U13 ( .A(round_inst_n7), .ZN(round_inst_n39) );
  INV_X2 round_inst_U12 ( .A(round_inst_n9), .ZN(round_inst_n42) );
  INV_X2 round_inst_U11 ( .A(round_inst_n36), .ZN(round_inst_n44) );
  INV_X2 round_inst_U10 ( .A(round_inst_n35), .ZN(round_inst_n52) );
  INV_X2 round_inst_U9 ( .A(round_inst_n28), .ZN(round_inst_n59) );
  INV_X2 round_inst_U8 ( .A(round_inst_n22), .ZN(round_inst_n46) );
  INV_X2 round_inst_U7 ( .A(round_inst_n21), .ZN(round_inst_n50) );
  INV_X2 round_inst_U6 ( .A(round_inst_n16), .ZN(round_inst_n48) );
  INV_X2 round_inst_U5 ( .A(round_inst_n11), .ZN(round_inst_n56) );
  INV_X2 round_inst_U4 ( .A(round_inst_n25), .ZN(round_inst_n54) );
  INV_X2 round_inst_U3 ( .A(round_inst_n31), .ZN(round_inst_n68) );
  INV_X2 round_inst_U2 ( .A(round_inst_n6), .ZN(cout[0]) );
  INV_X2 round_inst_U1 ( .A(round_inst_n14), .ZN(round_inst_n70) );
  XNOR2_X1 round_inst_A_0__aw_U4 ( .A(round_inst_A_0__aw_n3), .B(
        round_inst_srout_w[48]), .ZN(round_inst_aout_w[1]) );
  XNOR2_X1 round_inst_A_0__aw_U3 ( .A(round_inst_srout_w[49]), .B(
        round_inst_aout_w[3]), .ZN(round_inst_A_0__aw_n3) );
  INV_X1 round_inst_A_0__aw_U2 ( .A(round_inst_srout_w[49]), .ZN(
        round_inst_aout_w[0]) );
  INV_X1 round_inst_A_0__aw_U1 ( .A(round_inst_srout_w[51]), .ZN(
        round_inst_aout_w[2]) );
  XNOR2_X1 round_inst_A_0__ax_U2 ( .A(round_inst_A_0__ax_n1), .B(
        round_inst_srout_x[48]), .ZN(round_inst_aout_x[1]) );
  XNOR2_X1 round_inst_A_0__ax_U1 ( .A(round_inst_aout_x[0]), .B(
        round_inst_aout_x[3]), .ZN(round_inst_A_0__ax_n1) );
  XNOR2_X1 round_inst_A_0__ay_U2 ( .A(round_inst_A_0__ay_n3), .B(
        round_inst_srout_y[48]), .ZN(round_inst_aout_y[1]) );
  XNOR2_X1 round_inst_A_0__ay_U1 ( .A(round_inst_aout_y[0]), .B(
        round_inst_aout_y[3]), .ZN(round_inst_A_0__ay_n3) );
  XNOR2_X1 round_inst_A_0__az_U2 ( .A(round_inst_A_0__az_n3), .B(
        round_inst_srout_z[48]), .ZN(round_inst_aout_z[1]) );
  XNOR2_X1 round_inst_A_0__az_U1 ( .A(round_inst_aout_z[0]), .B(
        round_inst_aout_z[3]), .ZN(round_inst_A_0__az_n3) );
  XNOR2_X1 round_inst_A_1__aw_U4 ( .A(round_inst_A_1__aw_n5), .B(
        round_inst_srout_w[36]), .ZN(round_inst_aout_w[5]) );
  XNOR2_X1 round_inst_A_1__aw_U3 ( .A(round_inst_srout_w[37]), .B(
        round_inst_aout_w[7]), .ZN(round_inst_A_1__aw_n5) );
  INV_X1 round_inst_A_1__aw_U2 ( .A(round_inst_srout_w[37]), .ZN(
        round_inst_aout_w[4]) );
  INV_X1 round_inst_A_1__aw_U1 ( .A(round_inst_srout_w[39]), .ZN(
        round_inst_aout_w[6]) );
  XNOR2_X1 round_inst_A_1__ax_U2 ( .A(round_inst_A_1__ax_n3), .B(
        round_inst_srout_x[36]), .ZN(round_inst_aout_x[5]) );
  XNOR2_X1 round_inst_A_1__ax_U1 ( .A(round_inst_aout_x[4]), .B(
        round_inst_aout_x[7]), .ZN(round_inst_A_1__ax_n3) );
  XNOR2_X1 round_inst_A_1__ay_U2 ( .A(round_inst_A_1__ay_n3), .B(
        round_inst_srout_y[36]), .ZN(round_inst_aout_y[5]) );
  XNOR2_X1 round_inst_A_1__ay_U1 ( .A(round_inst_aout_y[4]), .B(
        round_inst_aout_y[7]), .ZN(round_inst_A_1__ay_n3) );
  XNOR2_X1 round_inst_A_1__az_U2 ( .A(round_inst_A_1__az_n3), .B(
        round_inst_srout_z[36]), .ZN(round_inst_aout_z[5]) );
  XNOR2_X1 round_inst_A_1__az_U1 ( .A(round_inst_aout_z[4]), .B(
        round_inst_aout_z[7]), .ZN(round_inst_A_1__az_n3) );
  XNOR2_X1 round_inst_A_2__aw_U4 ( .A(round_inst_A_2__aw_n5), .B(
        round_inst_srout_w[24]), .ZN(round_inst_aout_w[9]) );
  XNOR2_X1 round_inst_A_2__aw_U3 ( .A(round_inst_srout_w[25]), .B(
        round_inst_aout_w[11]), .ZN(round_inst_A_2__aw_n5) );
  INV_X1 round_inst_A_2__aw_U2 ( .A(round_inst_srout_w[25]), .ZN(
        round_inst_aout_w[8]) );
  INV_X1 round_inst_A_2__aw_U1 ( .A(round_inst_srout_w[27]), .ZN(
        round_inst_aout_w[10]) );
  XNOR2_X1 round_inst_A_2__ax_U2 ( .A(round_inst_A_2__ax_n3), .B(
        round_inst_srout_x[24]), .ZN(round_inst_aout_x[9]) );
  XNOR2_X1 round_inst_A_2__ax_U1 ( .A(round_inst_aout_x[8]), .B(
        round_inst_aout_x[11]), .ZN(round_inst_A_2__ax_n3) );
  XNOR2_X1 round_inst_A_2__ay_U2 ( .A(round_inst_A_2__ay_n3), .B(
        round_inst_srout_y[24]), .ZN(round_inst_aout_y[9]) );
  XNOR2_X1 round_inst_A_2__ay_U1 ( .A(round_inst_aout_y[8]), .B(
        round_inst_aout_y[11]), .ZN(round_inst_A_2__ay_n3) );
  XNOR2_X1 round_inst_A_2__az_U2 ( .A(round_inst_A_2__az_n3), .B(
        round_inst_srout_z[24]), .ZN(round_inst_aout_z[9]) );
  XNOR2_X1 round_inst_A_2__az_U1 ( .A(round_inst_aout_z[8]), .B(
        round_inst_aout_z[11]), .ZN(round_inst_A_2__az_n3) );
  XNOR2_X1 round_inst_A_3__aw_U4 ( .A(round_inst_A_3__aw_n5), .B(
        round_inst_srout_w[12]), .ZN(round_inst_aout_w[13]) );
  XNOR2_X1 round_inst_A_3__aw_U3 ( .A(round_inst_srout_w[13]), .B(
        round_inst_aout_w[15]), .ZN(round_inst_A_3__aw_n5) );
  INV_X1 round_inst_A_3__aw_U2 ( .A(round_inst_srout_w[13]), .ZN(
        round_inst_aout_w[12]) );
  INV_X1 round_inst_A_3__aw_U1 ( .A(round_inst_srout_w[15]), .ZN(
        round_inst_aout_w[14]) );
  XNOR2_X1 round_inst_A_3__ax_U2 ( .A(round_inst_A_3__ax_n3), .B(
        round_inst_srout_x[12]), .ZN(round_inst_aout_x[13]) );
  XNOR2_X1 round_inst_A_3__ax_U1 ( .A(round_inst_aout_x[12]), .B(
        round_inst_aout_x[15]), .ZN(round_inst_A_3__ax_n3) );
  XNOR2_X1 round_inst_A_3__ay_U2 ( .A(round_inst_A_3__ay_n3), .B(
        round_inst_srout_y[12]), .ZN(round_inst_aout_y[13]) );
  XNOR2_X1 round_inst_A_3__ay_U1 ( .A(round_inst_aout_y[12]), .B(
        round_inst_aout_y[15]), .ZN(round_inst_A_3__ay_n3) );
  XNOR2_X1 round_inst_A_3__az_U2 ( .A(round_inst_A_3__az_n3), .B(
        round_inst_srout_z[12]), .ZN(round_inst_aout_z[13]) );
  XNOR2_X1 round_inst_A_3__az_U1 ( .A(round_inst_aout_z[12]), .B(
        round_inst_aout_z[15]), .ZN(round_inst_A_3__az_n3) );
  XNOR2_X1 round_inst_A_4__aw_U4 ( .A(round_inst_A_4__aw_n5), .B(
        round_inst_srout_w[0]), .ZN(round_inst_aout_w[17]) );
  XNOR2_X1 round_inst_A_4__aw_U3 ( .A(round_inst_srout_w[1]), .B(
        round_inst_aout_w[19]), .ZN(round_inst_A_4__aw_n5) );
  INV_X1 round_inst_A_4__aw_U2 ( .A(round_inst_srout_w[1]), .ZN(
        round_inst_aout_w[16]) );
  INV_X1 round_inst_A_4__aw_U1 ( .A(round_inst_srout_w[3]), .ZN(
        round_inst_aout_w[18]) );
  XNOR2_X1 round_inst_A_4__ax_U2 ( .A(round_inst_A_4__ax_n3), .B(
        round_inst_srout_x[0]), .ZN(round_inst_aout_x[17]) );
  XNOR2_X1 round_inst_A_4__ax_U1 ( .A(round_inst_aout_x[16]), .B(
        round_inst_aout_x[19]), .ZN(round_inst_A_4__ax_n3) );
  XNOR2_X1 round_inst_A_4__ay_U2 ( .A(round_inst_A_4__ay_n3), .B(
        round_inst_srout_y[0]), .ZN(round_inst_aout_y[17]) );
  XNOR2_X1 round_inst_A_4__ay_U1 ( .A(round_inst_aout_y[16]), .B(
        round_inst_aout_y[19]), .ZN(round_inst_A_4__ay_n3) );
  XNOR2_X1 round_inst_A_4__az_U2 ( .A(round_inst_A_4__az_n3), .B(
        round_inst_srout_z[0]), .ZN(round_inst_aout_z[17]) );
  XNOR2_X1 round_inst_A_4__az_U1 ( .A(round_inst_aout_z[16]), .B(
        round_inst_aout_z[19]), .ZN(round_inst_A_4__az_n3) );
  XNOR2_X1 round_inst_A_5__aw_U4 ( .A(round_inst_A_5__aw_n5), .B(
        round_inst_srout_w[52]), .ZN(round_inst_aout_w[21]) );
  XNOR2_X1 round_inst_A_5__aw_U3 ( .A(round_inst_srout_w[53]), .B(
        round_inst_aout_w[23]), .ZN(round_inst_A_5__aw_n5) );
  INV_X1 round_inst_A_5__aw_U2 ( .A(round_inst_srout_w[53]), .ZN(
        round_inst_aout_w[20]) );
  INV_X1 round_inst_A_5__aw_U1 ( .A(round_inst_srout_w[55]), .ZN(
        round_inst_aout_w[22]) );
  XNOR2_X1 round_inst_A_5__ax_U2 ( .A(round_inst_A_5__ax_n3), .B(
        round_inst_srout_x[52]), .ZN(round_inst_aout_x[21]) );
  XNOR2_X1 round_inst_A_5__ax_U1 ( .A(round_inst_aout_x[20]), .B(
        round_inst_aout_x[23]), .ZN(round_inst_A_5__ax_n3) );
  XNOR2_X1 round_inst_A_5__ay_U2 ( .A(round_inst_A_5__ay_n3), .B(
        round_inst_srout_y[52]), .ZN(round_inst_aout_y[21]) );
  XNOR2_X1 round_inst_A_5__ay_U1 ( .A(round_inst_aout_y[20]), .B(
        round_inst_aout_y[23]), .ZN(round_inst_A_5__ay_n3) );
  XNOR2_X1 round_inst_A_5__az_U2 ( .A(round_inst_A_5__az_n3), .B(
        round_inst_srout_z[52]), .ZN(round_inst_aout_z[21]) );
  XNOR2_X1 round_inst_A_5__az_U1 ( .A(round_inst_aout_z[20]), .B(
        round_inst_aout_z[23]), .ZN(round_inst_A_5__az_n3) );
  XNOR2_X1 round_inst_A_6__aw_U4 ( .A(round_inst_A_6__aw_n5), .B(
        round_inst_srout_w[40]), .ZN(round_inst_aout_w[25]) );
  XNOR2_X1 round_inst_A_6__aw_U3 ( .A(round_inst_srout_w[41]), .B(
        round_inst_aout_w[27]), .ZN(round_inst_A_6__aw_n5) );
  INV_X1 round_inst_A_6__aw_U2 ( .A(round_inst_srout_w[41]), .ZN(
        round_inst_aout_w[24]) );
  INV_X1 round_inst_A_6__aw_U1 ( .A(round_inst_srout_w[43]), .ZN(
        round_inst_aout_w[26]) );
  XNOR2_X1 round_inst_A_6__ax_U2 ( .A(round_inst_A_6__ax_n3), .B(
        round_inst_srout_x[40]), .ZN(round_inst_aout_x[25]) );
  XNOR2_X1 round_inst_A_6__ax_U1 ( .A(round_inst_aout_x[24]), .B(
        round_inst_aout_x[27]), .ZN(round_inst_A_6__ax_n3) );
  XNOR2_X1 round_inst_A_6__ay_U2 ( .A(round_inst_A_6__ay_n3), .B(
        round_inst_srout_y[40]), .ZN(round_inst_aout_y[25]) );
  XNOR2_X1 round_inst_A_6__ay_U1 ( .A(round_inst_aout_y[24]), .B(
        round_inst_aout_y[27]), .ZN(round_inst_A_6__ay_n3) );
  XNOR2_X1 round_inst_A_6__az_U2 ( .A(round_inst_A_6__az_n3), .B(
        round_inst_srout_z[40]), .ZN(round_inst_aout_z[25]) );
  XNOR2_X1 round_inst_A_6__az_U1 ( .A(round_inst_aout_z[24]), .B(
        round_inst_aout_z[27]), .ZN(round_inst_A_6__az_n3) );
  XNOR2_X1 round_inst_A_7__aw_U4 ( .A(round_inst_A_7__aw_n5), .B(
        round_inst_srout_w[28]), .ZN(round_inst_aout_w[29]) );
  XNOR2_X1 round_inst_A_7__aw_U3 ( .A(round_inst_srout_w[29]), .B(
        round_inst_aout_w[31]), .ZN(round_inst_A_7__aw_n5) );
  INV_X1 round_inst_A_7__aw_U2 ( .A(round_inst_srout_w[29]), .ZN(
        round_inst_aout_w[28]) );
  INV_X1 round_inst_A_7__aw_U1 ( .A(round_inst_srout_w[31]), .ZN(
        round_inst_aout_w[30]) );
  XNOR2_X1 round_inst_A_7__ax_U2 ( .A(round_inst_A_7__ax_n3), .B(
        round_inst_srout_x[28]), .ZN(round_inst_aout_x[29]) );
  XNOR2_X1 round_inst_A_7__ax_U1 ( .A(round_inst_aout_x[28]), .B(
        round_inst_aout_x[31]), .ZN(round_inst_A_7__ax_n3) );
  XNOR2_X1 round_inst_A_7__ay_U2 ( .A(round_inst_A_7__ay_n3), .B(
        round_inst_srout_y[28]), .ZN(round_inst_aout_y[29]) );
  XNOR2_X1 round_inst_A_7__ay_U1 ( .A(round_inst_aout_y[28]), .B(
        round_inst_aout_y[31]), .ZN(round_inst_A_7__ay_n3) );
  XNOR2_X1 round_inst_A_7__az_U2 ( .A(round_inst_A_7__az_n3), .B(
        round_inst_srout_z[28]), .ZN(round_inst_aout_z[29]) );
  XNOR2_X1 round_inst_A_7__az_U1 ( .A(round_inst_aout_z[28]), .B(
        round_inst_aout_z[31]), .ZN(round_inst_A_7__az_n3) );
  XNOR2_X1 round_inst_A_8__aw_U4 ( .A(round_inst_A_8__aw_n5), .B(
        round_inst_srout_w[16]), .ZN(round_inst_aout_w[33]) );
  XNOR2_X1 round_inst_A_8__aw_U3 ( .A(round_inst_srout_w[17]), .B(
        round_inst_aout_w[35]), .ZN(round_inst_A_8__aw_n5) );
  INV_X1 round_inst_A_8__aw_U2 ( .A(round_inst_srout_w[17]), .ZN(
        round_inst_aout_w[32]) );
  INV_X1 round_inst_A_8__aw_U1 ( .A(round_inst_srout_w[19]), .ZN(
        round_inst_aout_w[34]) );
  XNOR2_X1 round_inst_A_8__ax_U2 ( .A(round_inst_A_8__ax_n3), .B(
        round_inst_srout_x[16]), .ZN(round_inst_aout_x[33]) );
  XNOR2_X1 round_inst_A_8__ax_U1 ( .A(round_inst_aout_x[32]), .B(
        round_inst_aout_x[35]), .ZN(round_inst_A_8__ax_n3) );
  XNOR2_X1 round_inst_A_8__ay_U2 ( .A(round_inst_A_8__ay_n3), .B(
        round_inst_srout_y[16]), .ZN(round_inst_aout_y[33]) );
  XNOR2_X1 round_inst_A_8__ay_U1 ( .A(round_inst_aout_y[32]), .B(
        round_inst_aout_y[35]), .ZN(round_inst_A_8__ay_n3) );
  XNOR2_X1 round_inst_A_8__az_U2 ( .A(round_inst_A_8__az_n3), .B(
        round_inst_srout_z[16]), .ZN(round_inst_aout_z[33]) );
  XNOR2_X1 round_inst_A_8__az_U1 ( .A(round_inst_aout_z[32]), .B(
        round_inst_aout_z[35]), .ZN(round_inst_A_8__az_n3) );
  XNOR2_X1 round_inst_A_9__aw_U4 ( .A(round_inst_A_9__aw_n5), .B(
        round_inst_srout_w[4]), .ZN(round_inst_aout_w[37]) );
  XNOR2_X1 round_inst_A_9__aw_U3 ( .A(round_inst_srout_w[5]), .B(
        round_inst_aout_w[39]), .ZN(round_inst_A_9__aw_n5) );
  INV_X1 round_inst_A_9__aw_U2 ( .A(round_inst_srout_w[5]), .ZN(
        round_inst_aout_w[36]) );
  INV_X1 round_inst_A_9__aw_U1 ( .A(round_inst_srout_w[7]), .ZN(
        round_inst_aout_w[38]) );
  XNOR2_X1 round_inst_A_9__ax_U2 ( .A(round_inst_A_9__ax_n3), .B(
        round_inst_srout_x[4]), .ZN(round_inst_aout_x[37]) );
  XNOR2_X1 round_inst_A_9__ax_U1 ( .A(round_inst_aout_x[36]), .B(
        round_inst_aout_x[39]), .ZN(round_inst_A_9__ax_n3) );
  XNOR2_X1 round_inst_A_9__ay_U2 ( .A(round_inst_A_9__ay_n3), .B(
        round_inst_srout_y[4]), .ZN(round_inst_aout_y[37]) );
  XNOR2_X1 round_inst_A_9__ay_U1 ( .A(round_inst_aout_y[36]), .B(
        round_inst_aout_y[39]), .ZN(round_inst_A_9__ay_n3) );
  XNOR2_X1 round_inst_A_9__az_U2 ( .A(round_inst_A_9__az_n3), .B(
        round_inst_srout_z[4]), .ZN(round_inst_aout_z[37]) );
  XNOR2_X1 round_inst_A_9__az_U1 ( .A(round_inst_aout_z[36]), .B(
        round_inst_aout_z[39]), .ZN(round_inst_A_9__az_n3) );
  XNOR2_X1 round_inst_A_10__aw_U4 ( .A(round_inst_A_10__aw_n5), .B(
        round_inst_srout_w[56]), .ZN(round_inst_aout_w[41]) );
  XNOR2_X1 round_inst_A_10__aw_U3 ( .A(round_inst_srout_w[57]), .B(
        round_inst_aout_w[43]), .ZN(round_inst_A_10__aw_n5) );
  INV_X1 round_inst_A_10__aw_U2 ( .A(round_inst_srout_w[57]), .ZN(
        round_inst_aout_w[40]) );
  INV_X1 round_inst_A_10__aw_U1 ( .A(round_inst_srout_w[59]), .ZN(
        round_inst_aout_w[42]) );
  XNOR2_X1 round_inst_A_10__ax_U2 ( .A(round_inst_A_10__ax_n3), .B(
        round_inst_srout_x[56]), .ZN(round_inst_aout_x[41]) );
  XNOR2_X1 round_inst_A_10__ax_U1 ( .A(round_inst_aout_x[40]), .B(
        round_inst_aout_x[43]), .ZN(round_inst_A_10__ax_n3) );
  XNOR2_X1 round_inst_A_10__ay_U2 ( .A(round_inst_A_10__ay_n3), .B(
        round_inst_srout_y[56]), .ZN(round_inst_aout_y[41]) );
  XNOR2_X1 round_inst_A_10__ay_U1 ( .A(round_inst_aout_y[40]), .B(
        round_inst_aout_y[43]), .ZN(round_inst_A_10__ay_n3) );
  XNOR2_X1 round_inst_A_10__az_U2 ( .A(round_inst_A_10__az_n3), .B(
        round_inst_srout_z[56]), .ZN(round_inst_aout_z[41]) );
  XNOR2_X1 round_inst_A_10__az_U1 ( .A(round_inst_aout_z[40]), .B(
        round_inst_aout_z[43]), .ZN(round_inst_A_10__az_n3) );
  XNOR2_X1 round_inst_A_11__aw_U4 ( .A(round_inst_A_11__aw_n5), .B(
        round_inst_srout_w[44]), .ZN(round_inst_aout_w[45]) );
  XNOR2_X1 round_inst_A_11__aw_U3 ( .A(round_inst_srout_w[45]), .B(
        round_inst_aout_w[47]), .ZN(round_inst_A_11__aw_n5) );
  INV_X1 round_inst_A_11__aw_U2 ( .A(round_inst_srout_w[45]), .ZN(
        round_inst_aout_w[44]) );
  INV_X1 round_inst_A_11__aw_U1 ( .A(round_inst_srout_w[47]), .ZN(
        round_inst_aout_w[46]) );
  XNOR2_X1 round_inst_A_11__ax_U2 ( .A(round_inst_A_11__ax_n3), .B(
        round_inst_srout_x[44]), .ZN(round_inst_aout_x[45]) );
  XNOR2_X1 round_inst_A_11__ax_U1 ( .A(round_inst_aout_x[44]), .B(
        round_inst_aout_x[47]), .ZN(round_inst_A_11__ax_n3) );
  XNOR2_X1 round_inst_A_11__ay_U2 ( .A(round_inst_A_11__ay_n3), .B(
        round_inst_srout_y[44]), .ZN(round_inst_aout_y[45]) );
  XNOR2_X1 round_inst_A_11__ay_U1 ( .A(round_inst_aout_y[44]), .B(
        round_inst_aout_y[47]), .ZN(round_inst_A_11__ay_n3) );
  XNOR2_X1 round_inst_A_11__az_U2 ( .A(round_inst_A_11__az_n3), .B(
        round_inst_srout_z[44]), .ZN(round_inst_aout_z[45]) );
  XNOR2_X1 round_inst_A_11__az_U1 ( .A(round_inst_aout_z[44]), .B(
        round_inst_aout_z[47]), .ZN(round_inst_A_11__az_n3) );
  XNOR2_X1 round_inst_A_12__aw_U4 ( .A(round_inst_A_12__aw_n5), .B(
        round_inst_srout_w[32]), .ZN(round_inst_aout_w[49]) );
  XNOR2_X1 round_inst_A_12__aw_U3 ( .A(round_inst_srout_w[33]), .B(
        round_inst_aout_w[51]), .ZN(round_inst_A_12__aw_n5) );
  INV_X1 round_inst_A_12__aw_U2 ( .A(round_inst_srout_w[33]), .ZN(
        round_inst_aout_w[48]) );
  INV_X1 round_inst_A_12__aw_U1 ( .A(round_inst_srout_w[35]), .ZN(
        round_inst_aout_w[50]) );
  XNOR2_X1 round_inst_A_12__ax_U2 ( .A(round_inst_A_12__ax_n3), .B(
        round_inst_srout_x[32]), .ZN(round_inst_aout_x[49]) );
  XNOR2_X1 round_inst_A_12__ax_U1 ( .A(round_inst_aout_x[48]), .B(
        round_inst_aout_x[51]), .ZN(round_inst_A_12__ax_n3) );
  XNOR2_X1 round_inst_A_12__ay_U2 ( .A(round_inst_A_12__ay_n3), .B(
        round_inst_srout_y[32]), .ZN(round_inst_aout_y[49]) );
  XNOR2_X1 round_inst_A_12__ay_U1 ( .A(round_inst_aout_y[48]), .B(
        round_inst_aout_y[51]), .ZN(round_inst_A_12__ay_n3) );
  XNOR2_X1 round_inst_A_12__az_U2 ( .A(round_inst_A_12__az_n3), .B(
        round_inst_srout_z[32]), .ZN(round_inst_aout_z[49]) );
  XNOR2_X1 round_inst_A_12__az_U1 ( .A(round_inst_aout_z[48]), .B(
        round_inst_aout_z[51]), .ZN(round_inst_A_12__az_n3) );
  XNOR2_X1 round_inst_A_13__aw_U4 ( .A(round_inst_A_13__aw_n5), .B(
        round_inst_srout_w[20]), .ZN(round_inst_aout_w[53]) );
  XNOR2_X1 round_inst_A_13__aw_U3 ( .A(round_inst_srout_w[21]), .B(
        round_inst_aout_w[55]), .ZN(round_inst_A_13__aw_n5) );
  INV_X1 round_inst_A_13__aw_U2 ( .A(round_inst_srout_w[23]), .ZN(
        round_inst_aout_w[54]) );
  INV_X1 round_inst_A_13__aw_U1 ( .A(round_inst_srout_w[21]), .ZN(
        round_inst_aout_w[52]) );
  XNOR2_X1 round_inst_A_13__ax_U2 ( .A(round_inst_A_13__ax_n3), .B(
        round_inst_srout_x[20]), .ZN(round_inst_aout_x[53]) );
  XNOR2_X1 round_inst_A_13__ax_U1 ( .A(round_inst_aout_x[52]), .B(
        round_inst_aout_x[55]), .ZN(round_inst_A_13__ax_n3) );
  XNOR2_X1 round_inst_A_13__ay_U2 ( .A(round_inst_A_13__ay_n3), .B(
        round_inst_srout_y[20]), .ZN(round_inst_aout_y[53]) );
  XNOR2_X1 round_inst_A_13__ay_U1 ( .A(round_inst_aout_y[52]), .B(
        round_inst_aout_y[55]), .ZN(round_inst_A_13__ay_n3) );
  XNOR2_X1 round_inst_A_13__az_U2 ( .A(round_inst_A_13__az_n3), .B(
        round_inst_srout_z[20]), .ZN(round_inst_aout_z[53]) );
  XNOR2_X1 round_inst_A_13__az_U1 ( .A(round_inst_aout_z[52]), .B(
        round_inst_aout_z[55]), .ZN(round_inst_A_13__az_n3) );
  XNOR2_X1 round_inst_A_14__aw_U4 ( .A(round_inst_A_14__aw_n5), .B(
        round_inst_srout_w[8]), .ZN(round_inst_aout_w[57]) );
  XNOR2_X1 round_inst_A_14__aw_U3 ( .A(round_inst_srout_w[9]), .B(
        round_inst_aout_w[59]), .ZN(round_inst_A_14__aw_n5) );
  INV_X1 round_inst_A_14__aw_U2 ( .A(round_inst_srout_w[9]), .ZN(
        round_inst_aout_w[56]) );
  INV_X1 round_inst_A_14__aw_U1 ( .A(round_inst_srout_w[11]), .ZN(
        round_inst_aout_w[58]) );
  XNOR2_X1 round_inst_A_14__ax_U2 ( .A(round_inst_A_14__ax_n3), .B(
        round_inst_srout_x[8]), .ZN(round_inst_aout_x[57]) );
  XNOR2_X1 round_inst_A_14__ax_U1 ( .A(round_inst_aout_x[56]), .B(
        round_inst_aout_x[59]), .ZN(round_inst_A_14__ax_n3) );
  XNOR2_X1 round_inst_A_14__ay_U2 ( .A(round_inst_A_14__ay_n3), .B(
        round_inst_srout_y[8]), .ZN(round_inst_aout_y[57]) );
  XNOR2_X1 round_inst_A_14__ay_U1 ( .A(round_inst_aout_y[56]), .B(
        round_inst_aout_y[59]), .ZN(round_inst_A_14__ay_n3) );
  XNOR2_X1 round_inst_A_14__az_U2 ( .A(round_inst_A_14__az_n3), .B(
        round_inst_srout_z[8]), .ZN(round_inst_aout_z[57]) );
  XNOR2_X1 round_inst_A_14__az_U1 ( .A(round_inst_aout_z[56]), .B(
        round_inst_aout_z[59]), .ZN(round_inst_A_14__az_n3) );
  XNOR2_X1 round_inst_A_15__aw_U4 ( .A(round_inst_A_15__aw_n5), .B(
        round_inst_srout_w[60]), .ZN(round_inst_aout_w[61]) );
  XNOR2_X1 round_inst_A_15__aw_U3 ( .A(round_inst_srout_w[61]), .B(
        round_inst_aout_w[63]), .ZN(round_inst_A_15__aw_n5) );
  INV_X1 round_inst_A_15__aw_U2 ( .A(round_inst_srout_w[63]), .ZN(
        round_inst_aout_w[62]) );
  INV_X1 round_inst_A_15__aw_U1 ( .A(round_inst_srout_w[61]), .ZN(
        round_inst_aout_w[60]) );
  XNOR2_X1 round_inst_A_15__ax_U2 ( .A(round_inst_A_15__ax_n3), .B(
        round_inst_srout_x[60]), .ZN(round_inst_aout_x[61]) );
  XNOR2_X1 round_inst_A_15__ax_U1 ( .A(round_inst_aout_x[60]), .B(
        round_inst_aout_x[63]), .ZN(round_inst_A_15__ax_n3) );
  XNOR2_X1 round_inst_A_15__ay_U2 ( .A(round_inst_A_15__ay_n3), .B(
        round_inst_srout_y[60]), .ZN(round_inst_aout_y[61]) );
  XNOR2_X1 round_inst_A_15__ay_U1 ( .A(round_inst_aout_y[60]), .B(
        round_inst_aout_y[63]), .ZN(round_inst_A_15__ay_n3) );
  XNOR2_X1 round_inst_A_15__az_U2 ( .A(round_inst_A_15__az_n3), .B(
        round_inst_srout_z[60]), .ZN(round_inst_aout_z[61]) );
  XNOR2_X1 round_inst_A_15__az_U1 ( .A(round_inst_aout_z[60]), .B(
        round_inst_aout_z[63]), .ZN(round_inst_A_15__az_n3) );
  MUX2_X1 round_inst_mux_inv_w_U68 ( .A(round_inst_aout_w[60]), .B(
        round_inst_xout_w[60]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[60]) );
  MUX2_X1 round_inst_mux_inv_w_U67 ( .A(round_inst_aout_w[56]), .B(
        round_inst_xout_w[56]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[56]) );
  MUX2_X1 round_inst_mux_inv_w_U66 ( .A(round_inst_aout_w[52]), .B(
        round_inst_xout_w[52]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[52]) );
  MUX2_X1 round_inst_mux_inv_w_U65 ( .A(round_inst_aout_w[48]), .B(
        round_inst_xout_w[48]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[48]) );
  MUX2_X1 round_inst_mux_inv_w_U64 ( .A(round_inst_aout_w[44]), .B(
        round_inst_xout_w[44]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[44]) );
  MUX2_X1 round_inst_mux_inv_w_U63 ( .A(round_inst_aout_w[40]), .B(
        round_inst_xout_w[40]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[40]) );
  MUX2_X1 round_inst_mux_inv_w_U62 ( .A(round_inst_aout_w[36]), .B(
        round_inst_xout_w[36]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[36]) );
  MUX2_X1 round_inst_mux_inv_w_U61 ( .A(round_inst_aout_w[32]), .B(
        round_inst_xout_w[32]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[32]) );
  MUX2_X1 round_inst_mux_inv_w_U60 ( .A(round_inst_aout_w[28]), .B(
        round_inst_xout_w[28]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[28]) );
  MUX2_X1 round_inst_mux_inv_w_U59 ( .A(round_inst_aout_w[24]), .B(
        round_inst_xout_w[24]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[24]) );
  MUX2_X1 round_inst_mux_inv_w_U58 ( .A(round_inst_aout_w[20]), .B(
        round_inst_xout_w[20]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[20]) );
  MUX2_X1 round_inst_mux_inv_w_U57 ( .A(round_inst_aout_w[16]), .B(
        round_inst_xout_w[16]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[16]) );
  MUX2_X1 round_inst_mux_inv_w_U56 ( .A(round_inst_aout_w[12]), .B(
        round_inst_xout_w[12]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[12]) );
  MUX2_X1 round_inst_mux_inv_w_U55 ( .A(round_inst_aout_w[8]), .B(
        round_inst_xout_w[8]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[8]) );
  MUX2_X1 round_inst_mux_inv_w_U54 ( .A(round_inst_aout_w[4]), .B(
        round_inst_xout_w[4]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[4]) );
  MUX2_X1 round_inst_mux_inv_w_U53 ( .A(round_inst_aout_w[0]), .B(
        round_inst_xout_w[0]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[0]) );
  MUX2_X1 round_inst_mux_inv_w_U52 ( .A(round_inst_aout_w[62]), .B(
        round_inst_xout_w[62]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[62]) );
  MUX2_X1 round_inst_mux_inv_w_U51 ( .A(round_inst_aout_w[58]), .B(
        round_inst_xout_w[58]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[58]) );
  MUX2_X1 round_inst_mux_inv_w_U50 ( .A(round_inst_aout_w[54]), .B(
        round_inst_xout_w[54]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[54]) );
  MUX2_X1 round_inst_mux_inv_w_U49 ( .A(round_inst_aout_w[42]), .B(
        round_inst_xout_w[42]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[42]) );
  MUX2_X1 round_inst_mux_inv_w_U48 ( .A(round_inst_aout_w[38]), .B(
        round_inst_xout_w[38]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[38]) );
  MUX2_X1 round_inst_mux_inv_w_U47 ( .A(round_inst_aout_w[34]), .B(
        round_inst_xout_w[34]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[34]) );
  MUX2_X1 round_inst_mux_inv_w_U46 ( .A(round_inst_aout_w[26]), .B(
        round_inst_xout_w[26]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[26]) );
  MUX2_X1 round_inst_mux_inv_w_U45 ( .A(round_inst_aout_w[22]), .B(
        round_inst_xout_w[22]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[22]) );
  MUX2_X1 round_inst_mux_inv_w_U44 ( .A(round_inst_aout_w[14]), .B(
        round_inst_xout_w[14]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[14]) );
  MUX2_X1 round_inst_mux_inv_w_U43 ( .A(round_inst_aout_w[46]), .B(
        round_inst_xout_w[46]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[46]) );
  MUX2_X1 round_inst_mux_inv_w_U42 ( .A(round_inst_aout_w[10]), .B(
        round_inst_xout_w[10]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[10]) );
  MUX2_X1 round_inst_mux_inv_w_U41 ( .A(round_inst_aout_w[2]), .B(
        round_inst_xout_w[2]), .S(round_inst_mux_inv_w_n266), .Z(
        round_inst_sin_w[2]) );
  MUX2_X1 round_inst_mux_inv_w_U40 ( .A(round_inst_aout_w[61]), .B(
        round_inst_xout_w[61]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[61]) );
  MUX2_X1 round_inst_mux_inv_w_U39 ( .A(round_inst_aout_w[63]), .B(
        round_inst_xout_w[63]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[63]) );
  MUX2_X1 round_inst_mux_inv_w_U38 ( .A(round_inst_aout_w[57]), .B(
        round_inst_xout_w[57]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[57]) );
  MUX2_X1 round_inst_mux_inv_w_U37 ( .A(round_inst_aout_w[59]), .B(
        round_inst_xout_w[59]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[59]) );
  MUX2_X1 round_inst_mux_inv_w_U36 ( .A(round_inst_aout_w[53]), .B(
        round_inst_xout_w[53]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[53]) );
  MUX2_X1 round_inst_mux_inv_w_U35 ( .A(round_inst_aout_w[55]), .B(
        round_inst_xout_w[55]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[55]) );
  MUX2_X1 round_inst_mux_inv_w_U34 ( .A(round_inst_aout_w[49]), .B(
        round_inst_xout_w[49]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[49]) );
  MUX2_X1 round_inst_mux_inv_w_U33 ( .A(round_inst_aout_w[51]), .B(
        round_inst_xout_w[51]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[51]) );
  MUX2_X1 round_inst_mux_inv_w_U32 ( .A(round_inst_aout_w[45]), .B(
        round_inst_xout_w[45]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[45]) );
  MUX2_X1 round_inst_mux_inv_w_U31 ( .A(round_inst_aout_w[47]), .B(
        round_inst_xout_w[47]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[47]) );
  MUX2_X1 round_inst_mux_inv_w_U30 ( .A(round_inst_aout_w[41]), .B(
        round_inst_xout_w[41]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[41]) );
  MUX2_X1 round_inst_mux_inv_w_U29 ( .A(round_inst_aout_w[43]), .B(
        round_inst_xout_w[43]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[43]) );
  MUX2_X1 round_inst_mux_inv_w_U28 ( .A(round_inst_aout_w[37]), .B(
        round_inst_xout_w[37]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[37]) );
  MUX2_X1 round_inst_mux_inv_w_U27 ( .A(round_inst_aout_w[39]), .B(
        round_inst_xout_w[39]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[39]) );
  MUX2_X1 round_inst_mux_inv_w_U26 ( .A(round_inst_aout_w[33]), .B(
        round_inst_xout_w[33]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[33]) );
  MUX2_X1 round_inst_mux_inv_w_U25 ( .A(round_inst_aout_w[35]), .B(
        round_inst_xout_w[35]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[35]) );
  MUX2_X1 round_inst_mux_inv_w_U24 ( .A(round_inst_aout_w[29]), .B(
        round_inst_xout_w[29]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[29]) );
  MUX2_X1 round_inst_mux_inv_w_U23 ( .A(round_inst_aout_w[31]), .B(
        round_inst_xout_w[31]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[31]) );
  MUX2_X1 round_inst_mux_inv_w_U22 ( .A(round_inst_aout_w[25]), .B(
        round_inst_xout_w[25]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[25]) );
  MUX2_X1 round_inst_mux_inv_w_U21 ( .A(round_inst_aout_w[21]), .B(
        round_inst_xout_w[21]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[21]) );
  MUX2_X1 round_inst_mux_inv_w_U20 ( .A(round_inst_aout_w[23]), .B(
        round_inst_xout_w[23]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[23]) );
  MUX2_X1 round_inst_mux_inv_w_U19 ( .A(round_inst_aout_w[17]), .B(
        round_inst_xout_w[17]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[17]) );
  MUX2_X1 round_inst_mux_inv_w_U18 ( .A(round_inst_aout_w[19]), .B(
        round_inst_xout_w[19]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[19]) );
  MUX2_X1 round_inst_mux_inv_w_U17 ( .A(round_inst_aout_w[13]), .B(
        round_inst_xout_w[13]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[13]) );
  MUX2_X1 round_inst_mux_inv_w_U16 ( .A(round_inst_aout_w[15]), .B(
        round_inst_xout_w[15]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[15]) );
  MUX2_X1 round_inst_mux_inv_w_U15 ( .A(round_inst_aout_w[9]), .B(
        round_inst_xout_w[9]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[9]) );
  MUX2_X1 round_inst_mux_inv_w_U14 ( .A(round_inst_aout_w[11]), .B(
        round_inst_xout_w[11]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[11]) );
  MUX2_X1 round_inst_mux_inv_w_U13 ( .A(round_inst_aout_w[5]), .B(
        round_inst_xout_w[5]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[5]) );
  MUX2_X1 round_inst_mux_inv_w_U12 ( .A(round_inst_aout_w[7]), .B(
        round_inst_xout_w[7]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[7]) );
  MUX2_X1 round_inst_mux_inv_w_U11 ( .A(round_inst_aout_w[1]), .B(
        round_inst_xout_w[1]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[1]) );
  MUX2_X1 round_inst_mux_inv_w_U10 ( .A(round_inst_aout_w[3]), .B(
        round_inst_xout_w[3]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[3]) );
  MUX2_X1 round_inst_mux_inv_w_U9 ( .A(round_inst_aout_w[50]), .B(
        round_inst_xout_w[50]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[50]) );
  MUX2_X1 round_inst_mux_inv_w_U8 ( .A(round_inst_aout_w[30]), .B(
        round_inst_xout_w[30]), .S(round_inst_mux_inv_w_n265), .Z(
        round_inst_sin_w[30]) );
  INV_X1 round_inst_mux_inv_w_U7 ( .A(round_inst_mux_inv_w_n263), .ZN(
        round_inst_mux_inv_w_n265) );
  MUX2_X1 round_inst_mux_inv_w_U6 ( .A(round_inst_aout_w[27]), .B(
        round_inst_xout_w[27]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[27]) );
  MUX2_X1 round_inst_mux_inv_w_U5 ( .A(round_inst_aout_w[18]), .B(
        round_inst_xout_w[18]), .S(round_inst_mux_inv_w_n264), .Z(
        round_inst_sin_w[18]) );
  INV_X1 round_inst_mux_inv_w_U4 ( .A(round_inst_mux_inv_w_n263), .ZN(
        round_inst_mux_inv_w_n264) );
  MUX2_X1 round_inst_mux_inv_w_U3 ( .A(round_inst_aout_w[6]), .B(
        round_inst_xout_w[6]), .S(inv_sig), .Z(round_inst_sin_w[6]) );
  INV_X1 round_inst_mux_inv_w_U2 ( .A(inv_sig), .ZN(round_inst_mux_inv_w_n263)
         );
  INV_X2 round_inst_mux_inv_w_U1 ( .A(round_inst_mux_inv_w_n263), .ZN(
        round_inst_mux_inv_w_n266) );
  MUX2_X1 round_inst_mux_inv_x_U68 ( .A(round_inst_aout_x[63]), .B(
        round_inst_aout_x[62]), .S(round_inst_mux_inv_x_n266), .Z(bout[3]) );
  MUX2_X1 round_inst_mux_inv_x_U67 ( .A(round_inst_aout_x[55]), .B(
        round_inst_aout_x[22]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[55]) );
  MUX2_X1 round_inst_mux_inv_x_U66 ( .A(round_inst_aout_x[51]), .B(
        round_inst_aout_x[2]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[51]) );
  MUX2_X1 round_inst_mux_inv_x_U65 ( .A(round_inst_aout_x[59]), .B(
        round_inst_aout_x[42]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[59]) );
  MUX2_X1 round_inst_mux_inv_x_U64 ( .A(round_inst_aout_x[31]), .B(
        round_inst_aout_x[30]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[31]) );
  MUX2_X1 round_inst_mux_inv_x_U63 ( .A(round_inst_aout_x[19]), .B(
        round_inst_aout_x[34]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[19]) );
  MUX2_X1 round_inst_mux_inv_x_U62 ( .A(round_inst_aout_x[47]), .B(
        round_inst_aout_x[46]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[47]) );
  MUX2_X1 round_inst_mux_inv_x_U61 ( .A(round_inst_aout_x[39]), .B(
        round_inst_aout_x[6]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[39]) );
  MUX2_X1 round_inst_mux_inv_x_U60 ( .A(round_inst_aout_x[35]), .B(
        round_inst_aout_x[50]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[35]) );
  MUX2_X1 round_inst_mux_inv_x_U59 ( .A(round_inst_aout_x[15]), .B(
        round_inst_aout_x[14]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[15]) );
  MUX2_X1 round_inst_mux_inv_x_U58 ( .A(round_inst_aout_x[43]), .B(
        round_inst_aout_x[26]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[43]) );
  MUX2_X1 round_inst_mux_inv_x_U57 ( .A(round_inst_aout_x[3]), .B(
        round_inst_aout_x[18]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[3]) );
  MUX2_X1 round_inst_mux_inv_x_U56 ( .A(round_inst_aout_x[23]), .B(
        round_inst_aout_x[54]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[23]) );
  MUX2_X1 round_inst_mux_inv_x_U55 ( .A(round_inst_aout_x[27]), .B(
        round_inst_aout_x[10]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[27]) );
  MUX2_X1 round_inst_mux_inv_x_U54 ( .A(round_inst_aout_x[11]), .B(
        round_inst_aout_x[58]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[11]) );
  MUX2_X1 round_inst_mux_inv_x_U53 ( .A(round_inst_aout_x[7]), .B(
        round_inst_aout_x[38]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[7]) );
  MUX2_X1 round_inst_mux_inv_x_U52 ( .A(round_inst_aout_x[62]), .B(
        round_inst_aout_x[63]), .S(round_inst_mux_inv_x_n266), .Z(bout[2]) );
  MUX2_X1 round_inst_mux_inv_x_U51 ( .A(round_inst_aout_x[61]), .B(
        round_inst_aout_x[60]), .S(round_inst_mux_inv_x_n266), .Z(bout[1]) );
  MUX2_X1 round_inst_mux_inv_x_U50 ( .A(round_inst_aout_x[60]), .B(
        round_inst_srout_x[60]), .S(round_inst_mux_inv_x_n266), .Z(bout[0]) );
  MUX2_X1 round_inst_mux_inv_x_U49 ( .A(round_inst_aout_x[58]), .B(
        round_inst_aout_x[43]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[58]) );
  MUX2_X1 round_inst_mux_inv_x_U48 ( .A(round_inst_aout_x[54]), .B(
        round_inst_aout_x[23]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[54]) );
  MUX2_X1 round_inst_mux_inv_x_U47 ( .A(round_inst_aout_x[50]), .B(
        round_inst_aout_x[3]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[50]) );
  MUX2_X1 round_inst_mux_inv_x_U46 ( .A(round_inst_aout_x[46]), .B(
        round_inst_aout_x[47]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[46]) );
  MUX2_X1 round_inst_mux_inv_x_U45 ( .A(round_inst_aout_x[45]), .B(
        round_inst_aout_x[44]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[45]) );
  MUX2_X1 round_inst_mux_inv_x_U44 ( .A(round_inst_aout_x[42]), .B(
        round_inst_aout_x[27]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[42]) );
  MUX2_X1 round_inst_mux_inv_x_U43 ( .A(round_inst_aout_x[38]), .B(
        round_inst_aout_x[7]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[38]) );
  MUX2_X1 round_inst_mux_inv_x_U42 ( .A(round_inst_aout_x[34]), .B(
        round_inst_aout_x[51]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[34]) );
  MUX2_X1 round_inst_mux_inv_x_U41 ( .A(round_inst_aout_x[30]), .B(
        round_inst_aout_x[31]), .S(round_inst_mux_inv_x_n266), .Z(
        round_inst_sin_x[30]) );
  MUX2_X1 round_inst_mux_inv_x_U40 ( .A(round_inst_aout_x[26]), .B(
        round_inst_aout_x[11]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[26]) );
  MUX2_X1 round_inst_mux_inv_x_U39 ( .A(round_inst_aout_x[25]), .B(
        round_inst_aout_x[8]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[25]) );
  MUX2_X1 round_inst_mux_inv_x_U38 ( .A(round_inst_aout_x[22]), .B(
        round_inst_aout_x[55]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[22]) );
  MUX2_X1 round_inst_mux_inv_x_U37 ( .A(round_inst_aout_x[18]), .B(
        round_inst_aout_x[35]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[18]) );
  MUX2_X1 round_inst_mux_inv_x_U36 ( .A(round_inst_aout_x[14]), .B(
        round_inst_aout_x[15]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[14]) );
  MUX2_X1 round_inst_mux_inv_x_U35 ( .A(round_inst_aout_x[13]), .B(
        round_inst_aout_x[12]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[13]) );
  MUX2_X1 round_inst_mux_inv_x_U34 ( .A(round_inst_aout_x[10]), .B(
        round_inst_aout_x[59]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[10]) );
  MUX2_X1 round_inst_mux_inv_x_U33 ( .A(round_inst_aout_x[6]), .B(
        round_inst_aout_x[39]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[6]) );
  MUX2_X1 round_inst_mux_inv_x_U32 ( .A(round_inst_aout_x[1]), .B(
        round_inst_aout_x[16]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[1]) );
  MUX2_X1 round_inst_mux_inv_x_U31 ( .A(round_inst_aout_x[57]), .B(
        round_inst_aout_x[40]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[57]) );
  MUX2_X1 round_inst_mux_inv_x_U30 ( .A(round_inst_aout_x[53]), .B(
        round_inst_aout_x[20]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[53]) );
  MUX2_X1 round_inst_mux_inv_x_U29 ( .A(round_inst_aout_x[49]), .B(
        round_inst_aout_x[0]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[49]) );
  MUX2_X1 round_inst_mux_inv_x_U28 ( .A(round_inst_aout_x[41]), .B(
        round_inst_aout_x[24]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[41]) );
  MUX2_X1 round_inst_mux_inv_x_U27 ( .A(round_inst_aout_x[37]), .B(
        round_inst_aout_x[4]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[37]) );
  MUX2_X1 round_inst_mux_inv_x_U26 ( .A(round_inst_aout_x[33]), .B(
        round_inst_aout_x[48]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[33]) );
  MUX2_X1 round_inst_mux_inv_x_U25 ( .A(round_inst_aout_x[29]), .B(
        round_inst_aout_x[28]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[29]) );
  MUX2_X1 round_inst_mux_inv_x_U24 ( .A(round_inst_aout_x[21]), .B(
        round_inst_aout_x[52]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[21]) );
  MUX2_X1 round_inst_mux_inv_x_U23 ( .A(round_inst_aout_x[17]), .B(
        round_inst_aout_x[32]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[17]) );
  MUX2_X1 round_inst_mux_inv_x_U22 ( .A(round_inst_aout_x[9]), .B(
        round_inst_aout_x[56]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[9]) );
  MUX2_X1 round_inst_mux_inv_x_U21 ( .A(round_inst_aout_x[5]), .B(
        round_inst_aout_x[36]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[5]) );
  MUX2_X1 round_inst_mux_inv_x_U20 ( .A(round_inst_aout_x[56]), .B(
        round_inst_srout_x[56]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[56]) );
  MUX2_X1 round_inst_mux_inv_x_U19 ( .A(round_inst_aout_x[52]), .B(
        round_inst_srout_x[52]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[52]) );
  MUX2_X1 round_inst_mux_inv_x_U18 ( .A(round_inst_aout_x[48]), .B(
        round_inst_srout_x[48]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[48]) );
  MUX2_X1 round_inst_mux_inv_x_U17 ( .A(round_inst_aout_x[36]), .B(
        round_inst_srout_x[36]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[36]) );
  MUX2_X1 round_inst_mux_inv_x_U16 ( .A(round_inst_aout_x[32]), .B(
        round_inst_srout_x[32]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[32]) );
  MUX2_X1 round_inst_mux_inv_x_U15 ( .A(round_inst_aout_x[28]), .B(
        round_inst_srout_x[28]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[28]) );
  MUX2_X1 round_inst_mux_inv_x_U14 ( .A(round_inst_aout_x[24]), .B(
        round_inst_srout_x[24]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[24]) );
  MUX2_X1 round_inst_mux_inv_x_U13 ( .A(round_inst_aout_x[20]), .B(
        round_inst_srout_x[20]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[20]) );
  MUX2_X1 round_inst_mux_inv_x_U12 ( .A(round_inst_aout_x[16]), .B(
        round_inst_srout_x[16]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[16]) );
  MUX2_X1 round_inst_mux_inv_x_U11 ( .A(round_inst_aout_x[8]), .B(
        round_inst_srout_x[8]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[8]) );
  MUX2_X1 round_inst_mux_inv_x_U10 ( .A(round_inst_aout_x[4]), .B(
        round_inst_srout_x[4]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[4]) );
  INV_X1 round_inst_mux_inv_x_U9 ( .A(round_inst_mux_inv_x_n263), .ZN(
        round_inst_mux_inv_x_n264) );
  MUX2_X1 round_inst_mux_inv_x_U8 ( .A(round_inst_aout_x[0]), .B(
        round_inst_srout_x[0]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[0]) );
  INV_X1 round_inst_mux_inv_x_U7 ( .A(round_inst_mux_inv_x_n263), .ZN(
        round_inst_mux_inv_x_n265) );
  INV_X1 round_inst_mux_inv_x_U6 ( .A(inv_sig), .ZN(round_inst_mux_inv_x_n263)
         );
  INV_X2 round_inst_mux_inv_x_U5 ( .A(round_inst_mux_inv_x_n263), .ZN(
        round_inst_mux_inv_x_n266) );
  MUX2_X2 round_inst_mux_inv_x_U4 ( .A(round_inst_aout_x[2]), .B(
        round_inst_aout_x[19]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[2]) );
  MUX2_X2 round_inst_mux_inv_x_U3 ( .A(round_inst_aout_x[40]), .B(
        round_inst_srout_x[40]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[40]) );
  MUX2_X2 round_inst_mux_inv_x_U2 ( .A(round_inst_aout_x[44]), .B(
        round_inst_srout_x[44]), .S(round_inst_mux_inv_x_n265), .Z(
        round_inst_sin_x[44]) );
  MUX2_X2 round_inst_mux_inv_x_U1 ( .A(round_inst_aout_x[12]), .B(
        round_inst_srout_x[12]), .S(round_inst_mux_inv_x_n264), .Z(
        round_inst_sin_x[12]) );
  MUX2_X1 round_inst_mux_inv_y_U70 ( .A(round_inst_aout_y[63]), .B(
        round_inst_aout_y[62]), .S(round_inst_mux_inv_y_n268), .Z(cout[3]) );
  MUX2_X1 round_inst_mux_inv_y_U69 ( .A(round_inst_aout_y[62]), .B(
        round_inst_aout_y[63]), .S(round_inst_mux_inv_y_n268), .Z(cout[2]) );
  MUX2_X1 round_inst_mux_inv_y_U68 ( .A(round_inst_aout_y[61]), .B(
        round_inst_aout_y[60]), .S(round_inst_mux_inv_y_n268), .Z(cout[1]) );
  MUX2_X1 round_inst_mux_inv_y_U67 ( .A(round_inst_aout_y[60]), .B(
        round_inst_srout_y[60]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_n72) );
  MUX2_X1 round_inst_mux_inv_y_U66 ( .A(round_inst_aout_y[56]), .B(
        round_inst_srout_y[56]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[56]) );
  MUX2_X1 round_inst_mux_inv_y_U65 ( .A(round_inst_aout_y[57]), .B(
        round_inst_aout_y[40]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[57]) );
  MUX2_X1 round_inst_mux_inv_y_U64 ( .A(round_inst_aout_y[52]), .B(
        round_inst_srout_y[52]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_mux_inv_y_n269) );
  MUX2_X1 round_inst_mux_inv_y_U63 ( .A(round_inst_aout_y[53]), .B(
        round_inst_aout_y[20]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[53]) );
  MUX2_X1 round_inst_mux_inv_y_U62 ( .A(round_inst_aout_y[48]), .B(
        round_inst_srout_y[48]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[48]) );
  MUX2_X1 round_inst_mux_inv_y_U61 ( .A(round_inst_aout_y[49]), .B(
        round_inst_aout_y[0]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[49]) );
  MUX2_X1 round_inst_mux_inv_y_U60 ( .A(round_inst_aout_y[44]), .B(
        round_inst_srout_y[44]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[44]) );
  MUX2_X1 round_inst_mux_inv_y_U59 ( .A(round_inst_aout_y[45]), .B(
        round_inst_aout_y[44]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[45]) );
  MUX2_X1 round_inst_mux_inv_y_U58 ( .A(round_inst_aout_y[40]), .B(
        round_inst_srout_y[40]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[40]) );
  MUX2_X1 round_inst_mux_inv_y_U57 ( .A(round_inst_aout_y[41]), .B(
        round_inst_aout_y[24]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[41]) );
  MUX2_X1 round_inst_mux_inv_y_U56 ( .A(round_inst_aout_y[36]), .B(
        round_inst_srout_y[36]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[36]) );
  MUX2_X1 round_inst_mux_inv_y_U55 ( .A(round_inst_aout_y[37]), .B(
        round_inst_aout_y[4]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[37]) );
  MUX2_X1 round_inst_mux_inv_y_U54 ( .A(round_inst_aout_y[32]), .B(
        round_inst_srout_y[32]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[32]) );
  MUX2_X1 round_inst_mux_inv_y_U53 ( .A(round_inst_aout_y[33]), .B(
        round_inst_aout_y[48]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[33]) );
  MUX2_X1 round_inst_mux_inv_y_U52 ( .A(round_inst_aout_y[28]), .B(
        round_inst_srout_y[28]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[28]) );
  MUX2_X1 round_inst_mux_inv_y_U51 ( .A(round_inst_aout_y[29]), .B(
        round_inst_aout_y[28]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[29]) );
  MUX2_X1 round_inst_mux_inv_y_U50 ( .A(round_inst_aout_y[24]), .B(
        round_inst_srout_y[24]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[24]) );
  MUX2_X1 round_inst_mux_inv_y_U49 ( .A(round_inst_aout_y[25]), .B(
        round_inst_aout_y[8]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[25]) );
  MUX2_X1 round_inst_mux_inv_y_U48 ( .A(round_inst_aout_y[20]), .B(
        round_inst_srout_y[20]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[20]) );
  MUX2_X1 round_inst_mux_inv_y_U47 ( .A(round_inst_aout_y[21]), .B(
        round_inst_aout_y[52]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[21]) );
  MUX2_X1 round_inst_mux_inv_y_U46 ( .A(round_inst_aout_y[16]), .B(
        round_inst_srout_y[16]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[16]) );
  MUX2_X1 round_inst_mux_inv_y_U45 ( .A(round_inst_aout_y[17]), .B(
        round_inst_aout_y[32]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[17]) );
  MUX2_X1 round_inst_mux_inv_y_U44 ( .A(round_inst_aout_y[12]), .B(
        round_inst_srout_y[12]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[12]) );
  MUX2_X1 round_inst_mux_inv_y_U43 ( .A(round_inst_aout_y[13]), .B(
        round_inst_aout_y[12]), .S(round_inst_mux_inv_y_n268), .Z(
        round_inst_sin_y[13]) );
  MUX2_X1 round_inst_mux_inv_y_U42 ( .A(round_inst_aout_y[8]), .B(
        round_inst_srout_y[8]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[8]) );
  MUX2_X1 round_inst_mux_inv_y_U41 ( .A(round_inst_aout_y[9]), .B(
        round_inst_aout_y[56]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[9]) );
  MUX2_X1 round_inst_mux_inv_y_U40 ( .A(round_inst_aout_y[5]), .B(
        round_inst_aout_y[36]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[5]) );
  MUX2_X1 round_inst_mux_inv_y_U39 ( .A(round_inst_aout_y[0]), .B(
        round_inst_srout_y[0]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[0]) );
  MUX2_X1 round_inst_mux_inv_y_U38 ( .A(round_inst_aout_y[1]), .B(
        round_inst_aout_y[16]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[1]) );
  MUX2_X1 round_inst_mux_inv_y_U37 ( .A(round_inst_aout_y[58]), .B(
        round_inst_aout_y[43]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[58]) );
  MUX2_X1 round_inst_mux_inv_y_U36 ( .A(round_inst_aout_y[54]), .B(
        round_inst_aout_y[23]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[54]) );
  MUX2_X1 round_inst_mux_inv_y_U35 ( .A(round_inst_aout_y[50]), .B(
        round_inst_aout_y[3]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[50]) );
  MUX2_X1 round_inst_mux_inv_y_U34 ( .A(round_inst_aout_y[46]), .B(
        round_inst_aout_y[47]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[46]) );
  MUX2_X1 round_inst_mux_inv_y_U33 ( .A(round_inst_aout_y[42]), .B(
        round_inst_aout_y[27]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[42]) );
  MUX2_X1 round_inst_mux_inv_y_U32 ( .A(round_inst_aout_y[38]), .B(
        round_inst_aout_y[7]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[38]) );
  MUX2_X1 round_inst_mux_inv_y_U31 ( .A(round_inst_aout_y[34]), .B(
        round_inst_aout_y[51]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[34]) );
  MUX2_X1 round_inst_mux_inv_y_U30 ( .A(round_inst_aout_y[30]), .B(
        round_inst_aout_y[31]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[30]) );
  MUX2_X1 round_inst_mux_inv_y_U29 ( .A(round_inst_aout_y[26]), .B(
        round_inst_aout_y[11]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[26]) );
  MUX2_X1 round_inst_mux_inv_y_U28 ( .A(round_inst_aout_y[22]), .B(
        round_inst_aout_y[55]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[22]) );
  MUX2_X1 round_inst_mux_inv_y_U27 ( .A(round_inst_aout_y[18]), .B(
        round_inst_aout_y[35]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[18]) );
  MUX2_X1 round_inst_mux_inv_y_U26 ( .A(round_inst_aout_y[14]), .B(
        round_inst_aout_y[15]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[14]) );
  MUX2_X1 round_inst_mux_inv_y_U25 ( .A(round_inst_aout_y[10]), .B(
        round_inst_aout_y[59]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[10]) );
  MUX2_X1 round_inst_mux_inv_y_U24 ( .A(round_inst_aout_y[6]), .B(
        round_inst_aout_y[39]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[6]) );
  MUX2_X1 round_inst_mux_inv_y_U23 ( .A(round_inst_aout_y[2]), .B(
        round_inst_aout_y[19]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[2]) );
  MUX2_X1 round_inst_mux_inv_y_U22 ( .A(round_inst_aout_y[59]), .B(
        round_inst_aout_y[42]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[59]) );
  MUX2_X1 round_inst_mux_inv_y_U21 ( .A(round_inst_aout_y[55]), .B(
        round_inst_aout_y[22]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[55]) );
  MUX2_X1 round_inst_mux_inv_y_U20 ( .A(round_inst_aout_y[51]), .B(
        round_inst_aout_y[2]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[51]) );
  MUX2_X1 round_inst_mux_inv_y_U19 ( .A(round_inst_aout_y[47]), .B(
        round_inst_aout_y[46]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[47]) );
  MUX2_X1 round_inst_mux_inv_y_U18 ( .A(round_inst_aout_y[43]), .B(
        round_inst_aout_y[26]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[43]) );
  MUX2_X1 round_inst_mux_inv_y_U17 ( .A(round_inst_aout_y[39]), .B(
        round_inst_aout_y[6]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[39]) );
  MUX2_X1 round_inst_mux_inv_y_U16 ( .A(round_inst_aout_y[35]), .B(
        round_inst_aout_y[50]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[35]) );
  MUX2_X1 round_inst_mux_inv_y_U15 ( .A(round_inst_aout_y[31]), .B(
        round_inst_aout_y[30]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[31]) );
  MUX2_X1 round_inst_mux_inv_y_U14 ( .A(round_inst_aout_y[27]), .B(
        round_inst_aout_y[10]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[27]) );
  MUX2_X1 round_inst_mux_inv_y_U13 ( .A(round_inst_aout_y[23]), .B(
        round_inst_aout_y[54]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[23]) );
  MUX2_X1 round_inst_mux_inv_y_U12 ( .A(round_inst_aout_y[19]), .B(
        round_inst_aout_y[34]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[19]) );
  MUX2_X1 round_inst_mux_inv_y_U11 ( .A(round_inst_aout_y[15]), .B(
        round_inst_aout_y[14]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[15]) );
  MUX2_X1 round_inst_mux_inv_y_U10 ( .A(round_inst_aout_y[11]), .B(
        round_inst_aout_y[58]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[11]) );
  MUX2_X1 round_inst_mux_inv_y_U9 ( .A(round_inst_aout_y[7]), .B(
        round_inst_aout_y[38]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[7]) );
  MUX2_X1 round_inst_mux_inv_y_U8 ( .A(round_inst_aout_y[3]), .B(
        round_inst_aout_y[18]), .S(round_inst_mux_inv_y_n266), .Z(
        round_inst_sin_y[3]) );
  INV_X1 round_inst_mux_inv_y_U7 ( .A(round_inst_mux_inv_y_n265), .ZN(
        round_inst_mux_inv_y_n266) );
  INV_X1 round_inst_mux_inv_y_U6 ( .A(round_inst_mux_inv_y_n265), .ZN(
        round_inst_mux_inv_y_n267) );
  INV_X1 round_inst_mux_inv_y_U5 ( .A(inv_sig), .ZN(round_inst_mux_inv_y_n265)
         );
  INV_X2 round_inst_mux_inv_y_U4 ( .A(round_inst_mux_inv_y_n263), .ZN(
        round_inst_sin_y[52]) );
  INV_X1 round_inst_mux_inv_y_U3 ( .A(round_inst_mux_inv_y_n269), .ZN(
        round_inst_mux_inv_y_n263) );
  INV_X2 round_inst_mux_inv_y_U2 ( .A(round_inst_mux_inv_y_n265), .ZN(
        round_inst_mux_inv_y_n268) );
  MUX2_X2 round_inst_mux_inv_y_U1 ( .A(round_inst_aout_y[4]), .B(
        round_inst_srout_y[4]), .S(round_inst_mux_inv_y_n267), .Z(
        round_inst_sin_y[4]) );
  MUX2_X1 round_inst_mux_inv_z_U69 ( .A(round_inst_aout_z[63]), .B(
        round_inst_aout_z[62]), .S(round_inst_mux_inv_z_n267), .Z(dout[3]) );
  MUX2_X1 round_inst_mux_inv_z_U68 ( .A(round_inst_aout_z[62]), .B(
        round_inst_aout_z[63]), .S(round_inst_mux_inv_z_n267), .Z(dout[2]) );
  MUX2_X1 round_inst_mux_inv_z_U67 ( .A(round_inst_aout_z[61]), .B(
        round_inst_aout_z[60]), .S(round_inst_mux_inv_z_n267), .Z(dout[1]) );
  MUX2_X1 round_inst_mux_inv_z_U66 ( .A(round_inst_aout_z[60]), .B(
        round_inst_srout_z[60]), .S(round_inst_mux_inv_z_n267), .Z(dout[0]) );
  MUX2_X1 round_inst_mux_inv_z_U65 ( .A(round_inst_aout_z[58]), .B(
        round_inst_aout_z[43]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[58]) );
  MUX2_X1 round_inst_mux_inv_z_U64 ( .A(round_inst_aout_z[59]), .B(
        round_inst_aout_z[42]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[59]) );
  MUX2_X1 round_inst_mux_inv_z_U63 ( .A(round_inst_aout_z[57]), .B(
        round_inst_aout_z[40]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[57]) );
  MUX2_X1 round_inst_mux_inv_z_U62 ( .A(round_inst_aout_z[54]), .B(
        round_inst_aout_z[23]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[54]) );
  MUX2_X1 round_inst_mux_inv_z_U61 ( .A(round_inst_aout_z[53]), .B(
        round_inst_aout_z[20]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[53]) );
  MUX2_X1 round_inst_mux_inv_z_U60 ( .A(round_inst_aout_z[50]), .B(
        round_inst_aout_z[3]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[50]) );
  MUX2_X1 round_inst_mux_inv_z_U59 ( .A(round_inst_aout_z[51]), .B(
        round_inst_aout_z[2]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[51]) );
  MUX2_X1 round_inst_mux_inv_z_U58 ( .A(round_inst_aout_z[49]), .B(
        round_inst_aout_z[0]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[49]) );
  MUX2_X1 round_inst_mux_inv_z_U57 ( .A(round_inst_aout_z[46]), .B(
        round_inst_aout_z[47]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[46]) );
  MUX2_X1 round_inst_mux_inv_z_U56 ( .A(round_inst_aout_z[42]), .B(
        round_inst_aout_z[27]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[42]) );
  MUX2_X1 round_inst_mux_inv_z_U55 ( .A(round_inst_aout_z[38]), .B(
        round_inst_aout_z[7]), .S(round_inst_mux_inv_z_n267), .Z(
        round_inst_sin_z[38]) );
  MUX2_X1 round_inst_mux_inv_z_U54 ( .A(round_inst_aout_z[39]), .B(
        round_inst_aout_z[6]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[39]) );
  MUX2_X1 round_inst_mux_inv_z_U53 ( .A(round_inst_aout_z[37]), .B(
        round_inst_aout_z[4]), .S(round_inst_mux_inv_z_n267), .Z(
        round_inst_sin_z[37]) );
  MUX2_X1 round_inst_mux_inv_z_U52 ( .A(round_inst_aout_z[34]), .B(
        round_inst_aout_z[51]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[34]) );
  MUX2_X1 round_inst_mux_inv_z_U51 ( .A(round_inst_aout_z[35]), .B(
        round_inst_aout_z[50]), .S(round_inst_mux_inv_z_n267), .Z(
        round_inst_sin_z[35]) );
  MUX2_X1 round_inst_mux_inv_z_U50 ( .A(round_inst_aout_z[33]), .B(
        round_inst_aout_z[48]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[33]) );
  MUX2_X1 round_inst_mux_inv_z_U49 ( .A(round_inst_aout_z[30]), .B(
        round_inst_aout_z[31]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[30]) );
  MUX2_X1 round_inst_mux_inv_z_U48 ( .A(round_inst_aout_z[31]), .B(
        round_inst_aout_z[30]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[31]) );
  INV_X1 round_inst_mux_inv_z_U47 ( .A(round_inst_mux_inv_z_n263), .ZN(
        round_inst_mux_inv_z_n266) );
  MUX2_X1 round_inst_mux_inv_z_U46 ( .A(round_inst_aout_z[29]), .B(
        round_inst_aout_z[28]), .S(round_inst_mux_inv_z_n267), .Z(
        round_inst_sin_z[29]) );
  MUX2_X1 round_inst_mux_inv_z_U45 ( .A(round_inst_aout_z[26]), .B(
        round_inst_aout_z[11]), .S(round_inst_mux_inv_z_n267), .Z(
        round_inst_sin_z[26]) );
  MUX2_X1 round_inst_mux_inv_z_U44 ( .A(round_inst_aout_z[27]), .B(
        round_inst_aout_z[10]), .S(round_inst_mux_inv_z_n267), .Z(
        round_inst_sin_z[27]) );
  INV_X1 round_inst_mux_inv_z_U43 ( .A(round_inst_mux_inv_z_n263), .ZN(
        round_inst_mux_inv_z_n267) );
  MUX2_X1 round_inst_mux_inv_z_U42 ( .A(round_inst_aout_z[22]), .B(
        round_inst_aout_z[55]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[22]) );
  MUX2_X1 round_inst_mux_inv_z_U41 ( .A(round_inst_aout_z[23]), .B(
        round_inst_aout_z[54]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[23]) );
  MUX2_X1 round_inst_mux_inv_z_U40 ( .A(round_inst_aout_z[21]), .B(
        round_inst_aout_z[52]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[21]) );
  MUX2_X1 round_inst_mux_inv_z_U39 ( .A(round_inst_aout_z[18]), .B(
        round_inst_aout_z[35]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[18]) );
  MUX2_X1 round_inst_mux_inv_z_U38 ( .A(round_inst_aout_z[19]), .B(
        round_inst_aout_z[34]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[19]) );
  MUX2_X1 round_inst_mux_inv_z_U37 ( .A(round_inst_aout_z[17]), .B(
        round_inst_aout_z[32]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[17]) );
  MUX2_X1 round_inst_mux_inv_z_U36 ( .A(round_inst_aout_z[14]), .B(
        round_inst_aout_z[15]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[14]) );
  MUX2_X1 round_inst_mux_inv_z_U35 ( .A(round_inst_aout_z[10]), .B(
        round_inst_aout_z[59]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[10]) );
  MUX2_X1 round_inst_mux_inv_z_U34 ( .A(round_inst_aout_z[11]), .B(
        round_inst_aout_z[58]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[11]) );
  MUX2_X1 round_inst_mux_inv_z_U33 ( .A(round_inst_aout_z[9]), .B(
        round_inst_aout_z[56]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[9]) );
  MUX2_X1 round_inst_mux_inv_z_U32 ( .A(round_inst_aout_z[6]), .B(
        round_inst_aout_z[39]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[6]) );
  MUX2_X1 round_inst_mux_inv_z_U31 ( .A(round_inst_aout_z[7]), .B(
        round_inst_aout_z[38]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[7]) );
  MUX2_X1 round_inst_mux_inv_z_U30 ( .A(round_inst_aout_z[2]), .B(
        round_inst_aout_z[19]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[2]) );
  MUX2_X1 round_inst_mux_inv_z_U29 ( .A(round_inst_aout_z[56]), .B(
        round_inst_srout_z[56]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[56]) );
  MUX2_X1 round_inst_mux_inv_z_U28 ( .A(round_inst_aout_z[52]), .B(
        round_inst_srout_z[52]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[52]) );
  MUX2_X1 round_inst_mux_inv_z_U27 ( .A(round_inst_aout_z[48]), .B(
        round_inst_srout_z[48]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[48]) );
  MUX2_X1 round_inst_mux_inv_z_U26 ( .A(round_inst_aout_z[44]), .B(
        round_inst_srout_z[44]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[44]) );
  MUX2_X1 round_inst_mux_inv_z_U25 ( .A(round_inst_aout_z[45]), .B(
        round_inst_aout_z[44]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[45]) );
  MUX2_X1 round_inst_mux_inv_z_U24 ( .A(round_inst_aout_z[40]), .B(
        round_inst_srout_z[40]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[40]) );
  MUX2_X1 round_inst_mux_inv_z_U23 ( .A(round_inst_aout_z[41]), .B(
        round_inst_aout_z[24]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[41]) );
  MUX2_X1 round_inst_mux_inv_z_U22 ( .A(round_inst_aout_z[36]), .B(
        round_inst_srout_z[36]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[36]) );
  MUX2_X1 round_inst_mux_inv_z_U21 ( .A(round_inst_aout_z[32]), .B(
        round_inst_srout_z[32]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[32]) );
  MUX2_X1 round_inst_mux_inv_z_U20 ( .A(round_inst_aout_z[28]), .B(
        round_inst_srout_z[28]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[28]) );
  MUX2_X1 round_inst_mux_inv_z_U19 ( .A(round_inst_aout_z[24]), .B(
        round_inst_srout_z[24]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[24]) );
  MUX2_X1 round_inst_mux_inv_z_U18 ( .A(round_inst_aout_z[25]), .B(
        round_inst_aout_z[8]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[25]) );
  MUX2_X1 round_inst_mux_inv_z_U17 ( .A(round_inst_aout_z[20]), .B(
        round_inst_srout_z[20]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[20]) );
  MUX2_X1 round_inst_mux_inv_z_U16 ( .A(round_inst_aout_z[16]), .B(
        round_inst_srout_z[16]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[16]) );
  MUX2_X1 round_inst_mux_inv_z_U15 ( .A(round_inst_aout_z[12]), .B(
        round_inst_srout_z[12]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[12]) );
  MUX2_X1 round_inst_mux_inv_z_U14 ( .A(round_inst_aout_z[13]), .B(
        round_inst_aout_z[12]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[13]) );
  MUX2_X1 round_inst_mux_inv_z_U13 ( .A(round_inst_aout_z[8]), .B(
        round_inst_srout_z[8]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[8]) );
  MUX2_X1 round_inst_mux_inv_z_U12 ( .A(round_inst_aout_z[4]), .B(
        round_inst_srout_z[4]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[4]) );
  MUX2_X1 round_inst_mux_inv_z_U11 ( .A(round_inst_aout_z[5]), .B(
        round_inst_aout_z[36]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[5]) );
  MUX2_X1 round_inst_mux_inv_z_U10 ( .A(round_inst_aout_z[0]), .B(
        round_inst_srout_z[0]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[0]) );
  MUX2_X1 round_inst_mux_inv_z_U9 ( .A(round_inst_aout_z[1]), .B(
        round_inst_aout_z[16]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[1]) );
  INV_X1 round_inst_mux_inv_z_U8 ( .A(round_inst_mux_inv_z_n263), .ZN(
        round_inst_mux_inv_z_n264) );
  INV_X1 round_inst_mux_inv_z_U7 ( .A(round_inst_mux_inv_z_n263), .ZN(
        round_inst_mux_inv_z_n265) );
  INV_X1 round_inst_mux_inv_z_U6 ( .A(inv_sig), .ZN(round_inst_mux_inv_z_n263)
         );
  MUX2_X2 round_inst_mux_inv_z_U5 ( .A(round_inst_aout_z[43]), .B(
        round_inst_aout_z[26]), .S(round_inst_mux_inv_z_n267), .Z(
        round_inst_sin_z[43]) );
  MUX2_X2 round_inst_mux_inv_z_U4 ( .A(round_inst_aout_z[15]), .B(
        round_inst_aout_z[14]), .S(round_inst_mux_inv_z_n264), .Z(
        round_inst_sin_z[15]) );
  MUX2_X2 round_inst_mux_inv_z_U3 ( .A(round_inst_aout_z[47]), .B(
        round_inst_aout_z[46]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[47]) );
  MUX2_X2 round_inst_mux_inv_z_U2 ( .A(round_inst_aout_z[55]), .B(
        round_inst_aout_z[22]), .S(round_inst_mux_inv_z_n266), .Z(
        round_inst_sin_z[55]) );
  MUX2_X2 round_inst_mux_inv_z_U1 ( .A(round_inst_aout_z[3]), .B(
        round_inst_aout_z[18]), .S(round_inst_mux_inv_z_n265), .Z(
        round_inst_sin_z[3]) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U149 ( .A(
        round_inst_sbox_inst0_com_w_inst_n160), .B(
        round_inst_sbox_inst0_com_w_inst_n159), .ZN(round_inst_sout_w[3]) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U148 ( .A(
        round_inst_sbox_inst0_com_w_inst_n158), .B(
        round_inst_sbox_inst0_com_w_inst_n157), .ZN(
        round_inst_sbox_inst0_com_w_inst_n159) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U147 ( .A(
        round_inst_sbox_inst0_com_w_inst_n156), .B(
        round_inst_sbox_inst0_com_w_inst_n155), .ZN(
        round_inst_sbox_inst0_com_w_inst_n157) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U146 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n154), .A2(round_inst_sin_z[0]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n155) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U145 ( .A(
        round_inst_sbox_inst0_com_w_inst_n153), .B(
        round_inst_sbox_inst0_com_w_inst_n152), .ZN(
        round_inst_sbox_inst0_com_w_inst_n156) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U144 ( .A(
        round_inst_sbox_inst0_com_w_inst_n151), .B(
        round_inst_sbox_inst0_com_w_inst_n150), .ZN(
        round_inst_sbox_inst0_com_w_inst_n152) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U143 ( .A(
        round_inst_sbox_inst0_com_w_inst_n149), .B(
        round_inst_sbox_inst0_com_w_inst_n148), .ZN(
        round_inst_sbox_inst0_com_w_inst_n150) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U142 ( .A(cin[3]), .B(din[3]), 
        .ZN(round_inst_sbox_inst0_com_w_inst_n148) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U141 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n147), .A2(
        round_inst_sbox_inst0_com_w_inst_n146), .ZN(
        round_inst_sbox_inst0_com_w_inst_n149) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U140 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n145), .A2(
        round_inst_sbox_inst0_com_w_inst_n144), .ZN(
        round_inst_sbox_inst0_com_w_inst_n147) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U139 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n143), .A2(
        round_inst_sbox_inst0_com_w_inst_n142), .ZN(
        round_inst_sbox_inst0_com_w_inst_n151) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U138 ( .A(
        round_inst_sbox_inst0_com_w_inst_n141), .B(
        round_inst_sbox_inst0_com_w_inst_n140), .ZN(
        round_inst_sbox_inst0_com_w_inst_n158) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U137 ( .A(
        round_inst_sbox_inst0_com_w_inst_n139), .B(
        round_inst_sbox_inst0_com_w_inst_n138), .ZN(
        round_inst_sbox_inst0_com_w_inst_n140) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U136 ( .A(
        round_inst_sbox_inst0_com_w_inst_n137), .B(
        round_inst_sbox_inst0_com_w_inst_n136), .Z(
        round_inst_sbox_inst0_com_w_inst_n138) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U135 ( .A(
        round_inst_sbox_inst0_com_w_inst_n135), .B(
        round_inst_sbox_inst0_com_w_inst_n134), .ZN(
        round_inst_sbox_inst0_com_w_inst_n136) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U134 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n133), .A2(round_inst_sin_z[2]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n134) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U133 ( .A(
        round_inst_sbox_inst0_com_w_inst_n132), .B(
        round_inst_sbox_inst0_com_w_inst_n131), .Z(
        round_inst_sbox_inst0_com_w_inst_n133) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U132 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n144), .A2(round_inst_n40), .ZN(
        round_inst_sbox_inst0_com_w_inst_n131) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U131 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n130), .A2(
        round_inst_sbox_inst0_com_w_inst_n129), .ZN(
        round_inst_sbox_inst0_com_w_inst_n135) );
  NAND3_X1 round_inst_sbox_inst0_com_w_inst_U130 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n144), .A2(round_inst_sin_y[2]), .A3(
        round_inst_sbox_inst0_com_w_inst_n128), .ZN(
        round_inst_sbox_inst0_com_w_inst_n137) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U129 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n127), .A2(
        round_inst_sbox_inst0_com_w_inst_n126), .ZN(
        round_inst_sbox_inst0_com_w_inst_n139) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U128 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n144), .A2(round_inst_sin_x[2]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n126) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U127 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n125), .A2(
        round_inst_sbox_inst0_com_w_inst_n124), .ZN(
        round_inst_sbox_inst0_com_w_inst_n141) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U126 ( .A(
        round_inst_sbox_inst0_com_w_inst_n123), .B(
        round_inst_sbox_inst0_com_w_inst_n143), .ZN(
        round_inst_sbox_inst0_com_w_inst_n125) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U125 ( .A1(round_inst_n40), .A2(
        round_inst_sin_x[2]), .ZN(round_inst_sbox_inst0_com_w_inst_n123) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U124 ( .A(
        round_inst_sbox_inst0_com_w_inst_n153), .B(
        round_inst_sbox_inst0_com_w_inst_n122), .ZN(round_inst_sout_w[1]) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U123 ( .A(
        round_inst_sbox_inst0_com_w_inst_n121), .B(
        round_inst_sbox_inst0_com_w_inst_n120), .ZN(
        round_inst_sbox_inst0_com_w_inst_n122) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U122 ( .A(
        round_inst_sbox_inst0_com_w_inst_n119), .B(
        round_inst_sbox_inst0_com_w_inst_n118), .ZN(
        round_inst_sbox_inst0_com_w_inst_n120) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U121 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n117), .A2(
        round_inst_sbox_inst0_com_w_inst_n124), .ZN(
        round_inst_sbox_inst0_com_w_inst_n119) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U120 ( .A(round_inst_sin_x[2]), 
        .B(round_inst_sin_z[2]), .ZN(round_inst_sbox_inst0_com_w_inst_n117) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U119 ( .A(
        round_inst_sbox_inst0_com_w_inst_n130), .B(
        round_inst_sbox_inst0_com_w_inst_n116), .ZN(
        round_inst_sbox_inst0_com_w_inst_n121) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U118 ( .A(
        round_inst_sbox_inst0_com_w_inst_n115), .B(
        round_inst_sbox_inst0_com_w_inst_n114), .ZN(
        round_inst_sbox_inst0_com_w_inst_n116) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U117 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n144), .A2(round_inst_sin_y[2]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n114) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U116 ( .A(din[1]), .B(cin[1]), 
        .ZN(round_inst_sbox_inst0_com_w_inst_n115) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U115 ( .A(
        round_inst_sbox_inst0_com_w_inst_n113), .B(
        round_inst_sbox_inst0_com_w_inst_n112), .ZN(round_inst_sout_w[0]) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U114 ( .A(
        round_inst_sbox_inst0_com_w_inst_n111), .B(
        round_inst_sbox_inst0_com_w_inst_n110), .ZN(
        round_inst_sbox_inst0_com_w_inst_n113) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U113 ( .A(
        round_inst_sbox_inst0_com_w_inst_n109), .B(
        round_inst_sbox_inst0_com_w_inst_n108), .ZN(
        round_inst_sbox_inst0_com_w_inst_n110) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U112 ( .A(round_inst_sin_x[2]), .B(
        round_inst_sbox_inst0_com_w_inst_n107), .Z(
        round_inst_sbox_inst0_com_w_inst_n108) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U111 ( .A(cin[0]), .B(din[0]), .Z(
        round_inst_sbox_inst0_com_w_inst_n109) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U110 ( .A(
        round_inst_sbox_inst0_com_w_inst_n153), .B(
        round_inst_sbox_inst0_com_w_inst_n154), .ZN(
        round_inst_sbox_inst0_com_w_inst_n111) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U109 ( .A(
        round_inst_sbox_inst0_com_w_inst_n106), .B(
        round_inst_sbox_inst0_com_w_inst_n143), .ZN(
        round_inst_sbox_inst0_com_w_inst_n154) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U108 ( .A(
        round_inst_sbox_inst0_com_w_inst_n105), .B(
        round_inst_sbox_inst0_com_w_inst_n104), .ZN(
        round_inst_sbox_inst0_com_w_inst_n106) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U107 ( .A(
        round_inst_sbox_inst0_com_w_inst_n103), .B(
        round_inst_sbox_inst0_com_w_inst_n102), .Z(
        round_inst_sbox_inst0_com_w_inst_n153) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U106 ( .A(
        round_inst_sbox_inst0_com_w_inst_n101), .B(
        round_inst_sbox_inst0_com_w_inst_n100), .ZN(
        round_inst_sbox_inst0_com_w_inst_n102) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U105 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n99), .A2(round_inst_sin_z[0]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n100) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U104 ( .A(
        round_inst_sbox_inst0_com_w_inst_n98), .B(
        round_inst_sbox_inst0_com_w_inst_n97), .ZN(
        round_inst_sbox_inst0_com_w_inst_n101) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U103 ( .A(
        round_inst_sbox_inst0_com_w_inst_n96), .B(
        round_inst_sbox_inst0_com_w_inst_n95), .ZN(
        round_inst_sbox_inst0_com_w_inst_n97) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U102 ( .A(
        round_inst_sbox_inst0_com_w_inst_n94), .B(
        round_inst_sbox_inst0_com_w_inst_n93), .Z(
        round_inst_sbox_inst0_com_w_inst_n95) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U101 ( .A1(round_inst_sin_y[2]), 
        .A2(round_inst_sbox_inst0_com_w_inst_n92), .ZN(
        round_inst_sbox_inst0_com_w_inst_n93) );
  MUX2_X1 round_inst_sbox_inst0_com_w_inst_U100 ( .A(
        round_inst_sbox_inst0_com_w_inst_n91), .B(
        round_inst_sbox_inst0_com_w_inst_n146), .S(
        round_inst_sbox_inst0_com_w_inst_n124), .Z(
        round_inst_sbox_inst0_com_w_inst_n92) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U99 ( .A1(round_inst_sin_z[2]), 
        .A2(round_inst_sbox_inst0_com_w_inst_n90), .ZN(
        round_inst_sbox_inst0_com_w_inst_n94) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U98 ( .A(
        round_inst_sbox_inst0_com_w_inst_n89), .B(
        round_inst_sbox_inst0_com_w_inst_n88), .ZN(
        round_inst_sbox_inst0_com_w_inst_n90) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U97 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n87), .A2(round_inst_sin_x[2]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n96) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U96 ( .A(
        round_inst_sbox_inst0_com_w_inst_n146), .B(
        round_inst_sbox_inst0_com_w_inst_n86), .Z(
        round_inst_sbox_inst0_com_w_inst_n87) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U95 ( .A(
        round_inst_sbox_inst0_com_w_inst_n85), .B(
        round_inst_sbox_inst0_com_w_inst_n84), .ZN(
        round_inst_sbox_inst0_com_w_inst_n86) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U94 ( .A1(round_inst_sin_y[0]), 
        .A2(round_inst_sin_z[1]), .ZN(round_inst_sbox_inst0_com_w_inst_n84) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U93 ( .A(
        round_inst_sbox_inst0_com_w_inst_n83), .B(
        round_inst_sbox_inst0_com_w_inst_n88), .ZN(
        round_inst_sbox_inst0_com_w_inst_n85) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U92 ( .A(
        round_inst_sbox_inst0_com_w_inst_n82), .B(
        round_inst_sbox_inst0_com_w_inst_n81), .Z(
        round_inst_sbox_inst0_com_w_inst_n98) );
  NAND3_X1 round_inst_sbox_inst0_com_w_inst_U91 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n146), .A2(round_inst_sin_z[2]), .A3(
        round_inst_sbox_inst0_com_w_inst_n142), .ZN(
        round_inst_sbox_inst0_com_w_inst_n81) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U90 ( .A(round_inst_sin_y[0]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n142) );
  NAND3_X1 round_inst_sbox_inst0_com_w_inst_U89 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n144), .A2(round_inst_sin_z[1]), .A3(
        round_inst_sin_y[2]), .ZN(round_inst_sbox_inst0_com_w_inst_n82) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U88 ( .A(
        round_inst_sbox_inst0_com_w_inst_n80), .B(
        round_inst_sbox_inst0_com_w_inst_n79), .Z(
        round_inst_sbox_inst0_com_w_inst_n103) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U87 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n78), .A2(
        round_inst_sbox_inst0_com_w_inst_n91), .ZN(
        round_inst_sbox_inst0_com_w_inst_n79) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U86 ( .A(
        round_inst_sbox_inst0_com_w_inst_n130), .B(
        round_inst_sbox_inst0_com_w_inst_n77), .Z(
        round_inst_sbox_inst0_com_w_inst_n78) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U85 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n144), .A2(round_inst_sin_z[2]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n77) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U84 ( .A1(round_inst_sin_y[0]), 
        .A2(round_inst_sin_x[2]), .ZN(round_inst_sbox_inst0_com_w_inst_n130)
         );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U83 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n76), .A2(round_inst_sin_y[2]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n80) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U82 ( .A(
        round_inst_sbox_inst0_com_w_inst_n75), .B(
        round_inst_sbox_inst0_com_w_inst_n88), .Z(
        round_inst_sbox_inst0_com_w_inst_n76) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U81 ( .A(
        round_inst_sbox_inst0_com_w_inst_n74), .B(
        round_inst_sbox_inst0_com_w_inst_n112), .Z(round_inst_xin_w[3]) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U80 ( .A(
        round_inst_sbox_inst0_com_w_inst_n73), .B(
        round_inst_sbox_inst0_com_w_inst_n72), .ZN(
        round_inst_sbox_inst0_com_w_inst_n112) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U79 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n71), .A2(
        round_inst_sbox_inst0_com_w_inst_n144), .ZN(
        round_inst_sbox_inst0_com_w_inst_n72) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U78 ( .A(
        round_inst_sbox_inst0_com_w_inst_n70), .B(
        round_inst_sbox_inst0_com_w_inst_n69), .ZN(
        round_inst_sbox_inst0_com_w_inst_n71) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U77 ( .A(
        round_inst_sbox_inst0_com_w_inst_n129), .B(
        round_inst_sbox_inst0_com_w_inst_n68), .Z(
        round_inst_sbox_inst0_com_w_inst_n70) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U76 ( .A(
        round_inst_sbox_inst0_com_w_inst_n67), .B(
        round_inst_sbox_inst0_com_w_inst_n145), .Z(
        round_inst_sbox_inst0_com_w_inst_n129) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U75 ( .A(
        round_inst_sbox_inst0_com_w_inst_n75), .B(
        round_inst_sbox_inst0_com_w_inst_n132), .ZN(
        round_inst_sbox_inst0_com_w_inst_n73) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U74 ( .A(
        round_inst_sbox_inst0_com_w_inst_n66), .B(
        round_inst_sbox_inst0_com_w_inst_n65), .ZN(
        round_inst_sbox_inst0_com_w_inst_n74) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U73 ( .A(
        round_inst_sbox_inst0_com_w_inst_n160), .B(
        round_inst_sbox_inst0_com_w_inst_n118), .ZN(
        round_inst_sbox_inst0_com_w_inst_n65) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U72 ( .A(
        round_inst_sbox_inst0_com_w_inst_n64), .B(
        round_inst_sbox_inst0_com_w_inst_n63), .Z(
        round_inst_sbox_inst0_com_w_inst_n118) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U71 ( .A(
        round_inst_sbox_inst0_com_w_inst_n62), .B(
        round_inst_sbox_inst0_com_w_inst_n61), .ZN(
        round_inst_sbox_inst0_com_w_inst_n63) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U70 ( .A(
        round_inst_sbox_inst0_com_w_inst_n60), .B(
        round_inst_sbox_inst0_com_w_inst_n59), .ZN(
        round_inst_sbox_inst0_com_w_inst_n61) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U69 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n69), .A2(
        round_inst_sbox_inst0_com_w_inst_n143), .ZN(
        round_inst_sbox_inst0_com_w_inst_n59) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U68 ( .A1(round_inst_sin_y[2]), 
        .A2(round_inst_sbox_inst0_com_w_inst_n145), .ZN(
        round_inst_sbox_inst0_com_w_inst_n143) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U67 ( .A(
        round_inst_sbox_inst0_com_w_inst_n58), .B(round_inst_sin_z[1]), .Z(
        round_inst_sbox_inst0_com_w_inst_n69) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U66 ( .A(
        round_inst_sbox_inst0_com_w_inst_n57), .B(
        round_inst_sbox_inst0_com_w_inst_n56), .ZN(
        round_inst_sbox_inst0_com_w_inst_n60) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U65 ( .A(
        round_inst_sbox_inst0_com_w_inst_n55), .B(
        round_inst_sbox_inst0_com_w_inst_n54), .ZN(
        round_inst_sbox_inst0_com_w_inst_n56) );
  NOR3_X1 round_inst_sbox_inst0_com_w_inst_U64 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n68), .A2(
        round_inst_sbox_inst0_com_w_inst_n53), .A3(
        round_inst_sbox_inst0_com_w_inst_n67), .ZN(
        round_inst_sbox_inst0_com_w_inst_n54) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U63 ( .A(round_inst_sin_x[2]), .B(
        round_inst_sin_y[2]), .ZN(round_inst_sbox_inst0_com_w_inst_n53) );
  NAND3_X1 round_inst_sbox_inst0_com_w_inst_U62 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n146), .A2(round_inst_n40), .A3(
        round_inst_sin_z[2]), .ZN(round_inst_sbox_inst0_com_w_inst_n55) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U61 ( .A(
        round_inst_sbox_inst0_com_w_inst_n52), .B(
        round_inst_sbox_inst0_com_w_inst_n51), .ZN(
        round_inst_sbox_inst0_com_w_inst_n57) );
  NOR3_X1 round_inst_sbox_inst0_com_w_inst_U60 ( .A1(round_inst_sin_z[2]), 
        .A2(round_inst_sbox_inst0_com_w_inst_n107), .A3(
        round_inst_sbox_inst0_com_w_inst_n58), .ZN(
        round_inst_sbox_inst0_com_w_inst_n51) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U59 ( .A(
        round_inst_sbox_inst0_com_w_inst_n50), .B(
        round_inst_sbox_inst0_com_w_inst_n49), .ZN(
        round_inst_sbox_inst0_com_w_inst_n52) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U58 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n105), .A2(
        round_inst_sbox_inst0_com_w_inst_n48), .ZN(
        round_inst_sbox_inst0_com_w_inst_n49) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U57 ( .A1(round_inst_sin_x[2]), 
        .A2(round_inst_sbox_inst0_com_w_inst_n128), .ZN(
        round_inst_sbox_inst0_com_w_inst_n105) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U56 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n99), .A2(
        round_inst_sbox_inst0_com_w_inst_n47), .ZN(
        round_inst_sbox_inst0_com_w_inst_n50) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U55 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n91), .A2(round_inst_sin_x[2]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n99) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U54 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n46), .A2(
        round_inst_sbox_inst0_com_w_inst_n146), .ZN(
        round_inst_sbox_inst0_com_w_inst_n62) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U53 ( .A(
        round_inst_sbox_inst0_com_w_inst_n128), .B(
        round_inst_sbox_inst0_com_w_inst_n45), .Z(
        round_inst_sbox_inst0_com_w_inst_n46) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U52 ( .A1(round_inst_sin_y[2]), 
        .A2(round_inst_sbox_inst0_com_w_inst_n107), .ZN(
        round_inst_sbox_inst0_com_w_inst_n45) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U51 ( .A(
        round_inst_sbox_inst0_com_w_inst_n67), .ZN(
        round_inst_sbox_inst0_com_w_inst_n128) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U50 ( .A(
        round_inst_sbox_inst0_com_w_inst_n44), .B(
        round_inst_sbox_inst0_com_w_inst_n43), .Z(
        round_inst_sbox_inst0_com_w_inst_n64) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U49 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n104), .A2(
        round_inst_sbox_inst0_com_w_inst_n42), .ZN(
        round_inst_sbox_inst0_com_w_inst_n43) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U48 ( .A(round_inst_sin_z[1]), .B(
        round_inst_sbox_inst0_com_w_inst_n146), .ZN(
        round_inst_sbox_inst0_com_w_inst_n42) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U47 ( .A1(round_inst_sin_x[2]), 
        .A2(round_inst_sbox_inst0_com_w_inst_n145), .ZN(
        round_inst_sbox_inst0_com_w_inst_n104) );
  NAND3_X1 round_inst_sbox_inst0_com_w_inst_U46 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n41), .A2(round_inst_sin_x[2]), .A3(
        round_inst_sbox_inst0_com_w_inst_n91), .ZN(
        round_inst_sbox_inst0_com_w_inst_n44) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U45 ( .A(round_inst_n40), .B(
        round_inst_sbox_inst0_com_w_inst_n107), .ZN(
        round_inst_sbox_inst0_com_w_inst_n41) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U44 ( .A(
        round_inst_sbox_inst0_com_w_inst_n40), .B(
        round_inst_sbox_inst0_com_w_inst_n39), .ZN(
        round_inst_sbox_inst0_com_w_inst_n160) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U43 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n38), .A2(round_inst_n40), .ZN(
        round_inst_sbox_inst0_com_w_inst_n39) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U42 ( .A(
        round_inst_sbox_inst0_com_w_inst_n83), .B(
        round_inst_sbox_inst0_com_w_inst_n37), .ZN(
        round_inst_sbox_inst0_com_w_inst_n38) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U41 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n144), .A2(round_inst_sin_z[1]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n37) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U40 ( .A(
        round_inst_sbox_inst0_com_w_inst_n36), .B(
        round_inst_sbox_inst0_com_w_inst_n75), .ZN(
        round_inst_sbox_inst0_com_w_inst_n83) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U39 ( .A(
        round_inst_sbox_inst0_com_w_inst_n35), .B(
        round_inst_sbox_inst0_com_w_inst_n89), .ZN(
        round_inst_sbox_inst0_com_w_inst_n36) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U38 ( .A(
        round_inst_sbox_inst0_com_w_inst_n34), .B(
        round_inst_sbox_inst0_com_w_inst_n33), .ZN(
        round_inst_sbox_inst0_com_w_inst_n40) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U37 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n32), .A2(
        round_inst_sbox_inst0_com_w_inst_n91), .ZN(
        round_inst_sbox_inst0_com_w_inst_n33) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U36 ( .A(
        round_inst_sbox_inst0_com_w_inst_n132), .B(
        round_inst_sbox_inst0_com_w_inst_n31), .Z(
        round_inst_sbox_inst0_com_w_inst_n32) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U35 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n144), .A2(round_inst_sin_z[3]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n31) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U34 ( .A(
        round_inst_sbox_inst0_com_w_inst_n30), .B(
        round_inst_sbox_inst0_com_w_inst_n29), .ZN(
        round_inst_sbox_inst0_com_w_inst_n34) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U33 ( .A(
        round_inst_sbox_inst0_com_w_inst_n28), .B(
        round_inst_sbox_inst0_com_w_inst_n27), .ZN(
        round_inst_sbox_inst0_com_w_inst_n29) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U32 ( .A(
        round_inst_sbox_inst0_com_w_inst_n26), .B(
        round_inst_sbox_inst0_com_w_inst_n25), .ZN(
        round_inst_sbox_inst0_com_w_inst_n27) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U31 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n127), .A2(
        round_inst_sbox_inst0_com_w_inst_n75), .ZN(
        round_inst_sbox_inst0_com_w_inst_n25) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U30 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n146), .A2(round_inst_sin_y[0]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n75) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U29 ( .A(
        round_inst_sbox_inst0_com_w_inst_n47), .B(
        round_inst_sbox_inst0_com_w_inst_n145), .Z(
        round_inst_sbox_inst0_com_w_inst_n127) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U28 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n48), .A2(
        round_inst_sbox_inst0_com_w_inst_n132), .ZN(
        round_inst_sbox_inst0_com_w_inst_n26) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U27 ( .A1(round_inst_sin_y[0]), 
        .A2(round_inst_sbox_inst0_com_w_inst_n145), .ZN(
        round_inst_sbox_inst0_com_w_inst_n132) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U26 ( .A(round_inst_sin_z[1]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n48) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U25 ( .A(
        round_inst_sbox_inst0_com_w_inst_n24), .B(
        round_inst_sbox_inst0_com_w_inst_n23), .ZN(
        round_inst_sbox_inst0_com_w_inst_n28) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U24 ( .A(
        round_inst_sbox_inst0_com_w_inst_n22), .B(
        round_inst_sbox_inst0_com_w_inst_n21), .Z(
        round_inst_sbox_inst0_com_w_inst_n23) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U23 ( .A1(round_inst_sin_z[3]), 
        .A2(round_inst_sbox_inst0_com_w_inst_n89), .ZN(
        round_inst_sbox_inst0_com_w_inst_n21) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U22 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n68), .A2(
        round_inst_sbox_inst0_com_w_inst_n124), .ZN(
        round_inst_sbox_inst0_com_w_inst_n89) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U21 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n88), .A2(
        round_inst_sbox_inst0_com_w_inst_n67), .ZN(
        round_inst_sbox_inst0_com_w_inst_n22) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U20 ( .A(round_inst_n40), .B(
        round_inst_sbox_inst0_com_w_inst_n47), .Z(
        round_inst_sbox_inst0_com_w_inst_n67) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U19 ( .A(round_inst_sin_z[3]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n47) );
  NOR2_X1 round_inst_sbox_inst0_com_w_inst_U18 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n107), .A2(
        round_inst_sbox_inst0_com_w_inst_n35), .ZN(
        round_inst_sbox_inst0_com_w_inst_n24) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U17 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n91), .A2(
        round_inst_sbox_inst0_com_w_inst_n144), .ZN(
        round_inst_sbox_inst0_com_w_inst_n35) );
  NAND3_X1 round_inst_sbox_inst0_com_w_inst_U16 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n20), .A2(
        round_inst_sbox_inst0_com_w_inst_n19), .A3(
        round_inst_sbox_inst0_com_w_inst_n145), .ZN(
        round_inst_sbox_inst0_com_w_inst_n30) );
  NAND3_X1 round_inst_sbox_inst0_com_w_inst_U15 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n91), .A2(round_inst_sin_z[0]), .A3(
        round_inst_sbox_inst0_com_w_inst_n68), .ZN(
        round_inst_sbox_inst0_com_w_inst_n19) );
  OR2_X1 round_inst_sbox_inst0_com_w_inst_U14 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n88), .A2(
        round_inst_sbox_inst0_com_w_inst_n91), .ZN(
        round_inst_sbox_inst0_com_w_inst_n20) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U13 ( .A(
        round_inst_sbox_inst0_com_w_inst_n58), .ZN(
        round_inst_sbox_inst0_com_w_inst_n91) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U12 ( .A(round_inst_sin_y[1]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n58) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U11 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n146), .A2(round_inst_sin_z[0]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n88) );
  XOR2_X1 round_inst_sbox_inst0_com_w_inst_U10 ( .A(
        round_inst_sbox_inst0_com_w_inst_n18), .B(cin[2]), .Z(
        round_inst_sbox_inst0_com_w_inst_n66) );
  XNOR2_X1 round_inst_sbox_inst0_com_w_inst_U9 ( .A(
        round_inst_sbox_inst0_com_w_inst_n17), .B(din[2]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n18) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U8 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n16), .A2(
        round_inst_sbox_inst0_com_w_inst_n144), .ZN(
        round_inst_sbox_inst0_com_w_inst_n17) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U7 ( .A(
        round_inst_sbox_inst0_com_w_inst_n124), .ZN(
        round_inst_sbox_inst0_com_w_inst_n144) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U6 ( .A(round_inst_sin_x[0]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n124) );
  NAND2_X1 round_inst_sbox_inst0_com_w_inst_U5 ( .A1(
        round_inst_sbox_inst0_com_w_inst_n145), .A2(
        round_inst_sbox_inst0_com_w_inst_n146), .ZN(
        round_inst_sbox_inst0_com_w_inst_n16) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U4 ( .A(
        round_inst_sbox_inst0_com_w_inst_n68), .ZN(
        round_inst_sbox_inst0_com_w_inst_n146) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U3 ( .A(round_inst_sin_x[1]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n68) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U2 ( .A(
        round_inst_sbox_inst0_com_w_inst_n107), .ZN(
        round_inst_sbox_inst0_com_w_inst_n145) );
  INV_X1 round_inst_sbox_inst0_com_w_inst_U1 ( .A(round_inst_sin_x[3]), .ZN(
        round_inst_sbox_inst0_com_w_inst_n107) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U145 ( .A(
        round_inst_sbox_inst0_com_x_inst_n299), .B(
        round_inst_sbox_inst0_com_x_inst_n298), .ZN(round_inst_sout_x[0]) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U144 ( .A(
        round_inst_sbox_inst0_com_x_inst_n297), .B(
        round_inst_sbox_inst0_com_x_inst_n296), .ZN(
        round_inst_sbox_inst0_com_x_inst_n299) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U143 ( .A(round_inst_n40), .B(
        round_inst_sbox_inst0_com_x_inst_n295), .ZN(
        round_inst_sbox_inst0_com_x_inst_n296) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U142 ( .A(din[0]), .B(
        round_inst_sbox_inst0_com_x_inst_n294), .Z(
        round_inst_sbox_inst0_com_x_inst_n297) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U141 ( .A(
        round_inst_sbox_inst0_com_x_inst_n293), .B(
        round_inst_sbox_inst0_com_x_inst_n292), .ZN(round_inst_srout2_x[18])
         );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U140 ( .A(
        round_inst_sbox_inst0_com_x_inst_n291), .B(
        round_inst_sbox_inst0_com_x_inst_n294), .ZN(
        round_inst_sbox_inst0_com_x_inst_n292) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U139 ( .A(
        round_inst_sbox_inst0_com_x_inst_n290), .B(
        round_inst_sbox_inst0_com_x_inst_n289), .ZN(
        round_inst_sbox_inst0_com_x_inst_n294) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U138 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n288), .A2(
        round_inst_sbox_inst0_com_x_inst_n287), .ZN(
        round_inst_sbox_inst0_com_x_inst_n289) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U137 ( .A(
        round_inst_sbox_inst0_com_x_inst_n286), .B(
        round_inst_sbox_inst0_com_x_inst_n285), .ZN(
        round_inst_sbox_inst0_com_x_inst_n290) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U136 ( .A(
        round_inst_sbox_inst0_com_x_inst_n284), .B(
        round_inst_sbox_inst0_com_x_inst_n283), .Z(
        round_inst_sbox_inst0_com_x_inst_n293) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U135 ( .A(
        round_inst_sbox_inst0_com_x_inst_n282), .B(
        round_inst_sbox_inst0_com_x_inst_n281), .ZN(
        round_inst_sbox_inst0_com_x_inst_n283) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U134 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n286), .A2(round_inst_sin_z[0]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n281) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U133 ( .A(
        round_inst_sbox_inst0_com_x_inst_n280), .B(
        round_inst_sbox_inst0_com_x_inst_n279), .Z(
        round_inst_sbox_inst0_com_x_inst_n282) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U132 ( .A(
        round_inst_sbox_inst0_com_x_inst_n278), .B(
        round_inst_sbox_inst0_com_x_inst_n277), .Z(
        round_inst_sbox_inst0_com_x_inst_n279) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U131 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n276), .A2(
        round_inst_sbox_inst0_com_x_inst_n275), .ZN(
        round_inst_sbox_inst0_com_x_inst_n277) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U130 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n274), .A2(
        round_inst_sbox_inst0_com_x_inst_n287), .ZN(
        round_inst_sbox_inst0_com_x_inst_n278) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U129 ( .A(
        round_inst_sbox_inst0_com_x_inst_n273), .B(
        round_inst_sbox_inst0_com_x_inst_n272), .ZN(
        round_inst_sbox_inst0_com_x_inst_n280) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U128 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n271), .A2(
        round_inst_sbox_inst0_com_x_inst_n270), .ZN(
        round_inst_sbox_inst0_com_x_inst_n272) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U127 ( .A(round_inst_sin_y[1]), 
        .B(din[3]), .ZN(round_inst_sbox_inst0_com_x_inst_n273) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U126 ( .A(
        round_inst_sbox_inst0_com_x_inst_n269), .B(
        round_inst_sbox_inst0_com_x_inst_n268), .ZN(
        round_inst_sbox_inst0_com_x_inst_n284) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U125 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n267), .A2(round_inst_sin_z[3]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n268) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U124 ( .A(
        round_inst_sbox_inst0_com_x_inst_n274), .B(
        round_inst_sbox_inst0_com_x_inst_n266), .Z(
        round_inst_sbox_inst0_com_x_inst_n267) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U123 ( .A1(round_inst_sin_w[0]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n295), .ZN(
        round_inst_sbox_inst0_com_x_inst_n266) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U122 ( .A(
        round_inst_sbox_inst0_com_x_inst_n265), .B(
        round_inst_sbox_inst0_com_x_inst_n264), .ZN(
        round_inst_sbox_inst0_com_x_inst_n269) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U121 ( .A(
        round_inst_sbox_inst0_com_x_inst_n263), .B(
        round_inst_sbox_inst0_com_x_inst_n262), .ZN(
        round_inst_sbox_inst0_com_x_inst_n264) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U120 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n261), .A2(
        round_inst_sbox_inst0_com_x_inst_n270), .ZN(
        round_inst_sbox_inst0_com_x_inst_n262) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U119 ( .A(
        round_inst_sbox_inst0_com_x_inst_n260), .B(
        round_inst_sbox_inst0_com_x_inst_n259), .ZN(
        round_inst_sbox_inst0_com_x_inst_n263) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U118 ( .A(
        round_inst_sbox_inst0_com_x_inst_n258), .B(
        round_inst_sbox_inst0_com_x_inst_n257), .Z(
        round_inst_sbox_inst0_com_x_inst_n259) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U117 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n275), .A2(
        round_inst_sbox_inst0_com_x_inst_n261), .ZN(
        round_inst_sbox_inst0_com_x_inst_n257) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U116 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n276), .A2(
        round_inst_sbox_inst0_com_x_inst_n270), .ZN(
        round_inst_sbox_inst0_com_x_inst_n258) );
  INV_X1 round_inst_sbox_inst0_com_x_inst_U115 ( .A(round_inst_sin_w[3]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n270) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U114 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n256), .A2(
        round_inst_sbox_inst0_com_x_inst_n255), .ZN(
        round_inst_sbox_inst0_com_x_inst_n260) );
  INV_X1 round_inst_sbox_inst0_com_x_inst_U113 ( .A(round_inst_sin_w[0]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n256) );
  NAND3_X1 round_inst_sbox_inst0_com_x_inst_U112 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n254), .A2(round_inst_sin_z[0]), .A3(
        round_inst_n40), .ZN(round_inst_sbox_inst0_com_x_inst_n265) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U111 ( .A(round_inst_sin_w[2]), .B(
        round_inst_sbox_inst0_com_x_inst_n295), .Z(
        round_inst_sbox_inst0_com_x_inst_n254) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U110 ( .A(
        round_inst_sbox_inst0_com_x_inst_n253), .B(
        round_inst_sbox_inst0_com_x_inst_n276), .ZN(round_inst_srout2_x[16])
         );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U109 ( .A1(round_inst_sin_y[0]), 
        .A2(round_inst_sin_z[2]), .ZN(round_inst_sbox_inst0_com_x_inst_n276)
         );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U108 ( .A(
        round_inst_sbox_inst0_com_x_inst_n252), .B(
        round_inst_sbox_inst0_com_x_inst_n251), .Z(
        round_inst_sbox_inst0_com_x_inst_n253) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U107 ( .A(
        round_inst_sbox_inst0_com_x_inst_n250), .B(
        round_inst_sbox_inst0_com_x_inst_n249), .ZN(
        round_inst_sbox_inst0_com_x_inst_n252) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U106 ( .A(
        round_inst_sbox_inst0_com_x_inst_n248), .B(
        round_inst_sbox_inst0_com_x_inst_n285), .ZN(
        round_inst_sbox_inst0_com_x_inst_n249) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U105 ( .A(
        round_inst_sbox_inst0_com_x_inst_n247), .B(
        round_inst_sbox_inst0_com_x_inst_n246), .ZN(
        round_inst_sbox_inst0_com_x_inst_n285) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U104 ( .A1(round_inst_sin_z[2]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n245), .ZN(
        round_inst_sbox_inst0_com_x_inst_n246) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U103 ( .A(
        round_inst_sbox_inst0_com_x_inst_n244), .B(
        round_inst_sbox_inst0_com_x_inst_n243), .Z(
        round_inst_sbox_inst0_com_x_inst_n247) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U102 ( .A(
        round_inst_sbox_inst0_com_x_inst_n242), .B(
        round_inst_sbox_inst0_com_x_inst_n241), .ZN(
        round_inst_sbox_inst0_com_x_inst_n243) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U101 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n295), .A2(
        round_inst_sbox_inst0_com_x_inst_n245), .ZN(
        round_inst_sbox_inst0_com_x_inst_n241) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U100 ( .A(
        round_inst_sbox_inst0_com_x_inst_n240), .B(
        round_inst_sbox_inst0_com_x_inst_n239), .ZN(
        round_inst_sbox_inst0_com_x_inst_n242) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U99 ( .A(
        round_inst_sbox_inst0_com_x_inst_n238), .B(
        round_inst_sbox_inst0_com_x_inst_n237), .ZN(
        round_inst_sbox_inst0_com_x_inst_n239) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U98 ( .A1(round_inst_sin_z[2]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n236), .ZN(
        round_inst_sbox_inst0_com_x_inst_n237) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U97 ( .A(
        round_inst_sbox_inst0_com_x_inst_n235), .B(
        round_inst_sbox_inst0_com_x_inst_n234), .Z(
        round_inst_sbox_inst0_com_x_inst_n238) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U96 ( .A(
        round_inst_sbox_inst0_com_x_inst_n233), .B(
        round_inst_sbox_inst0_com_x_inst_n232), .ZN(
        round_inst_sbox_inst0_com_x_inst_n234) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U95 ( .A1(round_inst_sin_z[2]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n231), .ZN(
        round_inst_sbox_inst0_com_x_inst_n232) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U94 ( .A(
        round_inst_sbox_inst0_com_x_inst_n230), .B(
        round_inst_sbox_inst0_com_x_inst_n229), .ZN(
        round_inst_sbox_inst0_com_x_inst_n231) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U93 ( .A1(round_inst_sin_w[0]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n228), .ZN(
        round_inst_sbox_inst0_com_x_inst_n230) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U92 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n227), .A2(
        round_inst_sbox_inst0_com_x_inst_n226), .ZN(
        round_inst_sbox_inst0_com_x_inst_n233) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U91 ( .A(round_inst_sin_z[0]), .B(
        round_inst_sin_w[0]), .Z(round_inst_sbox_inst0_com_x_inst_n226) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U90 ( .A1(round_inst_sin_z[1]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n295), .ZN(
        round_inst_sbox_inst0_com_x_inst_n227) );
  NOR3_X1 round_inst_sbox_inst0_com_x_inst_U89 ( .A1(round_inst_sin_z[0]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n225), .A3(
        round_inst_sbox_inst0_com_x_inst_n228), .ZN(
        round_inst_sbox_inst0_com_x_inst_n235) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U88 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n224), .A2(round_inst_sin_w[2]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n240) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U87 ( .A(
        round_inst_sbox_inst0_com_x_inst_n223), .B(
        round_inst_sbox_inst0_com_x_inst_n222), .Z(
        round_inst_sbox_inst0_com_x_inst_n224) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U86 ( .A(
        round_inst_sbox_inst0_com_x_inst_n229), .B(
        round_inst_sbox_inst0_com_x_inst_n245), .ZN(
        round_inst_sbox_inst0_com_x_inst_n223) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U85 ( .A(
        round_inst_sbox_inst0_com_x_inst_n221), .B(
        round_inst_sbox_inst0_com_x_inst_n220), .Z(
        round_inst_sbox_inst0_com_x_inst_n244) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U84 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n251), .A2(round_inst_n70), .ZN(
        round_inst_sbox_inst0_com_x_inst_n220) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U83 ( .A(
        round_inst_sbox_inst0_com_x_inst_n271), .B(
        round_inst_sbox_inst0_com_x_inst_n261), .Z(
        round_inst_sbox_inst0_com_x_inst_n251) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U82 ( .A1(round_inst_sin_y[0]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n295), .ZN(
        round_inst_sbox_inst0_com_x_inst_n261) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U81 ( .A1(round_inst_sin_z[0]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n295), .ZN(
        round_inst_sbox_inst0_com_x_inst_n271) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U80 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n295), .A2(
        round_inst_sbox_inst0_com_x_inst_n222), .ZN(
        round_inst_sbox_inst0_com_x_inst_n221) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U79 ( .A(
        round_inst_sbox_inst0_com_x_inst_n274), .B(din[1]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n250) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U78 ( .A1(round_inst_sin_y[0]), 
        .A2(round_inst_sin_w[2]), .ZN(round_inst_sbox_inst0_com_x_inst_n274)
         );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U77 ( .A(
        round_inst_sbox_inst0_com_x_inst_n219), .B(
        round_inst_sbox_inst0_com_x_inst_n298), .ZN(round_inst_srout2_x[19])
         );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U76 ( .A(
        round_inst_sbox_inst0_com_x_inst_n218), .B(
        round_inst_sbox_inst0_com_x_inst_n217), .ZN(
        round_inst_sbox_inst0_com_x_inst_n298) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U75 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n216), .A2(round_inst_sin_y[0]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n217) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U74 ( .A(
        round_inst_sbox_inst0_com_x_inst_n215), .B(
        round_inst_sbox_inst0_com_x_inst_n214), .ZN(
        round_inst_sbox_inst0_com_x_inst_n216) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U73 ( .A(round_inst_sin_z[1]), .B(
        round_inst_sin_y[1]), .ZN(round_inst_sbox_inst0_com_x_inst_n215) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U72 ( .A(
        round_inst_sbox_inst0_com_x_inst_n213), .B(
        round_inst_sbox_inst0_com_x_inst_n212), .ZN(
        round_inst_sbox_inst0_com_x_inst_n218) );
  INV_X1 round_inst_sbox_inst0_com_x_inst_U71 ( .A(
        round_inst_sbox_inst0_com_x_inst_n211), .ZN(
        round_inst_sbox_inst0_com_x_inst_n212) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U70 ( .A1(round_inst_n40), .A2(
        round_inst_sin_z[0]), .ZN(round_inst_sbox_inst0_com_x_inst_n213) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U69 ( .A(
        round_inst_sbox_inst0_com_x_inst_n210), .B(
        round_inst_sbox_inst0_com_x_inst_n209), .ZN(
        round_inst_sbox_inst0_com_x_inst_n219) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U68 ( .A(round_inst_sin_y[0]), .B(
        round_inst_sbox_inst0_com_x_inst_n291), .ZN(
        round_inst_sbox_inst0_com_x_inst_n209) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U67 ( .A(
        round_inst_sbox_inst0_com_x_inst_n208), .B(
        round_inst_sbox_inst0_com_x_inst_n207), .ZN(
        round_inst_sbox_inst0_com_x_inst_n291) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U66 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n236), .A2(round_inst_sin_z[3]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n207) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U65 ( .A(
        round_inst_sbox_inst0_com_x_inst_n206), .B(
        round_inst_sbox_inst0_com_x_inst_n222), .ZN(
        round_inst_sbox_inst0_com_x_inst_n236) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U64 ( .A(
        round_inst_sbox_inst0_com_x_inst_n205), .B(
        round_inst_sbox_inst0_com_x_inst_n204), .Z(
        round_inst_sbox_inst0_com_x_inst_n208) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U63 ( .A(
        round_inst_sbox_inst0_com_x_inst_n203), .B(
        round_inst_sbox_inst0_com_x_inst_n202), .ZN(
        round_inst_sbox_inst0_com_x_inst_n204) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U62 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n201), .A2(round_inst_sin_w[3]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n202) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U61 ( .A(
        round_inst_sbox_inst0_com_x_inst_n200), .B(
        round_inst_sbox_inst0_com_x_inst_n206), .Z(
        round_inst_sbox_inst0_com_x_inst_n201) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U60 ( .A(
        round_inst_sbox_inst0_com_x_inst_n199), .B(
        round_inst_sbox_inst0_com_x_inst_n198), .ZN(
        round_inst_sbox_inst0_com_x_inst_n203) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U59 ( .A(
        round_inst_sbox_inst0_com_x_inst_n197), .B(
        round_inst_sbox_inst0_com_x_inst_n196), .ZN(
        round_inst_sbox_inst0_com_x_inst_n198) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U58 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n222), .A2(round_inst_sin_w[3]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n196) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U57 ( .A(
        round_inst_sbox_inst0_com_x_inst_n195), .B(
        round_inst_sbox_inst0_com_x_inst_n194), .ZN(
        round_inst_sbox_inst0_com_x_inst_n197) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U56 ( .A(
        round_inst_sbox_inst0_com_x_inst_n193), .B(
        round_inst_sbox_inst0_com_x_inst_n192), .ZN(
        round_inst_sbox_inst0_com_x_inst_n194) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U55 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n191), .A2(round_inst_sin_z[3]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n192) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U54 ( .A(
        round_inst_sbox_inst0_com_x_inst_n245), .B(
        round_inst_sbox_inst0_com_x_inst_n190), .ZN(
        round_inst_sbox_inst0_com_x_inst_n191) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U53 ( .A1(round_inst_sin_y[1]), 
        .A2(round_inst_sin_w[0]), .ZN(round_inst_sbox_inst0_com_x_inst_n190)
         );
  INV_X1 round_inst_sbox_inst0_com_x_inst_U52 ( .A(
        round_inst_sbox_inst0_com_x_inst_n200), .ZN(
        round_inst_sbox_inst0_com_x_inst_n245) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U51 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n189), .A2(
        round_inst_sbox_inst0_com_x_inst_n188), .ZN(
        round_inst_sbox_inst0_com_x_inst_n193) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U50 ( .A(round_inst_sin_w[0]), .B(
        round_inst_sin_z[0]), .ZN(round_inst_sbox_inst0_com_x_inst_n189) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U49 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n187), .A2(round_inst_n40), .ZN(
        round_inst_sbox_inst0_com_x_inst_n195) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U48 ( .A(
        round_inst_sbox_inst0_com_x_inst_n211), .B(
        round_inst_sbox_inst0_com_x_inst_n200), .ZN(
        round_inst_sbox_inst0_com_x_inst_n187) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U47 ( .A1(round_inst_sin_y[0]), 
        .A2(round_inst_sin_z[1]), .ZN(round_inst_sbox_inst0_com_x_inst_n200)
         );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U46 ( .A(
        round_inst_sbox_inst0_com_x_inst_n229), .B(
        round_inst_sbox_inst0_com_x_inst_n206), .Z(
        round_inst_sbox_inst0_com_x_inst_n211) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U45 ( .A1(round_inst_sin_y[1]), 
        .A2(round_inst_sin_z[0]), .ZN(round_inst_sbox_inst0_com_x_inst_n206)
         );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U44 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n186), .A2(round_inst_n40), .ZN(
        round_inst_sbox_inst0_com_x_inst_n199) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U43 ( .A(
        round_inst_sbox_inst0_com_x_inst_n222), .B(
        round_inst_sbox_inst0_com_x_inst_n185), .Z(
        round_inst_sbox_inst0_com_x_inst_n186) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U42 ( .A1(round_inst_sin_z[0]), 
        .A2(round_inst_n70), .ZN(round_inst_sbox_inst0_com_x_inst_n185) );
  AND2_X1 round_inst_sbox_inst0_com_x_inst_U41 ( .A1(round_inst_sin_y[0]), 
        .A2(round_inst_sin_y[1]), .ZN(round_inst_sbox_inst0_com_x_inst_n222)
         );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U40 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n184), .A2(
        round_inst_sbox_inst0_com_x_inst_n229), .ZN(
        round_inst_sbox_inst0_com_x_inst_n205) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U39 ( .A1(round_inst_sin_y[0]), 
        .A2(round_inst_n70), .ZN(round_inst_sbox_inst0_com_x_inst_n229) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U38 ( .A(round_inst_sin_w[3]), .B(
        round_inst_sin_z[3]), .ZN(round_inst_sbox_inst0_com_x_inst_n184) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U37 ( .A(din[2]), .B(
        round_inst_sbox_inst0_com_x_inst_n248), .Z(
        round_inst_sbox_inst0_com_x_inst_n210) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U36 ( .A(
        round_inst_sbox_inst0_com_x_inst_n183), .B(
        round_inst_sbox_inst0_com_x_inst_n182), .ZN(
        round_inst_sbox_inst0_com_x_inst_n248) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U35 ( .A1(round_inst_sin_w[2]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n181), .ZN(
        round_inst_sbox_inst0_com_x_inst_n182) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U34 ( .A(
        round_inst_sbox_inst0_com_x_inst_n188), .B(
        round_inst_sbox_inst0_com_x_inst_n180), .Z(
        round_inst_sbox_inst0_com_x_inst_n181) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U33 ( .A1(round_inst_sin_y[1]), 
        .A2(round_inst_sin_w[3]), .ZN(round_inst_sbox_inst0_com_x_inst_n180)
         );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U32 ( .A(
        round_inst_sbox_inst0_com_x_inst_n179), .B(
        round_inst_sbox_inst0_com_x_inst_n178), .ZN(
        round_inst_sbox_inst0_com_x_inst_n183) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U31 ( .A(
        round_inst_sbox_inst0_com_x_inst_n177), .B(
        round_inst_sbox_inst0_com_x_inst_n176), .ZN(
        round_inst_sbox_inst0_com_x_inst_n178) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U30 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n286), .A2(round_inst_sin_z[1]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n176) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U29 ( .A(
        round_inst_sbox_inst0_com_x_inst_n175), .B(
        round_inst_sbox_inst0_com_x_inst_n255), .Z(
        round_inst_sbox_inst0_com_x_inst_n286) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U28 ( .A1(round_inst_n40), .A2(
        round_inst_sin_z[2]), .ZN(round_inst_sbox_inst0_com_x_inst_n255) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U27 ( .A1(round_inst_sin_z[3]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n295), .ZN(
        round_inst_sbox_inst0_com_x_inst_n175) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U26 ( .A(
        round_inst_sbox_inst0_com_x_inst_n174), .B(
        round_inst_sbox_inst0_com_x_inst_n173), .Z(
        round_inst_sbox_inst0_com_x_inst_n177) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U25 ( .A(
        round_inst_sbox_inst0_com_x_inst_n172), .B(
        round_inst_sbox_inst0_com_x_inst_n171), .ZN(
        round_inst_sbox_inst0_com_x_inst_n173) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U24 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n188), .A2(
        round_inst_sbox_inst0_com_x_inst_n295), .ZN(
        round_inst_sbox_inst0_com_x_inst_n171) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U23 ( .A1(round_inst_sin_z[1]), 
        .A2(round_inst_n40), .ZN(round_inst_sbox_inst0_com_x_inst_n188) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U22 ( .A(
        round_inst_sbox_inst0_com_x_inst_n170), .B(
        round_inst_sbox_inst0_com_x_inst_n169), .ZN(
        round_inst_sbox_inst0_com_x_inst_n172) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U21 ( .A(
        round_inst_sbox_inst0_com_x_inst_n168), .B(
        round_inst_sbox_inst0_com_x_inst_n167), .Z(
        round_inst_sbox_inst0_com_x_inst_n169) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U20 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n166), .A2(round_inst_sin_z[3]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n167) );
  INV_X1 round_inst_sbox_inst0_com_x_inst_U19 ( .A(
        round_inst_sbox_inst0_com_x_inst_n165), .ZN(
        round_inst_sbox_inst0_com_x_inst_n166) );
  NAND3_X1 round_inst_sbox_inst0_com_x_inst_U18 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n164), .A2(round_inst_sin_w[3]), .A3(
        round_inst_sbox_inst0_com_x_inst_n295), .ZN(
        round_inst_sbox_inst0_com_x_inst_n168) );
  XOR2_X1 round_inst_sbox_inst0_com_x_inst_U17 ( .A(round_inst_sin_z[1]), .B(
        round_inst_sin_y[1]), .Z(round_inst_sbox_inst0_com_x_inst_n164) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U16 ( .A(
        round_inst_sbox_inst0_com_x_inst_n163), .B(
        round_inst_sbox_inst0_com_x_inst_n162), .ZN(
        round_inst_sbox_inst0_com_x_inst_n170) );
  NAND3_X1 round_inst_sbox_inst0_com_x_inst_U15 ( .A1(round_inst_sin_z[3]), 
        .A2(round_inst_n70), .A3(round_inst_sbox_inst0_com_x_inst_n295), .ZN(
        round_inst_sbox_inst0_com_x_inst_n162) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U14 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n287), .A2(
        round_inst_sbox_inst0_com_x_inst_n165), .ZN(
        round_inst_sbox_inst0_com_x_inst_n163) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U13 ( .A1(round_inst_sin_y[1]), 
        .A2(round_inst_sin_z[2]), .ZN(round_inst_sbox_inst0_com_x_inst_n165)
         );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U12 ( .A(
        round_inst_sbox_inst0_com_x_inst_n161), .B(
        round_inst_sbox_inst0_com_x_inst_n160), .ZN(
        round_inst_sbox_inst0_com_x_inst_n174) );
  NAND3_X1 round_inst_sbox_inst0_com_x_inst_U11 ( .A1(round_inst_n40), .A2(
        round_inst_n70), .A3(round_inst_sin_z[2]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n160) );
  NOR2_X1 round_inst_sbox_inst0_com_x_inst_U10 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n225), .A2(
        round_inst_sbox_inst0_com_x_inst_n159), .ZN(
        round_inst_sbox_inst0_com_x_inst_n161) );
  OR2_X1 round_inst_sbox_inst0_com_x_inst_U9 ( .A1(
        round_inst_sbox_inst0_com_x_inst_n228), .A2(
        round_inst_sbox_inst0_com_x_inst_n275), .ZN(
        round_inst_sbox_inst0_com_x_inst_n159) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U8 ( .A(round_inst_n40), .B(
        round_inst_sin_z[3]), .ZN(round_inst_sbox_inst0_com_x_inst_n275) );
  INV_X1 round_inst_sbox_inst0_com_x_inst_U7 ( .A(round_inst_sin_y[1]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n228) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U6 ( .A(
        round_inst_sbox_inst0_com_x_inst_n295), .B(round_inst_sin_w[2]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n225) );
  INV_X1 round_inst_sbox_inst0_com_x_inst_U5 ( .A(
        round_inst_sbox_inst0_com_x_inst_n288), .ZN(
        round_inst_sbox_inst0_com_x_inst_n295) );
  INV_X1 round_inst_sbox_inst0_com_x_inst_U4 ( .A(round_inst_sin_y[2]), .ZN(
        round_inst_sbox_inst0_com_x_inst_n288) );
  NAND2_X1 round_inst_sbox_inst0_com_x_inst_U3 ( .A1(round_inst_sin_y[1]), 
        .A2(round_inst_sbox_inst0_com_x_inst_n214), .ZN(
        round_inst_sbox_inst0_com_x_inst_n179) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U2 ( .A(round_inst_sin_z[3]), .B(
        round_inst_sbox_inst0_com_x_inst_n287), .ZN(
        round_inst_sbox_inst0_com_x_inst_n214) );
  XNOR2_X1 round_inst_sbox_inst0_com_x_inst_U1 ( .A(round_inst_sin_w[3]), .B(
        round_inst_n40), .ZN(round_inst_sbox_inst0_com_x_inst_n287) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U144 ( .A(
        round_inst_sbox_inst0_com_y_inst_n155), .B(
        round_inst_sbox_inst0_com_y_inst_n154), .Z(round_inst_sout_y[0]) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U143 ( .A(
        round_inst_sbox_inst0_com_y_inst_n153), .B(
        round_inst_sbox_inst0_com_y_inst_n152), .ZN(
        round_inst_sbox_inst0_com_y_inst_n154) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U142 ( .A(
        round_inst_sbox_inst0_com_y_inst_n151), .B(round_inst_sin_z[3]), .Z(
        round_inst_sbox_inst0_com_y_inst_n152) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U141 ( .A(bin[0]), .B(
        round_inst_sbox_inst0_com_y_inst_n150), .Z(
        round_inst_sbox_inst0_com_y_inst_n153) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U140 ( .A(
        round_inst_sbox_inst0_com_y_inst_n149), .B(
        round_inst_sbox_inst0_com_y_inst_n148), .ZN(round_inst_srout2_y[18])
         );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U139 ( .A(
        round_inst_sbox_inst0_com_y_inst_n155), .B(
        round_inst_sbox_inst0_com_y_inst_n147), .ZN(
        round_inst_sbox_inst0_com_y_inst_n148) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U138 ( .A(
        round_inst_sbox_inst0_com_y_inst_n146), .B(
        round_inst_sbox_inst0_com_y_inst_n145), .ZN(
        round_inst_sbox_inst0_com_y_inst_n147) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U137 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n144), .A2(round_inst_sin_w[0]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n145) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U136 ( .A(
        round_inst_sbox_inst0_com_y_inst_n143), .B(bin[3]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n146) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U135 ( .A(
        round_inst_sbox_inst0_com_y_inst_n142), .B(
        round_inst_sbox_inst0_com_y_inst_n141), .ZN(
        round_inst_sbox_inst0_com_y_inst_n155) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U134 ( .A(
        round_inst_sbox_inst0_com_y_inst_n140), .B(
        round_inst_sbox_inst0_com_y_inst_n139), .ZN(
        round_inst_sbox_inst0_com_y_inst_n141) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U133 ( .A(
        round_inst_sbox_inst0_com_y_inst_n138), .B(
        round_inst_sbox_inst0_com_y_inst_n137), .Z(
        round_inst_sbox_inst0_com_y_inst_n140) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U132 ( .A(
        round_inst_sbox_inst0_com_y_inst_n136), .B(
        round_inst_sbox_inst0_com_y_inst_n135), .Z(
        round_inst_sbox_inst0_com_y_inst_n149) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U131 ( .A(
        round_inst_sbox_inst0_com_y_inst_n134), .B(
        round_inst_sbox_inst0_com_y_inst_n133), .ZN(
        round_inst_sbox_inst0_com_y_inst_n135) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U130 ( .A(
        round_inst_sbox_inst0_com_y_inst_n132), .B(
        round_inst_sbox_inst0_com_y_inst_n131), .Z(
        round_inst_sbox_inst0_com_y_inst_n133) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U129 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n130), .A2(
        round_inst_sbox_inst0_com_y_inst_n129), .ZN(
        round_inst_sbox_inst0_com_y_inst_n131) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U128 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n128), .A2(
        round_inst_sbox_inst0_com_y_inst_n127), .ZN(
        round_inst_sbox_inst0_com_y_inst_n132) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U127 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n126), .A2(round_inst_sin_x[0]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n134) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U126 ( .A(
        round_inst_sbox_inst0_com_y_inst_n139), .B(
        round_inst_sbox_inst0_com_y_inst_n137), .ZN(
        round_inst_sbox_inst0_com_y_inst_n126) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U125 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n151), .A2(
        round_inst_sbox_inst0_com_y_inst_n125), .ZN(
        round_inst_sbox_inst0_com_y_inst_n137) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U124 ( .A(
        round_inst_sbox_inst0_com_y_inst_n124), .B(
        round_inst_sbox_inst0_com_y_inst_n123), .ZN(
        round_inst_sbox_inst0_com_y_inst_n136) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U123 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n122), .A2(round_inst_sin_z[3]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n123) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U122 ( .A(
        round_inst_sbox_inst0_com_y_inst_n129), .B(
        round_inst_sbox_inst0_com_y_inst_n121), .Z(
        round_inst_sbox_inst0_com_y_inst_n122) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U121 ( .A1(round_inst_sin_w[2]), 
        .A2(round_inst_sin_x[0]), .ZN(round_inst_sbox_inst0_com_y_inst_n121)
         );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U120 ( .A(
        round_inst_sbox_inst0_com_y_inst_n120), .B(
        round_inst_sbox_inst0_com_y_inst_n119), .Z(
        round_inst_sbox_inst0_com_y_inst_n124) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U119 ( .A(
        round_inst_sbox_inst0_com_y_inst_n118), .B(
        round_inst_sbox_inst0_com_y_inst_n117), .ZN(
        round_inst_sbox_inst0_com_y_inst_n119) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U118 ( .A(
        round_inst_sbox_inst0_com_y_inst_n116), .B(
        round_inst_sbox_inst0_com_y_inst_n115), .Z(
        round_inst_sbox_inst0_com_y_inst_n117) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U117 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n114), .A2(
        round_inst_sbox_inst0_com_y_inst_n113), .ZN(
        round_inst_sbox_inst0_com_y_inst_n115) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U116 ( .A(
        round_inst_sbox_inst0_com_y_inst_n112), .B(
        round_inst_sbox_inst0_com_y_inst_n111), .ZN(
        round_inst_sbox_inst0_com_y_inst_n114) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U115 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n110), .A2(
        round_inst_sbox_inst0_com_y_inst_n109), .ZN(
        round_inst_sbox_inst0_com_y_inst_n112) );
  NAND3_X1 round_inst_sbox_inst0_com_y_inst_U114 ( .A1(round_inst_sin_z[0]), 
        .A2(round_inst_sbox_inst0_com_y_inst_n108), .A3(
        round_inst_sbox_inst0_com_y_inst_n107), .ZN(
        round_inst_sbox_inst0_com_y_inst_n116) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U113 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n106), .A2(
        round_inst_sbox_inst0_com_y_inst_n129), .ZN(
        round_inst_sbox_inst0_com_y_inst_n118) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U112 ( .A(
        round_inst_sbox_inst0_com_y_inst_n105), .B(
        round_inst_sbox_inst0_com_y_inst_n104), .ZN(round_inst_srout2_y[16])
         );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U111 ( .A(
        round_inst_sbox_inst0_com_y_inst_n103), .B(
        round_inst_sbox_inst0_com_y_inst_n102), .ZN(
        round_inst_sbox_inst0_com_y_inst_n104) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U110 ( .A(
        round_inst_sbox_inst0_com_y_inst_n142), .B(
        round_inst_sbox_inst0_com_y_inst_n101), .ZN(
        round_inst_sbox_inst0_com_y_inst_n102) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U109 ( .A(
        round_inst_sbox_inst0_com_y_inst_n100), .B(
        round_inst_sbox_inst0_com_y_inst_n99), .ZN(
        round_inst_sbox_inst0_com_y_inst_n142) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U108 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n98), .A2(round_inst_sin_z[1]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n99) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U107 ( .A(
        round_inst_sbox_inst0_com_y_inst_n97), .B(
        round_inst_sbox_inst0_com_y_inst_n127), .Z(
        round_inst_sbox_inst0_com_y_inst_n98) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U106 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n96), .A2(
        round_inst_sbox_inst0_com_y_inst_n108), .ZN(
        round_inst_sbox_inst0_com_y_inst_n97) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U105 ( .A(round_inst_sin_x[0]), .B(
        round_inst_sbox_inst0_com_y_inst_n95), .Z(
        round_inst_sbox_inst0_com_y_inst_n96) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U104 ( .A(
        round_inst_sbox_inst0_com_y_inst_n94), .B(
        round_inst_sbox_inst0_com_y_inst_n93), .ZN(
        round_inst_sbox_inst0_com_y_inst_n100) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U103 ( .A(
        round_inst_sbox_inst0_com_y_inst_n92), .B(
        round_inst_sbox_inst0_com_y_inst_n91), .Z(
        round_inst_sbox_inst0_com_y_inst_n93) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U102 ( .A(
        round_inst_sbox_inst0_com_y_inst_n90), .B(
        round_inst_sbox_inst0_com_y_inst_n89), .ZN(
        round_inst_sbox_inst0_com_y_inst_n91) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U101 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n88), .A2(round_inst_sin_x[2]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n89) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U100 ( .A(
        round_inst_sbox_inst0_com_y_inst_n87), .B(
        round_inst_sbox_inst0_com_y_inst_n86), .ZN(
        round_inst_sbox_inst0_com_y_inst_n90) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U99 ( .A(
        round_inst_sbox_inst0_com_y_inst_n85), .B(
        round_inst_sbox_inst0_com_y_inst_n84), .ZN(
        round_inst_sbox_inst0_com_y_inst_n86) );
  NAND3_X1 round_inst_sbox_inst0_com_y_inst_U98 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n83), .A2(round_inst_n70), .A3(
        round_inst_sbox_inst0_com_y_inst_n108), .ZN(
        round_inst_sbox_inst0_com_y_inst_n84) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U97 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n82), .A2(
        round_inst_sbox_inst0_com_y_inst_n81), .ZN(
        round_inst_sbox_inst0_com_y_inst_n85) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U96 ( .A(
        round_inst_sbox_inst0_com_y_inst_n80), .ZN(
        round_inst_sbox_inst0_com_y_inst_n81) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U95 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n79), .A2(
        round_inst_sbox_inst0_com_y_inst_n108), .ZN(
        round_inst_sbox_inst0_com_y_inst_n87) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U94 ( .A(
        round_inst_sbox_inst0_com_y_inst_n78), .B(
        round_inst_sbox_inst0_com_y_inst_n80), .Z(
        round_inst_sbox_inst0_com_y_inst_n79) );
  MUX2_X1 round_inst_sbox_inst0_com_y_inst_U93 ( .A(round_inst_sin_x[1]), .B(
        round_inst_n70), .S(round_inst_sbox_inst0_com_y_inst_n95), .Z(
        round_inst_sbox_inst0_com_y_inst_n78) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U92 ( .A1(round_inst_sin_w[2]), 
        .A2(round_inst_sbox_inst0_com_y_inst_n77), .ZN(
        round_inst_sbox_inst0_com_y_inst_n92) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U91 ( .A(
        round_inst_sbox_inst0_com_y_inst_n76), .B(
        round_inst_sbox_inst0_com_y_inst_n75), .ZN(
        round_inst_sbox_inst0_com_y_inst_n77) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U90 ( .A1(round_inst_sin_w[0]), 
        .A2(round_inst_sbox_inst0_com_y_inst_n143), .ZN(
        round_inst_sbox_inst0_com_y_inst_n76) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U89 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n82), .A2(
        round_inst_sbox_inst0_com_y_inst_n74), .ZN(
        round_inst_sbox_inst0_com_y_inst_n94) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U88 ( .A(
        round_inst_sbox_inst0_com_y_inst_n73), .B(
        round_inst_sbox_inst0_com_y_inst_n72), .ZN(
        round_inst_sbox_inst0_com_y_inst_n74) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U87 ( .A(
        round_inst_sbox_inst0_com_y_inst_n129), .B(bin[1]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n103) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U86 ( .A1(round_inst_sin_w[0]), 
        .A2(round_inst_sbox_inst0_com_y_inst_n108), .ZN(
        round_inst_sbox_inst0_com_y_inst_n129) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U85 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n71), .A2(round_inst_sin_z[0]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n105) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U84 ( .A(
        round_inst_sbox_inst0_com_y_inst_n82), .B(
        round_inst_sbox_inst0_com_y_inst_n151), .Z(
        round_inst_sbox_inst0_com_y_inst_n71) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U83 ( .A(
        round_inst_sbox_inst0_com_y_inst_n127), .B(round_inst_sin_w[2]), .Z(
        round_inst_sbox_inst0_com_y_inst_n82) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U82 ( .A(
        round_inst_sbox_inst0_com_y_inst_n101), .B(
        round_inst_sbox_inst0_com_y_inst_n70), .Z(round_inst_srout2_y[19]) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U81 ( .A(
        round_inst_sbox_inst0_com_y_inst_n69), .B(
        round_inst_sbox_inst0_com_y_inst_n68), .ZN(
        round_inst_sbox_inst0_com_y_inst_n70) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U80 ( .A(
        round_inst_sbox_inst0_com_y_inst_n113), .B(
        round_inst_sbox_inst0_com_y_inst_n120), .Z(
        round_inst_sbox_inst0_com_y_inst_n68) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U79 ( .A(
        round_inst_sbox_inst0_com_y_inst_n67), .B(
        round_inst_sbox_inst0_com_y_inst_n66), .ZN(
        round_inst_sbox_inst0_com_y_inst_n120) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U78 ( .A(
        round_inst_sbox_inst0_com_y_inst_n65), .B(
        round_inst_sbox_inst0_com_y_inst_n64), .ZN(
        round_inst_sbox_inst0_com_y_inst_n66) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U77 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n106), .A2(
        round_inst_sbox_inst0_com_y_inst_n75), .ZN(
        round_inst_sbox_inst0_com_y_inst_n64) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U76 ( .A(
        round_inst_sbox_inst0_com_y_inst_n63), .B(
        round_inst_sbox_inst0_com_y_inst_n62), .ZN(
        round_inst_sbox_inst0_com_y_inst_n65) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U75 ( .A(
        round_inst_sbox_inst0_com_y_inst_n61), .B(
        round_inst_sbox_inst0_com_y_inst_n60), .ZN(
        round_inst_sbox_inst0_com_y_inst_n62) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U74 ( .A(
        round_inst_sbox_inst0_com_y_inst_n59), .B(
        round_inst_sbox_inst0_com_y_inst_n58), .ZN(
        round_inst_sbox_inst0_com_y_inst_n60) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U73 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n57), .A2(
        round_inst_sbox_inst0_com_y_inst_n72), .ZN(
        round_inst_sbox_inst0_com_y_inst_n58) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U72 ( .A(
        round_inst_sbox_inst0_com_y_inst_n56), .B(round_inst_sin_x[3]), .Z(
        round_inst_sbox_inst0_com_y_inst_n57) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U71 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n56), .A2(
        round_inst_sbox_inst0_com_y_inst_n55), .ZN(
        round_inst_sbox_inst0_com_y_inst_n59) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U70 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n95), .A2(
        round_inst_sbox_inst0_com_y_inst_n54), .ZN(
        round_inst_sbox_inst0_com_y_inst_n55) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U69 ( .A(
        round_inst_sbox_inst0_com_y_inst_n53), .B(
        round_inst_sbox_inst0_com_y_inst_n52), .ZN(
        round_inst_sbox_inst0_com_y_inst_n61) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U68 ( .A(
        round_inst_sbox_inst0_com_y_inst_n51), .B(
        round_inst_sbox_inst0_com_y_inst_n50), .Z(
        round_inst_sbox_inst0_com_y_inst_n52) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U67 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n72), .A2(
        round_inst_sbox_inst0_com_y_inst_n106), .ZN(
        round_inst_sbox_inst0_com_y_inst_n50) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U66 ( .A1(round_inst_sin_z[1]), 
        .A2(round_inst_sin_x[0]), .ZN(round_inst_sbox_inst0_com_y_inst_n72) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U65 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n130), .A2(
        round_inst_sbox_inst0_com_y_inst_n73), .ZN(
        round_inst_sbox_inst0_com_y_inst_n51) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U64 ( .A(round_inst_sin_x[3]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n130) );
  NAND3_X1 round_inst_sbox_inst0_com_y_inst_U63 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n83), .A2(round_inst_n70), .A3(
        round_inst_sin_z[3]), .ZN(round_inst_sbox_inst0_com_y_inst_n53) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U62 ( .A(
        round_inst_sbox_inst0_com_y_inst_n113), .B(round_inst_sin_x[0]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n83) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U61 ( .A(
        round_inst_sbox_inst0_com_y_inst_n49), .B(
        round_inst_sbox_inst0_com_y_inst_n48), .Z(
        round_inst_sbox_inst0_com_y_inst_n63) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U60 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n88), .A2(
        round_inst_sbox_inst0_com_y_inst_n47), .ZN(
        round_inst_sbox_inst0_com_y_inst_n48) );
  NAND3_X1 round_inst_sbox_inst0_com_y_inst_U59 ( .A1(round_inst_sin_x[1]), 
        .A2(round_inst_sin_w[0]), .A3(round_inst_sin_z[3]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n49) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U58 ( .A(
        round_inst_sbox_inst0_com_y_inst_n46), .B(
        round_inst_sbox_inst0_com_y_inst_n45), .Z(
        round_inst_sbox_inst0_com_y_inst_n67) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U57 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n107), .A2(
        round_inst_sbox_inst0_com_y_inst_n80), .ZN(
        round_inst_sbox_inst0_com_y_inst_n45) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U56 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n113), .A2(
        round_inst_sbox_inst0_com_y_inst_n143), .ZN(
        round_inst_sbox_inst0_com_y_inst_n80) );
  NOR3_X1 round_inst_sbox_inst0_com_y_inst_U55 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n113), .A2(
        round_inst_sbox_inst0_com_y_inst_n106), .A3(
        round_inst_sbox_inst0_com_y_inst_n54), .ZN(
        round_inst_sbox_inst0_com_y_inst_n46) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U54 ( .A(round_inst_sin_z[0]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n113) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U53 ( .A(bin[2]), .B(
        round_inst_sbox_inst0_com_y_inst_n150), .Z(
        round_inst_sbox_inst0_com_y_inst_n69) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U52 ( .A(
        round_inst_sbox_inst0_com_y_inst_n44), .B(
        round_inst_sbox_inst0_com_y_inst_n43), .ZN(
        round_inst_sbox_inst0_com_y_inst_n150) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U51 ( .A(
        round_inst_sbox_inst0_com_y_inst_n42), .B(
        round_inst_sbox_inst0_com_y_inst_n41), .ZN(
        round_inst_sbox_inst0_com_y_inst_n43) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U50 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n40), .A2(round_inst_sin_z[0]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n41) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U49 ( .A(
        round_inst_sbox_inst0_com_y_inst_n39), .B(
        round_inst_sbox_inst0_com_y_inst_n125), .ZN(
        round_inst_sbox_inst0_com_y_inst_n40) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U48 ( .A(
        round_inst_sbox_inst0_com_y_inst_n47), .ZN(
        round_inst_sbox_inst0_com_y_inst_n125) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U47 ( .A(round_inst_sin_w[3]), .B(
        round_inst_sin_x[3]), .Z(round_inst_sbox_inst0_com_y_inst_n47) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U46 ( .A(round_inst_sin_z[1]), .B(
        round_inst_sin_z[3]), .Z(round_inst_sbox_inst0_com_y_inst_n39) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U45 ( .A(
        round_inst_sbox_inst0_com_y_inst_n73), .B(
        round_inst_sbox_inst0_com_y_inst_n128), .ZN(
        round_inst_sbox_inst0_com_y_inst_n42) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U44 ( .A1(round_inst_sin_w[0]), 
        .A2(round_inst_sin_z[3]), .ZN(round_inst_sbox_inst0_com_y_inst_n128)
         );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U43 ( .A1(round_inst_sin_z[0]), 
        .A2(round_inst_n70), .ZN(round_inst_sbox_inst0_com_y_inst_n73) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U42 ( .A(
        round_inst_sbox_inst0_com_y_inst_n75), .B(
        round_inst_sbox_inst0_com_y_inst_n88), .ZN(
        round_inst_sbox_inst0_com_y_inst_n44) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U41 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n143), .A2(
        round_inst_sbox_inst0_com_y_inst_n95), .ZN(
        round_inst_sbox_inst0_com_y_inst_n88) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U40 ( .A(round_inst_sin_w[0]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n95) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U39 ( .A1(round_inst_sin_z[0]), 
        .A2(round_inst_sin_x[1]), .ZN(round_inst_sbox_inst0_com_y_inst_n75) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U38 ( .A(
        round_inst_sbox_inst0_com_y_inst_n38), .B(
        round_inst_sbox_inst0_com_y_inst_n37), .ZN(
        round_inst_sbox_inst0_com_y_inst_n101) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U37 ( .A(
        round_inst_sbox_inst0_com_y_inst_n36), .B(
        round_inst_sbox_inst0_com_y_inst_n35), .ZN(
        round_inst_sbox_inst0_com_y_inst_n37) );
  NAND3_X1 round_inst_sbox_inst0_com_y_inst_U36 ( .A1(round_inst_n70), .A2(
        round_inst_sin_z[3]), .A3(round_inst_sbox_inst0_com_y_inst_n127), .ZN(
        round_inst_sbox_inst0_com_y_inst_n35) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U35 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n34), .A2(round_inst_sin_x[3]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n36) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U34 ( .A(
        round_inst_sbox_inst0_com_y_inst_n33), .B(
        round_inst_sbox_inst0_com_y_inst_n32), .ZN(
        round_inst_sbox_inst0_com_y_inst_n34) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U33 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n31), .A2(
        round_inst_sbox_inst0_com_y_inst_n151), .ZN(
        round_inst_sbox_inst0_com_y_inst_n32) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U32 ( .A(
        round_inst_sbox_inst0_com_y_inst_n143), .B(round_inst_sin_x[1]), .Z(
        round_inst_sbox_inst0_com_y_inst_n31) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U31 ( .A1(round_inst_sin_w[2]), 
        .A2(round_inst_sin_z[1]), .ZN(round_inst_sbox_inst0_com_y_inst_n33) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U30 ( .A(
        round_inst_sbox_inst0_com_y_inst_n30), .B(
        round_inst_sbox_inst0_com_y_inst_n29), .ZN(
        round_inst_sbox_inst0_com_y_inst_n38) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U29 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n54), .A2(
        round_inst_sbox_inst0_com_y_inst_n138), .ZN(
        round_inst_sbox_inst0_com_y_inst_n29) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U28 ( .A(
        round_inst_sbox_inst0_com_y_inst_n144), .ZN(
        round_inst_sbox_inst0_com_y_inst_n138) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U27 ( .A(round_inst_n70), .B(
        round_inst_sbox_inst0_com_y_inst_n143), .Z(
        round_inst_sbox_inst0_com_y_inst_n54) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U26 ( .A(round_inst_sin_z[1]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n143) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U25 ( .A(
        round_inst_sbox_inst0_com_y_inst_n28), .B(
        round_inst_sbox_inst0_com_y_inst_n27), .ZN(
        round_inst_sbox_inst0_com_y_inst_n30) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U24 ( .A(
        round_inst_sbox_inst0_com_y_inst_n26), .B(
        round_inst_sbox_inst0_com_y_inst_n25), .ZN(
        round_inst_sbox_inst0_com_y_inst_n27) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U23 ( .A(
        round_inst_sbox_inst0_com_y_inst_n24), .B(
        round_inst_sbox_inst0_com_y_inst_n23), .Z(
        round_inst_sbox_inst0_com_y_inst_n25) );
  NAND3_X1 round_inst_sbox_inst0_com_y_inst_U22 ( .A1(round_inst_sin_z[1]), 
        .A2(round_inst_sin_w[3]), .A3(round_inst_sin_w[2]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n23) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U21 ( .A1(round_inst_sin_x[1]), 
        .A2(round_inst_sbox_inst0_com_y_inst_n144), .ZN(
        round_inst_sbox_inst0_com_y_inst_n24) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U20 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n110), .A2(
        round_inst_sbox_inst0_com_y_inst_n56), .ZN(
        round_inst_sbox_inst0_com_y_inst_n144) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U19 ( .A(round_inst_sin_w[2]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n110) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U18 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n22), .A2(round_inst_sin_z[1]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n26) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U17 ( .A(
        round_inst_sbox_inst0_com_y_inst_n21), .B(
        round_inst_sbox_inst0_com_y_inst_n111), .ZN(
        round_inst_sbox_inst0_com_y_inst_n22) );
  NOR2_X1 round_inst_sbox_inst0_com_y_inst_U16 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n20), .A2(
        round_inst_sbox_inst0_com_y_inst_n106), .ZN(
        round_inst_sbox_inst0_com_y_inst_n111) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U15 ( .A(
        round_inst_sbox_inst0_com_y_inst_n127), .B(
        round_inst_sbox_inst0_com_y_inst_n108), .Z(
        round_inst_sbox_inst0_com_y_inst_n20) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U14 ( .A(round_inst_sin_x[2]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n127) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U13 ( .A(
        round_inst_sbox_inst0_com_y_inst_n139), .B(
        round_inst_sbox_inst0_com_y_inst_n109), .ZN(
        round_inst_sbox_inst0_com_y_inst_n21) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U12 ( .A(
        round_inst_sbox_inst0_com_y_inst_n106), .B(
        round_inst_sbox_inst0_com_y_inst_n107), .Z(
        round_inst_sbox_inst0_com_y_inst_n109) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U11 ( .A(
        round_inst_sbox_inst0_com_y_inst_n56), .B(round_inst_sin_x[3]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n107) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U10 ( .A(round_inst_sin_w[3]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n106) );
  NAND2_X1 round_inst_sbox_inst0_com_y_inst_U9 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n108), .A2(round_inst_sin_z[3]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n139) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U8 ( .A(
        round_inst_sbox_inst0_com_y_inst_n19), .B(
        round_inst_sbox_inst0_com_y_inst_n18), .Z(
        round_inst_sbox_inst0_com_y_inst_n28) );
  NAND3_X1 round_inst_sbox_inst0_com_y_inst_U7 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n108), .A2(round_inst_sin_x[3]), .A3(
        round_inst_n70), .ZN(round_inst_sbox_inst0_com_y_inst_n18) );
  NAND3_X1 round_inst_sbox_inst0_com_y_inst_U6 ( .A1(
        round_inst_sbox_inst0_com_y_inst_n17), .A2(
        round_inst_sbox_inst0_com_y_inst_n108), .A3(
        round_inst_sbox_inst0_com_y_inst_n16), .ZN(
        round_inst_sbox_inst0_com_y_inst_n19) );
  XNOR2_X1 round_inst_sbox_inst0_com_y_inst_U5 ( .A(
        round_inst_sbox_inst0_com_y_inst_n56), .B(round_inst_sin_w[3]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n16) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U4 ( .A(round_inst_sin_z[3]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n56) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U3 ( .A(
        round_inst_sbox_inst0_com_y_inst_n151), .ZN(
        round_inst_sbox_inst0_com_y_inst_n108) );
  INV_X1 round_inst_sbox_inst0_com_y_inst_U2 ( .A(round_inst_sin_z[2]), .ZN(
        round_inst_sbox_inst0_com_y_inst_n151) );
  XOR2_X1 round_inst_sbox_inst0_com_y_inst_U1 ( .A(round_inst_n70), .B(
        round_inst_sin_x[1]), .Z(round_inst_sbox_inst0_com_y_inst_n17) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U135 ( .A(
        round_inst_sbox_inst0_com_z_inst_n274), .B(
        round_inst_sbox_inst0_com_z_inst_n273), .ZN(round_inst_sout_z[0]) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U134 ( .A(round_inst_sin_w[3]), 
        .B(round_inst_sbox_inst0_com_z_inst_n272), .ZN(
        round_inst_sbox_inst0_com_z_inst_n273) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U133 ( .A(
        round_inst_sbox_inst0_com_z_inst_n271), .B(
        round_inst_sbox_inst0_com_z_inst_n270), .ZN(
        round_inst_sbox_inst0_com_z_inst_n274) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U132 ( .A(
        round_inst_sbox_inst0_com_z_inst_n269), .B(
        round_inst_sbox_inst0_com_z_inst_n268), .ZN(
        round_inst_sbox_inst0_com_z_inst_n271) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U131 ( .A(cin[0]), .B(bin[0]), .Z(
        round_inst_sbox_inst0_com_z_inst_n268) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U130 ( .A(
        round_inst_sbox_inst0_com_z_inst_n267), .B(
        round_inst_sbox_inst0_com_z_inst_n269), .ZN(round_inst_srout2_z[18])
         );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U129 ( .A(
        round_inst_sbox_inst0_com_z_inst_n266), .B(
        round_inst_sbox_inst0_com_z_inst_n265), .ZN(
        round_inst_sbox_inst0_com_z_inst_n269) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U128 ( .A(
        round_inst_sbox_inst0_com_z_inst_n264), .B(
        round_inst_sbox_inst0_com_z_inst_n263), .Z(
        round_inst_sbox_inst0_com_z_inst_n265) );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U127 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n262), .A2(
        round_inst_sbox_inst0_com_z_inst_n270), .ZN(
        round_inst_sbox_inst0_com_z_inst_n266) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U126 ( .A(
        round_inst_sbox_inst0_com_z_inst_n261), .B(
        round_inst_sbox_inst0_com_z_inst_n260), .ZN(
        round_inst_sbox_inst0_com_z_inst_n267) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U125 ( .A(
        round_inst_sbox_inst0_com_z_inst_n259), .B(cin[3]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n260) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U124 ( .A(
        round_inst_sbox_inst0_com_z_inst_n258), .B(
        round_inst_sbox_inst0_com_z_inst_n257), .Z(
        round_inst_sbox_inst0_com_z_inst_n261) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U123 ( .A(
        round_inst_sbox_inst0_com_z_inst_n256), .B(
        round_inst_sbox_inst0_com_z_inst_n255), .ZN(
        round_inst_sbox_inst0_com_z_inst_n257) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U122 ( .A(
        round_inst_sbox_inst0_com_z_inst_n254), .B(
        round_inst_sbox_inst0_com_z_inst_n253), .ZN(
        round_inst_sbox_inst0_com_z_inst_n255) );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U121 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n252), .A2(
        round_inst_sbox_inst0_com_z_inst_n251), .ZN(
        round_inst_sbox_inst0_com_z_inst_n253) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U120 ( .A(round_inst_n70), .B(
        bin[3]), .ZN(round_inst_sbox_inst0_com_z_inst_n254) );
  NAND3_X1 round_inst_sbox_inst0_com_z_inst_U119 ( .A1(round_inst_sin_w[0]), 
        .A2(round_inst_sin_x[2]), .A3(round_inst_sin_x[3]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n256) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U118 ( .A(
        round_inst_sbox_inst0_com_z_inst_n250), .B(
        round_inst_sbox_inst0_com_z_inst_n249), .ZN(
        round_inst_sbox_inst0_com_z_inst_n258) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U117 ( .A(
        round_inst_sbox_inst0_com_z_inst_n248), .B(
        round_inst_sbox_inst0_com_z_inst_n247), .Z(
        round_inst_sbox_inst0_com_z_inst_n249) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U116 ( .A(
        round_inst_sbox_inst0_com_z_inst_n246), .B(
        round_inst_sbox_inst0_com_z_inst_n245), .ZN(
        round_inst_sbox_inst0_com_z_inst_n247) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U115 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n264), .A2(round_inst_sin_y[0]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n245) );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U114 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n262), .A2(
        round_inst_sbox_inst0_com_z_inst_n244), .ZN(
        round_inst_sbox_inst0_com_z_inst_n246) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U113 ( .A1(round_inst_sin_w[0]), 
        .A2(round_inst_sin_x[2]), .ZN(round_inst_sbox_inst0_com_z_inst_n244)
         );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U112 ( .A(round_inst_sin_w[3]), 
        .B(round_inst_n40), .ZN(round_inst_sbox_inst0_com_z_inst_n262) );
  NAND3_X1 round_inst_sbox_inst0_com_z_inst_U111 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n243), .A2(round_inst_sin_w[3]), .A3(
        round_inst_sin_x[0]), .ZN(round_inst_sbox_inst0_com_z_inst_n248) );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U110 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n242), .A2(
        round_inst_sbox_inst0_com_z_inst_n241), .ZN(
        round_inst_sbox_inst0_com_z_inst_n250) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U109 ( .A(
        round_inst_sbox_inst0_com_z_inst_n240), .B(
        round_inst_sbox_inst0_com_z_inst_n239), .ZN(round_inst_srout2_z[16])
         );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U108 ( .A(
        round_inst_sbox_inst0_com_z_inst_n241), .B(cin[1]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n239) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U107 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n238), .A2(round_inst_sin_w[2]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n241) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U106 ( .A(bin[1]), .B(
        round_inst_sbox_inst0_com_z_inst_n237), .ZN(
        round_inst_sbox_inst0_com_z_inst_n240) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U105 ( .A(
        round_inst_sbox_inst0_com_z_inst_n236), .B(
        round_inst_sbox_inst0_com_z_inst_n235), .ZN(
        round_inst_sbox_inst0_com_z_inst_n237) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U104 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n243), .A2(round_inst_sin_w[0]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n235) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U103 ( .A(
        round_inst_sbox_inst0_com_z_inst_n234), .B(
        round_inst_sbox_inst0_com_z_inst_n263), .Z(
        round_inst_sbox_inst0_com_z_inst_n236) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U102 ( .A(
        round_inst_sbox_inst0_com_z_inst_n233), .B(
        round_inst_sbox_inst0_com_z_inst_n232), .ZN(
        round_inst_sbox_inst0_com_z_inst_n263) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U101 ( .A(
        round_inst_sbox_inst0_com_z_inst_n231), .B(
        round_inst_sbox_inst0_com_z_inst_n230), .Z(
        round_inst_sbox_inst0_com_z_inst_n232) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U100 ( .A1(round_inst_sin_x[2]), 
        .A2(round_inst_sbox_inst0_com_z_inst_n229), .ZN(
        round_inst_sbox_inst0_com_z_inst_n230) );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U99 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n228), .A2(
        round_inst_sbox_inst0_com_z_inst_n270), .ZN(
        round_inst_sbox_inst0_com_z_inst_n231) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U98 ( .A(
        round_inst_sbox_inst0_com_z_inst_n227), .B(
        round_inst_sbox_inst0_com_z_inst_n226), .ZN(
        round_inst_sbox_inst0_com_z_inst_n233) );
  NAND3_X1 round_inst_sbox_inst0_com_z_inst_U97 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n225), .A2(round_inst_sin_x[0]), .A3(
        round_inst_sin_w[2]), .ZN(round_inst_sbox_inst0_com_z_inst_n226) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U96 ( .A(round_inst_sin_y[1]), .B(
        round_inst_sin_x[1]), .Z(round_inst_sbox_inst0_com_z_inst_n225) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U95 ( .A(
        round_inst_sbox_inst0_com_z_inst_n224), .B(
        round_inst_sbox_inst0_com_z_inst_n223), .ZN(
        round_inst_sbox_inst0_com_z_inst_n227) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U94 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n243), .A2(
        round_inst_sbox_inst0_com_z_inst_n222), .ZN(
        round_inst_sbox_inst0_com_z_inst_n223) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U93 ( .A(round_inst_sin_x[2]), .B(
        round_inst_sbox_inst0_com_z_inst_n252), .ZN(
        round_inst_sbox_inst0_com_z_inst_n243) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U92 ( .A(
        round_inst_sbox_inst0_com_z_inst_n221), .B(
        round_inst_sbox_inst0_com_z_inst_n220), .Z(
        round_inst_sbox_inst0_com_z_inst_n224) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U91 ( .A(
        round_inst_sbox_inst0_com_z_inst_n219), .B(
        round_inst_sbox_inst0_com_z_inst_n218), .ZN(
        round_inst_sbox_inst0_com_z_inst_n220) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U90 ( .A1(round_inst_sin_w[2]), 
        .A2(round_inst_sbox_inst0_com_z_inst_n217), .ZN(
        round_inst_sbox_inst0_com_z_inst_n218) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U89 ( .A(
        round_inst_sbox_inst0_com_z_inst_n216), .B(
        round_inst_sbox_inst0_com_z_inst_n215), .Z(
        round_inst_sbox_inst0_com_z_inst_n219) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U88 ( .A(
        round_inst_sbox_inst0_com_z_inst_n214), .B(
        round_inst_sbox_inst0_com_z_inst_n213), .ZN(
        round_inst_sbox_inst0_com_z_inst_n215) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U87 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n212), .A2(round_inst_sin_w[2]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n213) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U86 ( .A(
        round_inst_sbox_inst0_com_z_inst_n211), .B(
        round_inst_sbox_inst0_com_z_inst_n210), .ZN(
        round_inst_sbox_inst0_com_z_inst_n212) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U85 ( .A(
        round_inst_sbox_inst0_com_z_inst_n209), .B(
        round_inst_sbox_inst0_com_z_inst_n208), .Z(
        round_inst_sbox_inst0_com_z_inst_n211) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U84 ( .A1(round_inst_sin_x[1]), 
        .A2(round_inst_sin_y[0]), .ZN(round_inst_sbox_inst0_com_z_inst_n208)
         );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U83 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n207), .A2(round_inst_sin_y[0]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n214) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U82 ( .A(
        round_inst_sbox_inst0_com_z_inst_n206), .B(
        round_inst_sbox_inst0_com_z_inst_n205), .ZN(
        round_inst_sbox_inst0_com_z_inst_n216) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U81 ( .A1(round_inst_n70), .A2(
        round_inst_sin_y[2]), .ZN(round_inst_sbox_inst0_com_z_inst_n205) );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U80 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n204), .A2(
        round_inst_sbox_inst0_com_z_inst_n210), .ZN(
        round_inst_sbox_inst0_com_z_inst_n206) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U79 ( .A(round_inst_sin_x[2]), .B(
        round_inst_sbox_inst0_com_z_inst_n252), .Z(
        round_inst_sbox_inst0_com_z_inst_n204) );
  INV_X1 round_inst_sbox_inst0_com_z_inst_U78 ( .A(round_inst_sin_y[2]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n252) );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U77 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n203), .A2(
        round_inst_sbox_inst0_com_z_inst_n202), .ZN(
        round_inst_sbox_inst0_com_z_inst_n221) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U76 ( .A(
        round_inst_sbox_inst0_com_z_inst_n270), .B(round_inst_sin_y[2]), .Z(
        round_inst_sbox_inst0_com_z_inst_n203) );
  INV_X1 round_inst_sbox_inst0_com_z_inst_U75 ( .A(round_inst_sin_w[2]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n270) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U74 ( .A(
        round_inst_sbox_inst0_com_z_inst_n201), .B(
        round_inst_sbox_inst0_com_z_inst_n200), .ZN(round_inst_srout2_z[19])
         );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U73 ( .A(
        round_inst_sbox_inst0_com_z_inst_n199), .B(
        round_inst_sbox_inst0_com_z_inst_n198), .ZN(
        round_inst_sbox_inst0_com_z_inst_n200) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U72 ( .A(round_inst_sin_w[0]), .B(
        round_inst_sbox_inst0_com_z_inst_n234), .ZN(
        round_inst_sbox_inst0_com_z_inst_n198) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U71 ( .A(
        round_inst_sbox_inst0_com_z_inst_n197), .B(
        round_inst_sbox_inst0_com_z_inst_n196), .ZN(
        round_inst_sbox_inst0_com_z_inst_n234) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U70 ( .A(
        round_inst_sbox_inst0_com_z_inst_n195), .B(
        round_inst_sbox_inst0_com_z_inst_n194), .ZN(
        round_inst_sbox_inst0_com_z_inst_n196) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U69 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n193), .A2(round_inst_n40), .ZN(
        round_inst_sbox_inst0_com_z_inst_n194) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U68 ( .A(
        round_inst_sbox_inst0_com_z_inst_n192), .B(
        round_inst_sbox_inst0_com_z_inst_n191), .ZN(
        round_inst_sbox_inst0_com_z_inst_n193) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U67 ( .A1(round_inst_sin_x[3]), 
        .A2(round_inst_sbox_inst0_com_z_inst_n192), .ZN(
        round_inst_sbox_inst0_com_z_inst_n195) );
  INV_X1 round_inst_sbox_inst0_com_z_inst_U66 ( .A(
        round_inst_sbox_inst0_com_z_inst_n207), .ZN(
        round_inst_sbox_inst0_com_z_inst_n192) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U65 ( .A1(round_inst_n70), .A2(
        round_inst_sin_x[2]), .ZN(round_inst_sbox_inst0_com_z_inst_n207) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U64 ( .A(
        round_inst_sbox_inst0_com_z_inst_n190), .B(
        round_inst_sbox_inst0_com_z_inst_n189), .ZN(
        round_inst_sbox_inst0_com_z_inst_n197) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U63 ( .A1(round_inst_sin_x[1]), 
        .A2(round_inst_sin_w[3]), .ZN(round_inst_sbox_inst0_com_z_inst_n189)
         );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U62 ( .A(
        round_inst_sbox_inst0_com_z_inst_n188), .B(
        round_inst_sbox_inst0_com_z_inst_n187), .ZN(
        round_inst_sbox_inst0_com_z_inst_n190) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U61 ( .A1(round_inst_sin_w[3]), 
        .A2(round_inst_sbox_inst0_com_z_inst_n186), .ZN(
        round_inst_sbox_inst0_com_z_inst_n187) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U60 ( .A(
        round_inst_sbox_inst0_com_z_inst_n185), .B(
        round_inst_sbox_inst0_com_z_inst_n184), .Z(
        round_inst_sbox_inst0_com_z_inst_n186) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U59 ( .A1(round_inst_sin_x[1]), 
        .A2(round_inst_sin_y[2]), .ZN(round_inst_sbox_inst0_com_z_inst_n184)
         );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U58 ( .A(
        round_inst_sbox_inst0_com_z_inst_n183), .B(
        round_inst_sbox_inst0_com_z_inst_n182), .ZN(
        round_inst_sbox_inst0_com_z_inst_n188) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U57 ( .A(
        round_inst_sbox_inst0_com_z_inst_n181), .B(
        round_inst_sbox_inst0_com_z_inst_n180), .ZN(
        round_inst_sbox_inst0_com_z_inst_n182) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U56 ( .A(
        round_inst_sbox_inst0_com_z_inst_n179), .B(
        round_inst_sbox_inst0_com_z_inst_n178), .Z(
        round_inst_sbox_inst0_com_z_inst_n180) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U55 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n264), .A2(round_inst_sin_y[1]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n178) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U54 ( .A(
        round_inst_sbox_inst0_com_z_inst_n177), .B(
        round_inst_sbox_inst0_com_z_inst_n176), .Z(
        round_inst_sbox_inst0_com_z_inst_n264) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U53 ( .A1(round_inst_sin_x[3]), 
        .A2(round_inst_sin_w[2]), .ZN(round_inst_sbox_inst0_com_z_inst_n176)
         );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U52 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n175), .A2(
        round_inst_sbox_inst0_com_z_inst_n185), .ZN(
        round_inst_sbox_inst0_com_z_inst_n179) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U51 ( .A1(round_inst_n70), .A2(
        round_inst_sin_w[2]), .ZN(round_inst_sbox_inst0_com_z_inst_n185) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U50 ( .A(
        round_inst_sbox_inst0_com_z_inst_n174), .B(
        round_inst_sbox_inst0_com_z_inst_n173), .ZN(
        round_inst_sbox_inst0_com_z_inst_n181) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U49 ( .A(
        round_inst_sbox_inst0_com_z_inst_n172), .B(
        round_inst_sbox_inst0_com_z_inst_n171), .Z(
        round_inst_sbox_inst0_com_z_inst_n173) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U48 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n170), .A2(round_inst_n70), .ZN(
        round_inst_sbox_inst0_com_z_inst_n171) );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U47 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n169), .A2(
        round_inst_sbox_inst0_com_z_inst_n191), .ZN(
        round_inst_sbox_inst0_com_z_inst_n172) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U46 ( .A1(round_inst_sin_x[1]), 
        .A2(round_inst_sin_w[2]), .ZN(round_inst_sbox_inst0_com_z_inst_n191)
         );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U45 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n177), .A2(
        round_inst_sbox_inst0_com_z_inst_n228), .ZN(
        round_inst_sbox_inst0_com_z_inst_n174) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U44 ( .A1(round_inst_sin_w[3]), 
        .A2(round_inst_sin_x[2]), .ZN(round_inst_sbox_inst0_com_z_inst_n177)
         );
  NAND3_X1 round_inst_sbox_inst0_com_z_inst_U43 ( .A1(round_inst_n70), .A2(
        round_inst_sbox_inst0_com_z_inst_n170), .A3(round_inst_sin_y[2]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n183) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U42 ( .A(bin[2]), .B(cin[2]), .Z(
        round_inst_sbox_inst0_com_z_inst_n199) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U41 ( .A(
        round_inst_sbox_inst0_com_z_inst_n272), .B(
        round_inst_sbox_inst0_com_z_inst_n259), .ZN(
        round_inst_sbox_inst0_com_z_inst_n201) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U40 ( .A(
        round_inst_sbox_inst0_com_z_inst_n168), .B(
        round_inst_sbox_inst0_com_z_inst_n167), .ZN(
        round_inst_sbox_inst0_com_z_inst_n259) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U39 ( .A(
        round_inst_sbox_inst0_com_z_inst_n166), .B(
        round_inst_sbox_inst0_com_z_inst_n165), .ZN(
        round_inst_sbox_inst0_com_z_inst_n167) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U38 ( .A(
        round_inst_sbox_inst0_com_z_inst_n164), .B(
        round_inst_sbox_inst0_com_z_inst_n163), .Z(
        round_inst_sbox_inst0_com_z_inst_n165) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U37 ( .A(
        round_inst_sbox_inst0_com_z_inst_n162), .B(
        round_inst_sbox_inst0_com_z_inst_n161), .ZN(
        round_inst_sbox_inst0_com_z_inst_n163) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U36 ( .A1(round_inst_n40), .A2(
        round_inst_sbox_inst0_com_z_inst_n217), .ZN(
        round_inst_sbox_inst0_com_z_inst_n161) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U35 ( .A(
        round_inst_sbox_inst0_com_z_inst_n160), .B(
        round_inst_sbox_inst0_com_z_inst_n159), .Z(
        round_inst_sbox_inst0_com_z_inst_n162) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U34 ( .A(
        round_inst_sbox_inst0_com_z_inst_n158), .B(
        round_inst_sbox_inst0_com_z_inst_n157), .ZN(
        round_inst_sbox_inst0_com_z_inst_n159) );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U33 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n156), .A2(
        round_inst_sbox_inst0_com_z_inst_n228), .ZN(
        round_inst_sbox_inst0_com_z_inst_n157) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U32 ( .A(round_inst_n70), .B(
        round_inst_sin_x[1]), .ZN(round_inst_sbox_inst0_com_z_inst_n228) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U31 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n155), .A2(round_inst_sin_x[3]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n158) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U30 ( .A(
        round_inst_sbox_inst0_com_z_inst_n209), .B(
        round_inst_sbox_inst0_com_z_inst_n154), .ZN(
        round_inst_sbox_inst0_com_z_inst_n155) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U29 ( .A(
        round_inst_sbox_inst0_com_z_inst_n217), .B(
        round_inst_sbox_inst0_com_z_inst_n153), .ZN(
        round_inst_sbox_inst0_com_z_inst_n154) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U28 ( .A1(round_inst_n70), .A2(
        round_inst_sin_y[0]), .ZN(round_inst_sbox_inst0_com_z_inst_n153) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U27 ( .A(
        round_inst_sbox_inst0_com_z_inst_n152), .B(
        round_inst_sbox_inst0_com_z_inst_n151), .ZN(
        round_inst_sbox_inst0_com_z_inst_n160) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U26 ( .A(
        round_inst_sbox_inst0_com_z_inst_n150), .B(
        round_inst_sbox_inst0_com_z_inst_n149), .Z(
        round_inst_sbox_inst0_com_z_inst_n151) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U25 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n229), .A2(round_inst_sin_x[3]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n149) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U24 ( .A1(round_inst_sin_y[1]), 
        .A2(round_inst_sbox_inst0_com_z_inst_n148), .ZN(
        round_inst_sbox_inst0_com_z_inst_n150) );
  NAND3_X1 round_inst_sbox_inst0_com_z_inst_U23 ( .A1(round_inst_sin_x[1]), 
        .A2(round_inst_sin_y[0]), .A3(round_inst_sin_w[3]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n152) );
  NAND3_X1 round_inst_sbox_inst0_com_z_inst_U22 ( .A1(round_inst_n70), .A2(
        round_inst_n40), .A3(round_inst_sbox_inst0_com_z_inst_n238), .ZN(
        round_inst_sbox_inst0_com_z_inst_n164) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U21 ( .A(round_inst_sin_x[0]), .B(
        round_inst_sin_w[0]), .Z(round_inst_sbox_inst0_com_z_inst_n238) );
  NOR2_X1 round_inst_sbox_inst0_com_z_inst_U20 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n175), .A2(
        round_inst_sbox_inst0_com_z_inst_n210), .ZN(
        round_inst_sbox_inst0_com_z_inst_n166) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U19 ( .A(round_inst_n40), .B(
        round_inst_sin_x[3]), .ZN(round_inst_sbox_inst0_com_z_inst_n175) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U18 ( .A1(
        round_inst_sbox_inst0_com_z_inst_n147), .A2(round_inst_sin_w[3]), .ZN(
        round_inst_sbox_inst0_com_z_inst_n168) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U17 ( .A(
        round_inst_sbox_inst0_com_z_inst_n217), .B(
        round_inst_sbox_inst0_com_z_inst_n146), .Z(
        round_inst_sbox_inst0_com_z_inst_n147) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U16 ( .A(
        round_inst_sbox_inst0_com_z_inst_n222), .B(
        round_inst_sbox_inst0_com_z_inst_n145), .ZN(
        round_inst_sbox_inst0_com_z_inst_n272) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U15 ( .A(
        round_inst_sbox_inst0_com_z_inst_n144), .B(
        round_inst_sbox_inst0_com_z_inst_n146), .ZN(
        round_inst_sbox_inst0_com_z_inst_n145) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U14 ( .A(
        round_inst_sbox_inst0_com_z_inst_n210), .B(
        round_inst_sbox_inst0_com_z_inst_n229), .Z(
        round_inst_sbox_inst0_com_z_inst_n146) );
  INV_X1 round_inst_sbox_inst0_com_z_inst_U13 ( .A(
        round_inst_sbox_inst0_com_z_inst_n202), .ZN(
        round_inst_sbox_inst0_com_z_inst_n229) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U12 ( .A1(round_inst_n70), .A2(
        round_inst_sin_w[0]), .ZN(round_inst_sbox_inst0_com_z_inst_n202) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U11 ( .A1(round_inst_sin_w[0]), 
        .A2(round_inst_sin_y[1]), .ZN(round_inst_sbox_inst0_com_z_inst_n210)
         );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U10 ( .A(
        round_inst_sbox_inst0_com_z_inst_n251), .B(
        round_inst_sbox_inst0_com_z_inst_n148), .Z(
        round_inst_sbox_inst0_com_z_inst_n144) );
  INV_X1 round_inst_sbox_inst0_com_z_inst_U9 ( .A(
        round_inst_sbox_inst0_com_z_inst_n156), .ZN(
        round_inst_sbox_inst0_com_z_inst_n148) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U8 ( .A1(round_inst_sin_x[0]), 
        .A2(round_inst_sin_w[3]), .ZN(round_inst_sbox_inst0_com_z_inst_n156)
         );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U7 ( .A1(round_inst_sin_w[0]), 
        .A2(round_inst_sbox_inst0_com_z_inst_n170), .ZN(
        round_inst_sbox_inst0_com_z_inst_n251) );
  INV_X1 round_inst_sbox_inst0_com_z_inst_U6 ( .A(
        round_inst_sbox_inst0_com_z_inst_n242), .ZN(
        round_inst_sbox_inst0_com_z_inst_n170) );
  XOR2_X1 round_inst_sbox_inst0_com_z_inst_U5 ( .A(round_inst_n40), .B(
        round_inst_sbox_inst0_com_z_inst_n169), .Z(
        round_inst_sbox_inst0_com_z_inst_n242) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U4 ( .A(round_inst_sin_w[3]), .B(
        round_inst_sin_x[3]), .ZN(round_inst_sbox_inst0_com_z_inst_n169) );
  XNOR2_X1 round_inst_sbox_inst0_com_z_inst_U3 ( .A(
        round_inst_sbox_inst0_com_z_inst_n209), .B(
        round_inst_sbox_inst0_com_z_inst_n217), .ZN(
        round_inst_sbox_inst0_com_z_inst_n222) );
  AND2_X1 round_inst_sbox_inst0_com_z_inst_U2 ( .A1(round_inst_sin_w[0]), .A2(
        round_inst_sin_x[1]), .ZN(round_inst_sbox_inst0_com_z_inst_n217) );
  NAND2_X1 round_inst_sbox_inst0_com_z_inst_U1 ( .A1(round_inst_n70), .A2(
        round_inst_sin_x[0]), .ZN(round_inst_sbox_inst0_com_z_inst_n209) );
  INV_X1 round_inst_S_1__sbox_inst_U2 ( .A(round_inst_sin_z[5]), .ZN(
        round_inst_S_1__sbox_inst_n2) );
  INV_X2 round_inst_S_1__sbox_inst_U1 ( .A(round_inst_S_1__sbox_inst_n2), .ZN(
        round_inst_S_1__sbox_inst_n1) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U148 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n538), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n537), .ZN(round_inst_sout_w[7])
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U147 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n536), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n535), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n537) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U146 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n534), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n533), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n535) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U145 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n531), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n536) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U144 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U143 ( .A1(round_inst_sin_z[6]), .A2(round_inst_S_1__sbox_inst_com_w_inst_n528), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U142 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n533), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n528) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n526), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n525), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n524), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n523), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n525) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U139 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n521), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n523) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n519), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n521) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U137 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n518), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n519) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n516), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n520) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n514), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n516) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n513), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n512), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n522) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U133 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n514), .A2(round_inst_sin_y[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n511), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n514) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U131 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n517), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n513) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U130 ( .A(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n509) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U129 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n508), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n507), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n524) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U128 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n508) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U127 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U126 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n503), .B(round_inst_sin_z[3]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n504) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U125 ( .A(round_inst_sin_x[5]), 
        .B(round_inst_n40), .ZN(round_inst_S_1__sbox_inst_com_w_inst_n503) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n502), .A2(round_inst_sin_z[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n505) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n501), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n500), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n502) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U122 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n499), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n498), .ZN(round_inst_sout_w[5])
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U121 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n496), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n498) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U120 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n496) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U119 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n493), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n492), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n510), .B(round_inst_sin_z[6]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n491), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n490), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n491) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U115 ( .A(round_inst_sin_y[1]), 
        .B(round_inst_sin_z[1]), .ZN(round_inst_S_1__sbox_inst_com_w_inst_n490) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n526), .ZN(round_inst_sout_w[4])
         );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U113 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n488), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n501), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n526) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n494), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n500), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n500) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U110 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n485), .A2(round_inst_n41), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n486) );
  AND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U109 ( .A1(round_inst_sin_x[6]), 
        .A2(round_inst_S_1__sbox_inst_com_w_inst_n484), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n487) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n483), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n482), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n482) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U106 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n479), .A2(round_inst_sin_z[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n480) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U105 ( .A1(round_inst_sin_x[5]), .A2(round_inst_sin_z[6]), .ZN(round_inst_S_1__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U104 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n478), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n477), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n481) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U103 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n510), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n477) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n475), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n474), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U101 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n473), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n472), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U100 ( .A1(
        round_inst_S_1__sbox_inst_n1), .A2(round_inst_sin_y[4]), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n472) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U99 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n471), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n470), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n478) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U98 ( .A(round_inst_sin_z[4]), 
        .B(round_inst_S_1__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n470) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n469), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n468), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n483) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U96 ( .A1(round_inst_sin_z[6]), 
        .A2(round_inst_S_1__sbox_inst_com_w_inst_n467), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n468) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n466), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n465), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n469) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U94 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n464), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n463), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n465) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U93 ( .A1(round_inst_sin_z[4]), 
        .A2(round_inst_S_1__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n463) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n461), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n460), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n462) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n460) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n458), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n457), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n464) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n517), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U88 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n492), .A2(round_inst_n41), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n517) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U87 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n455), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n454), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n466) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U85 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n474), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n534), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n452) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U84 ( .A(round_inst_n41), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n534) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U83 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n507), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n453) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U82 ( .A1(round_inst_sin_y[4]), 
        .A2(round_inst_sin_x[6]), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n507) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n450), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n489) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U80 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n449), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n448), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n450) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U79 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n447), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n448) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U78 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n446), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n501) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U77 ( .A(round_inst_sin_z[0]), 
        .B(round_inst_sin_y[0]), .ZN(round_inst_S_1__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n445), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n444), .ZN(round_inst_xin_w[7])
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n443), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n442), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n444) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n492), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n451), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n442) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U73 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n441), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n451) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U72 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n439), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n492), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n440) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U71 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U70 ( .A(
        round_inst_S_1__sbox_inst_n1), .B(round_inst_sin_x[5]), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n438) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U69 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n467), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n533), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n441) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n485), .A2(round_inst_sin_y[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n533) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U67 ( .A(round_inst_sin_y[2]), 
        .B(round_inst_sin_z[2]), .Z(round_inst_S_1__sbox_inst_com_w_inst_n443)
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n538), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n445) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n437), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n436), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n435), .A2(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n434), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n433), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n435) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U62 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n471), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n461), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n433) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U61 ( .A1(
        round_inst_S_1__sbox_inst_n1), .A2(round_inst_sin_x[6]), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U60 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n431), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n437) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U59 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n430), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n429), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n431) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U58 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n506), .A2(round_inst_sin_x[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n429) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U57 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n485), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n484), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n506) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U56 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n428), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n427), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n430) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U55 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n426), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n425), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U54 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n423), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n425) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n422), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n421), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n423) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U52 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n518), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n461), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U51 ( .A1(round_inst_sin_x[5]), 
        .A2(round_inst_n41), .ZN(round_inst_S_1__sbox_inst_com_w_inst_n461) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U50 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n455), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n420), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n422) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U49 ( .A(round_inst_n41), .B(
        round_inst_sin_z[6]), .ZN(round_inst_S_1__sbox_inst_com_w_inst_n455)
         );
  NAND3_X1 round_inst_S_1__sbox_inst_com_w_inst_U48 ( .A1(round_inst_sin_y[7]), 
        .A2(round_inst_sin_x[6]), .A3(
        round_inst_S_1__sbox_inst_com_w_inst_n419), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n424) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_w_inst_U47 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n485), .A2(round_inst_n41), .A3(
        round_inst_S_1__sbox_inst_n1), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n426) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U46 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n518), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n471), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n428) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U45 ( .A1(round_inst_sin_x[5]), 
        .A2(round_inst_sin_x[6]), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n471) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U44 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n418), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n417), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U43 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n416), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n415), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n417) );
  NOR3_X1 round_inst_S_1__sbox_inst_com_w_inst_U42 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n414), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n459), .A3(
        round_inst_S_1__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n415) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U41 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n485), .A2(round_inst_sin_x[6]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n447) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U40 ( .A(round_inst_sin_y[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n459) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n510), .A2(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n414) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U38 ( .A(round_inst_sin_x[6]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n510) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_w_inst_U37 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n485), .A2(round_inst_sin_x[6]), 
        .A3(round_inst_S_1__sbox_inst_n1), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n416) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_w_inst_U36 ( .A1(round_inst_sin_x[5]), 
        .A2(round_inst_sin_z[6]), .A3(round_inst_sin_y[7]), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n418) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n538) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U34 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n412) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U33 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n515), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n454), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n410) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U32 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n485), .B(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n515) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U31 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n456), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n527), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n411) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U30 ( .A1(round_inst_sin_y[7]), 
        .A2(round_inst_S_1__sbox_inst_com_w_inst_n492), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n527) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U29 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n419), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n456) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U28 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n408), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n413) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U27 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n407), .A2(round_inst_sin_z[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n408) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U26 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n420), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U25 ( .A1(round_inst_sin_x[5]), 
        .A2(round_inst_S_1__sbox_inst_com_w_inst_n484), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n406) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U24 ( .A(round_inst_sin_y[7]), 
        .B(round_inst_n39), .Z(round_inst_S_1__sbox_inst_com_w_inst_n484) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U23 ( .A1(round_inst_sin_y[5]), 
        .A2(round_inst_S_1__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U22 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n405), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n404), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U21 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n402), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U20 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n401), .A2(round_inst_sin_y[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n402) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U19 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n454), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n401) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U18 ( .A1(round_inst_sin_x[5]), 
        .A2(round_inst_S_1__sbox_inst_com_w_inst_n492), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n454) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U17 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n400), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n403) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n399), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n398), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n400) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U15 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n473), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n397), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n398) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U14 ( .A1(round_inst_sin_z[4]), 
        .A2(round_inst_sin_x[5]), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n397) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U13 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n419), .A2(round_inst_sin_y[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n399) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U12 ( .A(round_inst_sin_y[5]), 
        .B(round_inst_S_1__sbox_inst_n1), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n419) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U11 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n396), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n395), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U10 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n467), .A2(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n395) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U9 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_1__sbox_inst_com_w_inst_n473), .Z(
        round_inst_S_1__sbox_inst_com_w_inst_n467) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U8 ( .A1(round_inst_sin_y[5]), 
        .A2(round_inst_S_1__sbox_inst_com_w_inst_n492), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n473) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U7 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n492) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U6 ( .A(round_inst_sin_x[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n511) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U5 ( .A1(
        round_inst_S_1__sbox_inst_com_w_inst_n518), .A2(
        round_inst_S_1__sbox_inst_com_w_inst_n474), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n396) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_w_inst_U4 ( .A1(round_inst_sin_x[5]), 
        .A2(round_inst_sin_y[4]), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n485), .B(round_inst_sin_y[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n518) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U2 ( .A(
        round_inst_S_1__sbox_inst_com_w_inst_n446), .ZN(
        round_inst_S_1__sbox_inst_com_w_inst_n485) );
  INV_X1 round_inst_S_1__sbox_inst_com_w_inst_U1 ( .A(round_inst_sin_x[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U136 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n512), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n511), .ZN(round_inst_sout_x[4])
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n510), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n509), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n511) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U134 ( .A(round_inst_n41), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U133 ( .A(round_inst_sin_z[0]), 
        .B(round_inst_S_1__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n510) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U132 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n512), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n506), .Z(round_inst_srout2_x[38]) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U130 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n503), .A2(round_inst_sin_z[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U129 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U127 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n498), .A2(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U126 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U125 ( .A1(round_inst_n41), 
        .A2(round_inst_sin_w[4]), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U124 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U122 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U121 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U118 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n508), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n487) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U115 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n481) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_x_inst_U114 ( .A1(round_inst_sin_z[6]), .A2(round_inst_sin_w[4]), .A3(round_inst_S_1__sbox_inst_com_x_inst_n508), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n489) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n478), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n475), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n477) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n474), .B(round_inst_sin_z[3]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n475) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_x_inst_U110 ( .A1(round_inst_sin_w[6]), .A2(round_inst_S_1__sbox_inst_com_x_inst_n508), .A3(round_inst_sin_z[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n473), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n478) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n470), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n473) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n468), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n512) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n467), .A2(round_inst_n41), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n468) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n467) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n469) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n465), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n463), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_srout2_x[36]) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U100 ( .A1(round_inst_sin_y[4]), .A2(round_inst_sin_z[6]), .ZN(round_inst_S_1__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[1]), 
        .B(round_inst_S_1__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n461), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n462) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n466), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n460) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n458), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n457), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_1__sbox_inst_n1), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n459), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n456), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n455), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n454), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n453), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n455) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n452), .A2(round_inst_sin_w[6]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n451), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n450), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n454) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n449), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n448), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n447), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n446), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n448) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n445), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n446) );
  MUX2_X1 round_inst_S_1__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n444), .B(round_inst_n41), .S(
        round_inst_sin_y[4]), .Z(round_inst_S_1__sbox_inst_com_x_inst_n445) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n443), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_1__sbox_inst_com_x_inst_U85 ( .A(round_inst_n41), .B(
        round_inst_sin_z[6]), .S(round_inst_sin_z[4]), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n443) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n442), .A2(round_inst_sin_w[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n449) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n441), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n440), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n451) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_w[4]), 
        .A3(round_inst_sin_z[6]), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n440) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n439), .A2(round_inst_sin_w[5]), 
        .A3(round_inst_n41), .ZN(round_inst_S_1__sbox_inst_com_x_inst_n441) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U80 ( .A(round_inst_sin_y[4]), 
        .B(round_inst_sin_z[4]), .Z(round_inst_S_1__sbox_inst_com_x_inst_n439)
         );
  NAND3_X1 round_inst_S_1__sbox_inst_com_x_inst_U79 ( .A1(round_inst_sin_y[4]), 
        .A2(round_inst_S_1__sbox_inst_com_x_inst_n444), .A3(
        round_inst_S_1__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n456) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n459) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U77 ( .A1(round_inst_sin_y[4]), 
        .A2(round_inst_n41), .ZN(round_inst_S_1__sbox_inst_com_x_inst_n482) );
  AND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U76 ( .A1(round_inst_n41), .A2(
        round_inst_sin_z[4]), .ZN(round_inst_S_1__sbox_inst_com_x_inst_n490)
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n461) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U74 ( .A1(round_inst_sin_y[4]), 
        .A2(round_inst_sin_w[6]), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n497) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n436), .ZN(
        round_inst_srout2_x[39]) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n435), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n434), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n436) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U71 ( .A(round_inst_sin_y[4]), 
        .B(round_inst_S_1__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n434) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n433), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n432), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U69 ( .A1(round_inst_sin_z[4]), 
        .A2(round_inst_S_1__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n432) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n431), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n430), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n433) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n429), .A2(round_inst_sin_y[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n428), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n427) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_1__sbox_inst_n1), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n431) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n452) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[2]), 
        .B(round_inst_S_1__sbox_inst_com_x_inst_n437), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n435) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n424), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n423), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n422), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n421), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n423) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n420), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n419), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n421) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n418), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n419) );
  NOR3_X1 round_inst_S_1__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n470), .A3(
        round_inst_S_1__sbox_inst_com_x_inst_n416), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n417) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n415), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n414), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n418) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n413), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n414) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U53 ( .A1(round_inst_n41), 
        .A2(round_inst_S_1__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n412) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U52 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n442), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_1__sbox_inst_n1), .A2(round_inst_n41), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n442) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_x_inst_U50 ( .A1(round_inst_n41), 
        .A2(round_inst_S_1__sbox_inst_com_x_inst_n476), .A3(
        round_inst_S_1__sbox_inst_com_x_inst_n411), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n420) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U49 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n410), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n422) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U48 ( .A1(round_inst_n41), 
        .A2(round_inst_n39), .ZN(round_inst_S_1__sbox_inst_com_x_inst_n464) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U47 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n410) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n409), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n407), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n406), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n405), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n404), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n406) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U43 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n465), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n404) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U42 ( .A(round_inst_sin_w[5]), 
        .B(round_inst_S_1__sbox_inst_n1), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n438) );
  AND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U41 ( .A1(round_inst_sin_z[6]), 
        .A2(round_inst_S_1__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n465) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U40 ( .A1(round_inst_n39), 
        .A2(round_inst_S_1__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n405) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n476), .A3(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n407) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U38 ( .A(round_inst_sin_z[6]), 
        .B(round_inst_sin_w[6]), .Z(round_inst_S_1__sbox_inst_com_x_inst_n444)
         );
  NOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U37 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n403), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n402), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U36 ( .A(round_inst_sin_w[6]), 
        .B(round_inst_n41), .Z(round_inst_S_1__sbox_inst_com_x_inst_n402) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U35 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n401), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n400), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n399), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n400) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U33 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n398) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U32 ( .A1(round_inst_sin_z[4]), 
        .A2(round_inst_S_1__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n425) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U31 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n479), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n471) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n508), .B(round_inst_n39), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n426), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n399) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U28 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n401) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_1__sbox_inst_n1), .A3(round_inst_sin_y[4]), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n396) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n411), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U23 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n392), .A2(round_inst_sin_w[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U21 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_x_inst_U19 ( .A1(round_inst_sin_z[4]), 
        .A2(round_inst_S_1__sbox_inst_com_x_inst_n508), .A3(
        round_inst_sin_w[5]), .ZN(round_inst_S_1__sbox_inst_com_x_inst_n388)
         );
  MUX2_X1 round_inst_S_1__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n411), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n508), .S(
        round_inst_S_1__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U17 ( .A1(round_inst_sin_y[4]), 
        .A2(round_inst_S_1__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n491), .B(round_inst_n39), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n411) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U15 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U14 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n384), .A2(round_inst_sin_z[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n403), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U10 ( .A(round_inst_sin_w[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U9 ( .A1(
        round_inst_S_1__sbox_inst_n1), .A2(
        round_inst_S_1__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n403) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U8 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n508) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U7 ( .A(round_inst_sin_y[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n413) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n382), .A2(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_1__sbox_inst_com_x_inst_n426), .Z(
        round_inst_S_1__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U4 ( .A1(round_inst_sin_y[4]), 
        .A2(round_inst_sin_w[5]), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n426) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_1__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_w[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_1__sbox_inst_com_x_inst_n416), .ZN(
        round_inst_S_1__sbox_inst_com_x_inst_n476) );
  INV_X1 round_inst_S_1__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_y[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_x_inst_n416) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n517), .Z(round_inst_sout_y[4])
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n516), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n514), .B(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n515) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U134 ( .A(round_inst_sin_x[0]), 
        .B(round_inst_S_1__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n512), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_srout2_y[38]) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n508), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n518) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n507), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n506), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n508) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n506) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n503), .A2(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n507) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_1__sbox_inst_com_y_inst_U125 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_1__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U124 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U123 ( .A1(round_inst_sin_x[7]), .A2(round_inst_S_1__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n492), .A2(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U121 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U120 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U119 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U118 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n486), .A2(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U117 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n503), .A2(round_inst_sin_w[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U112 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_1__sbox_inst_n1), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[3]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_y_inst_U109 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n514), .A2(round_inst_n39), .A3(
        round_inst_sin_x[4]), .ZN(round_inst_S_1__sbox_inst_com_y_inst_n476)
         );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U108 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_y_inst_U107 ( .A1(round_inst_sin_w[4]), .A2(round_inst_sin_w[7]), .A3(round_inst_S_1__sbox_inst_com_y_inst_n514), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_1__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_1__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U105 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[36]) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U104 ( .A1(round_inst_sin_x[6]), .A2(round_inst_S_1__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U98 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_1__sbox_inst_n1), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U95 ( .A1(round_inst_sin_x[4]), 
        .A2(round_inst_S_1__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_y_inst_U94 ( .A1(round_inst_sin_w[4]), 
        .A2(round_inst_sin_x[5]), .A3(
        round_inst_S_1__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U93 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U92 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n457), .A2(round_inst_sin_x[6]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U88 ( .A1(
        round_inst_S_1__sbox_inst_n1), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_1__sbox_inst_com_y_inst_U87 ( .A(round_inst_sin_x[6]), 
        .B(round_inst_S_1__sbox_inst_com_y_inst_n503), .S(
        round_inst_S_1__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_1__sbox_inst_n1), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n478), .B(round_inst_sin_x[1]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n438), .Z(round_inst_srout2_y[39]) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U71 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U70 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_x[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_1__sbox_inst_n1), .A2(round_inst_sin_w[4]), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[7]), 
        .A3(round_inst_S_1__sbox_inst_n1), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U66 ( .A(round_inst_sin_w[4]), 
        .B(round_inst_sin_x[4]), .Z(round_inst_S_1__sbox_inst_com_y_inst_n443)
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U59 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U58 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U55 ( .A(round_inst_sin_x[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U54 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n418), .A2(round_inst_n39), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U53 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U51 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U50 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n414), .B(round_inst_sin_x[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U49 ( .A(round_inst_sin_w[5]), 
        .B(round_inst_S_1__sbox_inst_n1), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U48 ( .A1(
        round_inst_S_1__sbox_inst_n1), .A2(round_inst_sin_x[4]), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_1__sbox_inst_n1), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U46 ( .A(round_inst_sin_x[2]), 
        .B(round_inst_S_1__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n513) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[5]), 
        .B(round_inst_sin_x[7]), .Z(round_inst_S_1__sbox_inst_com_y_inst_n409)
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U41 ( .A(round_inst_sin_x[5]), 
        .B(round_inst_S_1__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[4]), 
        .Z(round_inst_S_1__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U36 ( .A(round_inst_sin_z[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_1__sbox_inst_n1), .B(round_inst_n39), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U28 ( .A(round_inst_sin_x[6]), 
        .B(round_inst_S_1__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U27 ( .A1(round_inst_sin_w[5]), 
        .A2(round_inst_n39), .ZN(round_inst_S_1__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n514), .A2(round_inst_sin_w[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_1__sbox_inst_n1), .A2(round_inst_sin_w[7]), .A3(
        round_inst_sin_x[6]), .ZN(round_inst_S_1__sbox_inst_com_y_inst_n403)
         );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_1__sbox_inst_n1), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n504), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_1__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U18 ( .A(round_inst_n39), .B(
        round_inst_sin_w[7]), .ZN(round_inst_S_1__sbox_inst_com_y_inst_n395)
         );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U17 ( .A(round_inst_n39), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[7]), 
        .B(round_inst_sin_x[7]), .ZN(round_inst_S_1__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_y_inst_U13 ( .A1(round_inst_sin_x[5]), 
        .A2(round_inst_sin_w[7]), .A3(
        round_inst_S_1__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_y_inst_U12 ( .A1(round_inst_n39), 
        .A2(round_inst_S_1__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_1__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[5]), 
        .B(round_inst_sin_x[5]), .S(round_inst_S_1__sbox_inst_com_y_inst_n503), 
        .Z(round_inst_S_1__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_1__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_y_inst_U9 ( .A1(round_inst_sin_x[5]), 
        .A2(round_inst_S_1__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_1__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U8 ( .A(round_inst_n39), .B(
        round_inst_sin_x[7]), .Z(round_inst_S_1__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_1__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_1__sbox_inst_n1), .A3(round_inst_sin_x[7]), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_1__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n503) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[6]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_1__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_1__sbox_inst_com_y_inst_n514) );
  INV_X1 round_inst_S_1__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[6]), 
        .ZN(round_inst_S_1__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U132 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n517), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n516), .ZN(round_inst_sout_z[4])
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n515), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n514), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U130 ( .A(round_inst_sin_w[6]), 
        .B(round_inst_sin_w[7]), .ZN(round_inst_S_1__sbox_inst_com_z_inst_n514) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_x[0]), 
        .B(round_inst_sin_y[0]), .Z(round_inst_S_1__sbox_inst_com_z_inst_n515)
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U128 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n512), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n517) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_srout2_z[38]) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n510), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n509), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n511) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n508), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n507), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n509) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U124 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n506), .A2(round_inst_sin_y[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U123 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n505), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n504), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n508) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n503), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n502), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U121 ( .A(round_inst_sin_w[5]), 
        .B(round_inst_sin_x[3]), .ZN(round_inst_S_1__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U120 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n501), .B(round_inst_n40), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n503) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U119 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n500), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n499), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n501) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U118 ( .A1(round_inst_n41), 
        .A2(round_inst_S_1__sbox_inst_com_z_inst_n498), .A3(
        round_inst_S_1__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n499) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U117 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_x[4]), 
        .A3(round_inst_sin_w[7]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n500) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U116 ( .A(round_inst_sin_x[6]), 
        .B(round_inst_n41), .Z(round_inst_S_1__sbox_inst_com_z_inst_n496) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U115 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n497), .A2(round_inst_sin_x[6]), 
        .A3(round_inst_sin_x[7]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n505) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U114 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n495), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n494), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n493), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n492), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n494) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n491), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n490), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n492) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U111 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n489), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n488), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n490) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n487), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n491) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U109 ( .A1(round_inst_sin_w[6]), .A2(round_inst_sin_x[7]), .A3(round_inst_sin_y[4]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n493) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U108 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n485), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n513) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U107 ( .A1(round_inst_sin_w[6]), .A2(round_inst_S_1__sbox_inst_com_z_inst_n498), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n486) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U106 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n484), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n506), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n482), .Z(round_inst_srout2_z[36]) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n481), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n480), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n479), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n484), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n478), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n477), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n484) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U101 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n476), .A2(round_inst_sin_x[4]), 
        .A3(round_inst_sin_w[6]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n477) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U100 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n475), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n474), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n478) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U99 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n473), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n497), .A3(round_inst_n41), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n474) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U98 ( .A(round_inst_sin_w[5]), 
        .B(round_inst_sin_y[5]), .Z(round_inst_S_1__sbox_inst_com_z_inst_n473)
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U97 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n472), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n471), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n475) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U96 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n470), .A2(round_inst_sin_x[6]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n471) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U95 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n469), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n468), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n467), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n466), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n465), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n464), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n466) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n463), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n462), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U91 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n461), .A2(round_inst_n41), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n462) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U90 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n460), .A2(round_inst_sin_x[6]), 
        .A3(round_inst_S_1__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n463) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U89 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n459), .A2(round_inst_sin_y[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n465) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_w[6]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U87 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n469) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U85 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n453), .A2(round_inst_n41), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n454) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U84 ( .A(round_inst_sin_w[5]), 
        .B(round_inst_S_1__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U83 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n451), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U82 ( .A1(round_inst_sin_w[6]), 
        .A2(round_inst_sin_x[4]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U81 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n488), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n448) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U79 ( .A(round_inst_sin_y[1]), 
        .B(round_inst_sin_x[1]), .Z(round_inst_S_1__sbox_inst_com_z_inst_n447)
         );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U78 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n497), .A2(round_inst_sin_x[6]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n488) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n446), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n483) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U76 ( .A(round_inst_sin_w[6]), 
        .B(round_inst_n41), .ZN(round_inst_S_1__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U75 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_srout2_z[39]) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n495), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n512), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U72 ( .A1(round_inst_sin_x[4]), 
        .A2(round_inst_sin_w[7]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n441) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U71 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n458), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n440), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n442) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U70 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n498), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U69 ( .A(round_inst_sin_w[7]), 
        .B(round_inst_S_1__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n498) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U68 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n495) );
  MUX2_X1 round_inst_S_1__sbox_inst_com_z_inst_U67 ( .A(round_inst_sin_x[7]), 
        .B(round_inst_sin_w[7]), .S(round_inst_S_1__sbox_inst_com_z_inst_n436), 
        .Z(round_inst_S_1__sbox_inst_com_z_inst_n437) );
  OR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U66 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n436) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U65 ( .A(round_inst_sin_x[4]), 
        .B(round_inst_S_1__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n487) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U64 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n438) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U63 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n497), .A2(round_inst_sin_x[7]), 
        .A3(round_inst_S_1__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U62 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n430), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n429) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U59 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n426), .A2(round_inst_sin_w[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U58 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n422), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n424) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U56 ( .A1(round_inst_sin_x[4]), 
        .A2(round_inst_S_1__sbox_inst_com_z_inst_n460), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U55 ( .A1(round_inst_sin_y[5]), 
        .A2(round_inst_sin_x[4]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n425) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U54 ( .A1(round_inst_sin_y[4]), 
        .A2(round_inst_sin_x[7]), .A3(round_inst_sin_w[5]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n428) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U53 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_y[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U52 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n461), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n423), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n470) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U50 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n497), .A2(round_inst_sin_y[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n423) );
  AND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U49 ( .A1(round_inst_sin_w[5]), 
        .A2(round_inst_sin_x[4]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n461) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U48 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n421) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U47 ( .A1(round_inst_sin_w[5]), 
        .A2(round_inst_S_1__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U46 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n460), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n419), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n418), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n432) );
  INV_X1 round_inst_S_1__sbox_inst_com_z_inst_U44 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U43 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n497), .B(round_inst_sin_y[4]), 
        .Z(round_inst_S_1__sbox_inst_com_z_inst_n451) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n417), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U41 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n497), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n449) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U39 ( .A1(round_inst_sin_w[7]), 
        .A2(round_inst_S_1__sbox_inst_com_z_inst_n413), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n414) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U38 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n415) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U35 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n506), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n460), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n409) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U34 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n407) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U32 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n405) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n404) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U30 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n506), .A2(round_inst_sin_y[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n402) );
  AND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U29 ( .A1(round_inst_sin_x[6]), 
        .A2(round_inst_sin_w[7]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n506) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n401), .A2(round_inst_n41), .A3(
        round_inst_sin_w[5]), .ZN(round_inst_S_1__sbox_inst_com_z_inst_n403)
         );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U27 ( .A(round_inst_sin_w[7]), 
        .B(round_inst_sin_x[7]), .Z(round_inst_S_1__sbox_inst_com_z_inst_n401)
         );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U26 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n399), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n406) );
  MUX2_X1 round_inst_S_1__sbox_inst_com_z_inst_U25 ( .A(round_inst_sin_y[7]), 
        .B(round_inst_S_1__sbox_inst_com_z_inst_n398), .S(
        round_inst_S_1__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U24 ( .A1(round_inst_sin_w[5]), 
        .A2(round_inst_sin_x[6]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U23 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n398) );
  INV_X1 round_inst_S_1__sbox_inst_com_z_inst_U22 ( .A(round_inst_sin_x[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n397) );
  NOR3_X1 round_inst_S_1__sbox_inst_com_z_inst_U21 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n489), .A3(
        round_inst_S_1__sbox_inst_com_z_inst_n395), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U20 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n394), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n395) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U19 ( .A(round_inst_sin_w[7]), 
        .B(round_inst_sin_y[7]), .ZN(round_inst_S_1__sbox_inst_com_z_inst_n489) );
  AND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U18 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n459), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U17 ( .A1(round_inst_sin_w[6]), 
        .A2(round_inst_S_1__sbox_inst_com_z_inst_n460), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n459) );
  INV_X1 round_inst_S_1__sbox_inst_com_z_inst_U16 ( .A(round_inst_sin_w[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U15 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n393), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U14 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n391), .A2(round_inst_n41), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U13 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_1__sbox_inst_com_z_inst_n390), .Z(
        round_inst_S_1__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U12 ( .A1(round_inst_sin_w[5]), 
        .A2(round_inst_sin_y[7]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n390) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U11 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n460), .A2(round_inst_sin_w[7]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n418) );
  NOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U10 ( .A1(
        round_inst_S_1__sbox_inst_com_z_inst_n439), .A2(
        round_inst_S_1__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_1__sbox_inst_com_z_inst_U9 ( .A1(round_inst_sin_w[6]), 
        .A2(round_inst_sin_w[5]), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n456) );
  XNOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U8 ( .A(round_inst_sin_x[7]), 
        .B(round_inst_sin_y[7]), .ZN(round_inst_S_1__sbox_inst_com_z_inst_n439) );
  NAND3_X1 round_inst_S_1__sbox_inst_com_z_inst_U7 ( .A1(round_inst_sin_w[6]), 
        .A2(round_inst_sin_x[7]), .A3(
        round_inst_S_1__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U6 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n460), .B(round_inst_sin_y[5]), 
        .Z(round_inst_S_1__sbox_inst_com_z_inst_n476) );
  INV_X1 round_inst_S_1__sbox_inst_com_z_inst_U5 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n394), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n460) );
  INV_X1 round_inst_S_1__sbox_inst_com_z_inst_U4 ( .A(round_inst_sin_x[5]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n394) );
  INV_X1 round_inst_S_1__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_1__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_1__sbox_inst_com_z_inst_n497) );
  INV_X1 round_inst_S_1__sbox_inst_com_z_inst_U2 ( .A(round_inst_sin_w[4]), 
        .ZN(round_inst_S_1__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_1__sbox_inst_com_z_inst_U1 ( .A(round_inst_sin_y[2]), 
        .B(round_inst_sin_x[2]), .Z(round_inst_S_1__sbox_inst_com_z_inst_n417)
         );
  INV_X1 round_inst_S_2__sbox_inst_U6 ( .A(round_inst_sin_x[10]), .ZN(
        round_inst_S_2__sbox_inst_n6) );
  INV_X1 round_inst_S_2__sbox_inst_U5 ( .A(round_inst_sin_z[9]), .ZN(
        round_inst_S_2__sbox_inst_n2) );
  INV_X1 round_inst_S_2__sbox_inst_U4 ( .A(round_inst_sin_z[11]), .ZN(
        round_inst_S_2__sbox_inst_n4) );
  INV_X2 round_inst_S_2__sbox_inst_U3 ( .A(round_inst_S_2__sbox_inst_n4), .ZN(
        round_inst_S_2__sbox_inst_n3) );
  INV_X2 round_inst_S_2__sbox_inst_U2 ( .A(round_inst_S_2__sbox_inst_n2), .ZN(
        round_inst_S_2__sbox_inst_n1) );
  INV_X2 round_inst_S_2__sbox_inst_U1 ( .A(round_inst_S_2__sbox_inst_n6), .ZN(
        round_inst_S_2__sbox_inst_n5) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n531), .ZN(round_inst_sout_w[11])
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U139 ( .A1(round_inst_sin_z[8]), .A2(round_inst_S_2__sbox_inst_com_w_inst_n528), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n526), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n524), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n526) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[10]), .A2(round_inst_S_2__sbox_inst_com_w_inst_n523), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n525) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n518), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n516), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n518) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n514), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n513), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n512), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n513) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_w_inst_U128 ( .A1(
        round_inst_S_2__sbox_inst_n5), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n510), .A3(
        round_inst_S_2__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n511) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U127 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n508), .A2(round_inst_n42), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n507), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U125 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n507) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_2__sbox_inst_n3), .A2(round_inst_n43), .A3(
        round_inst_S_2__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U122 ( .A(round_inst_sin_y[7]), 
        .B(round_inst_S_2__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U121 ( .A(round_inst_n61), .B(
        round_inst_n39), .Z(round_inst_S_2__sbox_inst_com_w_inst_n501) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U120 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[9])
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[5]), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[5]), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U113 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[8])
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_2__sbox_inst_n5), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U110 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n528), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U105 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_2__sbox_inst_n5), .B(round_inst_sin_z[10]), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_2__sbox_inst_n1), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U99 ( .A1(round_inst_n43), 
        .A2(round_inst_S_2__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_2__sbox_inst_n5), .A2(round_inst_n42), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n506) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U94 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[10]), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n461), .A2(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[10]), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U88 ( .A1(round_inst_sin_z[8]), 
        .A2(round_inst_S_2__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_w_inst_U85 ( .A1(round_inst_sin_y[9]), 
        .A2(round_inst_n42), .A3(round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_w_inst_U84 ( .A1(round_inst_n43), 
        .A2(round_inst_n61), .A3(round_inst_n42), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n528) );
  OR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_2__sbox_inst_n5), .B(round_inst_n43), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U80 ( .A(round_inst_sin_y[4]), 
        .B(round_inst_sin_z[4]), .Z(round_inst_S_2__sbox_inst_com_w_inst_n484)
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U79 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[11])
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U73 ( .A1(
        round_inst_S_2__sbox_inst_n3), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U71 ( .A1(round_inst_n43), 
        .A2(round_inst_n61), .ZN(round_inst_S_2__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_2__sbox_inst_n5), .A2(round_inst_sin_y[9]), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U69 ( .A1(
        round_inst_S_2__sbox_inst_n1), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n508), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_2__sbox_inst_n5), .A2(round_inst_S_2__sbox_inst_n1), .A3(
        round_inst_S_2__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n439), .A2(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n508), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_2__sbox_inst_n3), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n504) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U62 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n508) );
  INV_X1 round_inst_S_2__sbox_inst_com_w_inst_U61 ( .A(round_inst_n43), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U60 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U58 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U57 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U56 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U55 ( .A(round_inst_sin_y[9]), 
        .B(round_inst_S_2__sbox_inst_n1), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U54 ( .A1(
        round_inst_S_2__sbox_inst_n3), .A2(round_inst_S_2__sbox_inst_n1), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U52 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_w_inst_U51 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n505), .A3(
        round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U50 ( .A(round_inst_sin_y[9]), 
        .B(round_inst_n61), .Z(round_inst_S_2__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_w_inst_U49 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n505), .A2(round_inst_sin_y[9]), 
        .A3(round_inst_S_2__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U48 ( .A(round_inst_n43), .B(
        round_inst_sin_z[10]), .ZN(round_inst_S_2__sbox_inst_com_w_inst_n465)
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U47 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n520) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U45 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n421), .A2(
        round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U44 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U43 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n419), .A2(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U42 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U40 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_2__sbox_inst_n1), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n521) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U38 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U37 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U36 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n510), .B(round_inst_sin_z[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n498), .A2(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U33 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U32 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U31 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U30 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U29 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U28 ( .A1(round_inst_n61), 
        .A2(round_inst_sin_z[8]), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U27 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n522), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U26 ( .A(round_inst_n61), .B(
        round_inst_S_2__sbox_inst_n1), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U24 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n510), .A2(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U22 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[9]), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U21 ( .A(round_inst_n42), .B(
        round_inst_sin_z[8]), .Z(round_inst_S_2__sbox_inst_com_w_inst_n418) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U20 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U19 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U17 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n398), .A2(
        round_inst_S_2__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U15 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n498), .B(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_2__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_2__sbox_inst_com_w_inst_U13 ( .A(round_inst_sin_y[11]), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_2__sbox_inst_n1), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U11 ( .A(
        round_inst_S_2__sbox_inst_n3), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n505), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U9 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_2__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_2__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U8 ( .A1(round_inst_n61), .A2(
        round_inst_n42), .ZN(round_inst_S_2__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U7 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n510), .A2(round_inst_sin_y[9]), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n477) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_w_inst_U6 ( .A1(
        round_inst_S_2__sbox_inst_com_w_inst_n505), .A2(round_inst_n42), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n522) );
  INV_X1 round_inst_S_2__sbox_inst_com_w_inst_U5 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n505) );
  INV_X1 round_inst_S_2__sbox_inst_com_w_inst_U4 ( .A(round_inst_sin_x[11]), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n486) );
  INV_X1 round_inst_S_2__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_2__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_2__sbox_inst_com_w_inst_n510) );
  INV_X1 round_inst_S_2__sbox_inst_com_w_inst_U2 ( .A(round_inst_sin_x[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_w_inst_n489) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_w_inst_U1 ( .A(round_inst_n41), .B(
        round_inst_sin_z[6]), .Z(round_inst_S_2__sbox_inst_com_w_inst_n402) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n510), .ZN(round_inst_sout_x[8])
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n509), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n510) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U133 ( .A(round_inst_n43), .B(
        round_inst_sin_y[11]), .ZN(round_inst_S_2__sbox_inst_com_x_inst_n508)
         );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U132 ( .A(round_inst_sin_z[4]), 
        .B(round_inst_S_2__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n506), .Z(round_inst_srout2_x[58]) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U130 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U129 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n503), .A2(round_inst_sin_z[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U127 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U126 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U125 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U124 ( .A1(round_inst_n43), 
        .A2(round_inst_sin_w[8]), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U122 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U121 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U118 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_sin_y[11]), .A2(round_inst_S_2__sbox_inst_com_x_inst_n490), 
        .ZN(round_inst_S_2__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U115 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n487) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_x_inst_U114 ( .A1(
        round_inst_sin_z[10]), .A2(round_inst_sin_w[8]), .A3(
        round_inst_sin_y[11]), .ZN(round_inst_S_2__sbox_inst_com_x_inst_n489)
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n478), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n476), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n478) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n475), .B(round_inst_n39), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n476) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_w[10]), .A2(round_inst_sin_y[11]), .A3(
        round_inst_sin_z[8]), .ZN(round_inst_S_2__sbox_inst_com_x_inst_n475)
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n474), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n473), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n473) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n470), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n469), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n511) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n468), .A2(round_inst_n43), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n469) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n468) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n467), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n464), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_srout2_x[56]) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U100 ( .A1(round_inst_n42), 
        .A2(round_inst_sin_z[10]), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[5]), 
        .B(round_inst_S_2__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n464) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n462), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n460), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n467), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n461) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n458), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n467) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_2__sbox_inst_n1), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n457), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n459) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n455), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n454), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n456) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n453), .A2(round_inst_sin_w[10]), 
        .ZN(round_inst_S_2__sbox_inst_com_x_inst_n454) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n451), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n455) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n450), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n449), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n451) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n448), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n447), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n449) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n446), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_2__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n445), .B(round_inst_n43), .S(
        round_inst_n42), .Z(round_inst_S_2__sbox_inst_com_x_inst_n446) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n444), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n448) );
  MUX2_X1 round_inst_S_2__sbox_inst_com_x_inst_U85 ( .A(round_inst_n43), .B(
        round_inst_sin_z[10]), .S(round_inst_sin_z[8]), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n443), .A2(round_inst_sin_w[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n442), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n441), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n452) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[8]), 
        .A3(round_inst_sin_z[10]), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n441) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n440), .A2(round_inst_sin_w[9]), 
        .A3(round_inst_n43), .ZN(round_inst_S_2__sbox_inst_com_x_inst_n442) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U80 ( .A(round_inst_n42), .B(
        round_inst_sin_z[8]), .Z(round_inst_S_2__sbox_inst_com_x_inst_n440) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_x_inst_U79 ( .A1(round_inst_n42), 
        .A2(round_inst_S_2__sbox_inst_com_x_inst_n445), .A3(
        round_inst_S_2__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n460) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U77 ( .A1(round_inst_n42), 
        .A2(round_inst_n43), .ZN(round_inst_S_2__sbox_inst_com_x_inst_n482) );
  AND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U76 ( .A1(round_inst_n43), .A2(
        round_inst_sin_z[8]), .ZN(round_inst_S_2__sbox_inst_com_x_inst_n490)
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n462) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U74 ( .A1(round_inst_n42), 
        .A2(round_inst_sin_w[10]), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n497) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_srout2_x[59]) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n436), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n435), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U71 ( .A(round_inst_n42), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n435) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n434), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n433), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U69 ( .A1(round_inst_sin_z[8]), 
        .A2(round_inst_sin_y[11]), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n433) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n432), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n431), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n434) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n430), .A2(round_inst_n42), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n431) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n429), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n428), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_2__sbox_inst_n1), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n453), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n432) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[6]), 
        .B(round_inst_S_2__sbox_inst_com_x_inst_n438), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n436) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n425), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n424), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n423), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n422), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n421), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n420), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n422) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n419), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n420) );
  NOR3_X1 round_inst_S_2__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n471), .A3(
        round_inst_S_2__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n418) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n416), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n419) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n414), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U53 ( .A1(round_inst_n43), 
        .A2(round_inst_S_2__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n413) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U52 ( .A(round_inst_sin_y[11]), 
        .ZN(round_inst_S_2__sbox_inst_com_x_inst_n414) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n443), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n416) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U50 ( .A1(
        round_inst_S_2__sbox_inst_n1), .A2(round_inst_n43), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n443) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_x_inst_U49 ( .A1(round_inst_n43), 
        .A2(round_inst_S_2__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_2__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n421) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n411), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n423) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U47 ( .A1(round_inst_n43), 
        .A2(round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n465) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n411) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n410), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n407), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U43 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n406), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n405), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n407) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U42 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n466), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n405) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U41 ( .A(round_inst_sin_w[9]), 
        .B(round_inst_S_2__sbox_inst_n1), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n439) );
  AND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U40 ( .A1(round_inst_sin_z[10]), 
        .A2(round_inst_sin_y[11]), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_2__sbox_inst_n3), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n406) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_x_inst_U38 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U37 ( .A(round_inst_sin_z[10]), 
        .B(round_inst_sin_w[10]), .Z(round_inst_S_2__sbox_inst_com_x_inst_n445) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U36 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n404), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n410) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U35 ( .A(round_inst_sin_w[10]), 
        .B(round_inst_n43), .Z(round_inst_S_2__sbox_inst_com_x_inst_n403) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n402), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n401), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U33 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n400), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n399), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n401) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U32 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n399) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U31 ( .A1(round_inst_sin_z[8]), 
        .A2(round_inst_S_2__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n426) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n427), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n400) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U28 ( .A(round_inst_sin_y[11]), 
        .B(round_inst_S_2__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n471) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n402) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_2__sbox_inst_n1), .A3(round_inst_n42), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n396) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n398), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n481) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U23 ( .A(round_inst_sin_y[11]), 
        .B(round_inst_S_2__sbox_inst_n3), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U21 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n392), .A2(round_inst_sin_w[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n404), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_x_inst_U17 ( .A1(round_inst_sin_z[8]), 
        .A2(round_inst_sin_y[11]), .A3(round_inst_sin_w[9]), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n388) );
  MUX2_X1 round_inst_S_2__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n412), .B(round_inst_sin_y[11]), 
        .S(round_inst_S_2__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U15 ( .A1(round_inst_n42), 
        .A2(round_inst_S_2__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U14 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n491), .B(
        round_inst_S_2__sbox_inst_n3), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n412) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n384), .A2(round_inst_sin_z[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U10 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_2__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U9 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_w[11]), 
        .ZN(round_inst_S_2__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U7 ( .A1(
        round_inst_S_2__sbox_inst_n1), .A2(round_inst_sin_y[11]), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n404) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_2__sbox_inst_com_x_inst_n427), .Z(
        round_inst_S_2__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U4 ( .A1(round_inst_n42), .A2(
        round_inst_sin_w[9]), .ZN(round_inst_S_2__sbox_inst_com_x_inst_n427)
         );
  NAND2_X1 round_inst_S_2__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_2__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_2__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_2__sbox_inst_com_x_inst_n477) );
  INV_X1 round_inst_S_2__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_y[9]), 
        .ZN(round_inst_S_2__sbox_inst_com_x_inst_n417) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n517), .Z(round_inst_sout_y[8])
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n516), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n515) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U134 ( .A(round_inst_sin_x[4]), 
        .B(round_inst_S_2__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n512), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_srout2_y[58]) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n508), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n518) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n507), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n506), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n508) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n506) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n507) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_2__sbox_inst_com_y_inst_U125 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_2__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U124 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U123 ( .A1(
        round_inst_sin_x[11]), .A2(round_inst_S_2__sbox_inst_com_y_inst_n493), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n492), .A2(
        round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U121 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U120 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U119 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U118 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n486), .A2(
        round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U117 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n503), .A2(round_inst_sin_w[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U112 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_2__sbox_inst_n1), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[7]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_y_inst_U109 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_2__sbox_inst_n3), .A3(round_inst_sin_x[8]), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U108 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_y_inst_U107 ( .A1(round_inst_sin_w[8]), .A2(round_inst_sin_w[11]), .A3(round_inst_S_2__sbox_inst_com_y_inst_n514), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_2__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_2__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U105 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[56]) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U104 ( .A1(
        round_inst_S_2__sbox_inst_n5), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U98 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_2__sbox_inst_n1), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U95 ( .A1(round_inst_sin_x[8]), 
        .A2(round_inst_S_2__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_y_inst_U94 ( .A1(round_inst_sin_w[8]), 
        .A2(round_inst_n61), .A3(round_inst_S_2__sbox_inst_com_y_inst_n514), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U93 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U92 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U88 ( .A1(
        round_inst_S_2__sbox_inst_n1), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_2__sbox_inst_com_y_inst_U87 ( .A(
        round_inst_S_2__sbox_inst_n5), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n503), .S(
        round_inst_S_2__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_2__sbox_inst_n1), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n478), .B(round_inst_sin_x[5]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n438), .Z(round_inst_srout2_y[59]) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U71 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[11]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U70 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n483), .A2(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_2__sbox_inst_n1), .A2(round_inst_sin_w[8]), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[11]), 
        .A3(round_inst_S_2__sbox_inst_n1), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U66 ( .A(round_inst_sin_w[8]), 
        .B(round_inst_sin_x[8]), .Z(round_inst_S_2__sbox_inst_com_y_inst_n443)
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U59 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[11]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U58 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[9]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U55 ( .A(round_inst_sin_x[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U54 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n418), .A2(
        round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U53 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U51 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U50 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n414), .B(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U49 ( .A(round_inst_sin_w[9]), 
        .B(round_inst_S_2__sbox_inst_n1), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U48 ( .A1(
        round_inst_S_2__sbox_inst_n1), .A2(round_inst_sin_x[8]), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_2__sbox_inst_n1), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U46 ( .A(round_inst_sin_x[6]), 
        .B(round_inst_S_2__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n513) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[9]), 
        .B(round_inst_sin_x[11]), .Z(round_inst_S_2__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U41 ( .A(round_inst_n61), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[11]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[8]), 
        .Z(round_inst_S_2__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U36 ( .A(round_inst_sin_z[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_2__sbox_inst_n1), .B(round_inst_S_2__sbox_inst_n3), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_2__sbox_inst_n5), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U27 ( .A1(round_inst_sin_w[9]), 
        .A2(round_inst_S_2__sbox_inst_n3), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n514), .A2(round_inst_sin_w[9]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_2__sbox_inst_n1), .A2(round_inst_sin_w[11]), .A3(
        round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_2__sbox_inst_n1), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n504), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_2__sbox_inst_n3), .B(round_inst_sin_w[11]), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U17 ( .A(
        round_inst_S_2__sbox_inst_n3), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[11]), 
        .B(round_inst_sin_x[11]), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_y_inst_U13 ( .A1(round_inst_n61), 
        .A2(round_inst_sin_w[11]), .A3(
        round_inst_S_2__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_y_inst_U12 ( .A1(
        round_inst_S_2__sbox_inst_n3), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_2__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[9]), 
        .B(round_inst_n61), .S(round_inst_S_2__sbox_inst_com_y_inst_n503), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_y_inst_U9 ( .A1(round_inst_n61), .A2(
        round_inst_S_2__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_2__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_2__sbox_inst_n3), .B(round_inst_sin_x[11]), .Z(
        round_inst_S_2__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_2__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_2__sbox_inst_n1), .A3(round_inst_sin_x[11]), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_2__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n503) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[10]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_2__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_2__sbox_inst_com_y_inst_n514) );
  INV_X1 round_inst_S_2__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[10]), 
        .ZN(round_inst_S_2__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n516), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n515), .ZN(round_inst_sout_z[8])
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n514), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n513), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_w[10]), .B(round_inst_sin_w[11]), .ZN(round_inst_S_2__sbox_inst_com_z_inst_n513) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U128 ( .A(round_inst_sin_x[4]), 
        .B(round_inst_sin_y[4]), .Z(round_inst_S_2__sbox_inst_com_z_inst_n514)
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n510), .ZN(
        round_inst_srout2_z[58]) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n509), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n508), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U124 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n507), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n506), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n508) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U123 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n505), .A2(round_inst_n42), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n506) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n504), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n503), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n502), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n501), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n503) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U120 ( .A(round_inst_sin_w[9]), 
        .B(round_inst_sin_x[7]), .ZN(round_inst_S_2__sbox_inst_com_z_inst_n501) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U119 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n500), .B(round_inst_sin_y[7]), 
        .Z(round_inst_S_2__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U118 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n499), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n498), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n500) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U117 ( .A1(round_inst_n43), 
        .A2(round_inst_S_2__sbox_inst_com_z_inst_n497), .A3(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n498) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U116 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n495), .A2(round_inst_sin_x[8]), 
        .A3(round_inst_sin_w[11]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n499) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U115 ( .A(
        round_inst_S_2__sbox_inst_n5), .B(round_inst_n43), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n495) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U114 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_2__sbox_inst_n5), .A3(round_inst_sin_x[11]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n509) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n491), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n493) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U111 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n490), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n489), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n491) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n488), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n486), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n490) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U108 ( .A1(
        round_inst_sin_w[10]), .A2(round_inst_sin_x[11]), .A3(round_inst_n42), 
        .ZN(round_inst_S_2__sbox_inst_com_z_inst_n492) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U107 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n484), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U106 ( .A1(
        round_inst_sin_w[10]), .A2(round_inst_S_2__sbox_inst_com_z_inst_n497), 
        .ZN(round_inst_S_2__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n505), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n484) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n482), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n481), .Z(round_inst_srout2_z[56]) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n479), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n478), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n483), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U101 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n483) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U100 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n475), .A2(round_inst_sin_x[8]), 
        .A3(round_inst_sin_w[10]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U99 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n474), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n477) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U98 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n472), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .A3(round_inst_n43), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n473) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U97 ( .A(round_inst_sin_w[9]), 
        .B(round_inst_sin_y[9]), .Z(round_inst_S_2__sbox_inst_com_z_inst_n472)
         );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U96 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n471), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n474) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U95 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n469), .A2(
        round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n470) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n467), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n471) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n466), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n465), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n464), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n463), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U91 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n462), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n461), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U90 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n460), .A2(round_inst_n43), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n461) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U89 ( .A1(round_inst_n61), 
        .A2(round_inst_S_2__sbox_inst_n5), .A3(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n462) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n459), .A2(round_inst_n42), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U87 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_w[10]), 
        .ZN(round_inst_S_2__sbox_inst_com_z_inst_n466) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U85 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U84 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n453), .A2(round_inst_n43), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n454) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U83 ( .A(round_inst_sin_w[9]), 
        .B(round_inst_S_2__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n451), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U81 ( .A1(round_inst_sin_w[10]), .A2(round_inst_sin_x[8]), .ZN(round_inst_S_2__sbox_inst_com_z_inst_n478) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U79 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n487), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n448) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U78 ( .A(round_inst_sin_y[5]), 
        .B(round_inst_sin_x[5]), .Z(round_inst_S_2__sbox_inst_com_z_inst_n447)
         );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n487) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U76 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n446), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U75 ( .A(round_inst_sin_w[10]), 
        .B(round_inst_n43), .ZN(round_inst_S_2__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_srout2_z[59]) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n511), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U72 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n511) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U71 ( .A1(round_inst_sin_x[8]), 
        .A2(round_inst_sin_w[11]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n441) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U70 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n458), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n440), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n442) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U69 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U68 ( .A(round_inst_sin_w[11]), 
        .B(round_inst_S_2__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n497) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n494) );
  MUX2_X1 round_inst_S_2__sbox_inst_com_z_inst_U66 ( .A(round_inst_sin_x[11]), 
        .B(round_inst_sin_w[11]), .S(round_inst_S_2__sbox_inst_com_z_inst_n436), .Z(round_inst_S_2__sbox_inst_com_z_inst_n437) );
  OR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U65 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n436) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U64 ( .A(round_inst_sin_x[8]), 
        .B(round_inst_S_2__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n486) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U63 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n438) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U62 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_x[11]), 
        .A3(round_inst_S_2__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n430), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U59 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n429) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U58 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n426), .A2(round_inst_sin_w[11]), 
        .ZN(round_inst_S_2__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U56 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n422), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n424) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U55 ( .A1(round_inst_sin_x[8]), 
        .A2(round_inst_n61), .ZN(round_inst_S_2__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U54 ( .A1(round_inst_sin_y[9]), 
        .A2(round_inst_sin_x[8]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n425) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U53 ( .A1(round_inst_n42), 
        .A2(round_inst_sin_x[11]), .A3(round_inst_sin_w[9]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n428) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U52 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_y[11]), 
        .ZN(round_inst_S_2__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U50 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n460), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n423), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n469) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U49 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_y[9]), 
        .ZN(round_inst_S_2__sbox_inst_com_z_inst_n423) );
  AND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U48 ( .A1(round_inst_sin_w[9]), 
        .A2(round_inst_sin_x[8]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n460) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U47 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n421) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U46 ( .A1(round_inst_sin_w[9]), 
        .A2(round_inst_S_2__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .A2(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U44 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n419), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n418), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n432) );
  INV_X1 round_inst_S_2__sbox_inst_com_z_inst_U43 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .B(round_inst_n42), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n451) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U41 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n417), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n496), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U39 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n449) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U38 ( .A1(round_inst_sin_w[11]), .A2(round_inst_S_2__sbox_inst_com_z_inst_n413), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n414) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n415) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U35 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U34 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n505), .A2(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n409) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U32 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n407) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n405) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U30 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n404) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n505), .A2(round_inst_sin_y[9]), 
        .ZN(round_inst_S_2__sbox_inst_com_z_inst_n402) );
  AND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_S_2__sbox_inst_n5), .A2(round_inst_sin_w[11]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n505) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U27 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n401), .A2(round_inst_n43), .A3(
        round_inst_sin_w[9]), .ZN(round_inst_S_2__sbox_inst_com_z_inst_n403)
         );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U26 ( .A(round_inst_sin_w[11]), 
        .B(round_inst_sin_x[11]), .Z(round_inst_S_2__sbox_inst_com_z_inst_n401) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U25 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n399), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n406) );
  MUX2_X1 round_inst_S_2__sbox_inst_com_z_inst_U24 ( .A(round_inst_sin_y[11]), 
        .B(round_inst_S_2__sbox_inst_com_z_inst_n398), .S(
        round_inst_S_2__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U23 ( .A1(round_inst_sin_w[9]), 
        .A2(round_inst_S_2__sbox_inst_n5), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n398) );
  INV_X1 round_inst_S_2__sbox_inst_com_z_inst_U21 ( .A(round_inst_sin_x[11]), 
        .ZN(round_inst_S_2__sbox_inst_com_z_inst_n397) );
  NOR3_X1 round_inst_S_2__sbox_inst_com_z_inst_U20 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n488), .A3(
        round_inst_S_2__sbox_inst_com_z_inst_n395), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U19 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n394), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n395) );
  INV_X1 round_inst_S_2__sbox_inst_com_z_inst_U18 ( .A(round_inst_n61), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n394) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U17 ( .A(round_inst_sin_w[11]), 
        .B(round_inst_sin_y[11]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n488) );
  AND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U16 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n459), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U15 ( .A1(round_inst_sin_w[10]), .A2(round_inst_n61), .ZN(round_inst_S_2__sbox_inst_com_z_inst_n459) );
  INV_X1 round_inst_S_2__sbox_inst_com_z_inst_U14 ( .A(round_inst_sin_w[9]), 
        .ZN(round_inst_S_2__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U13 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n393), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U12 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n391), .A2(round_inst_n43), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U11 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_2__sbox_inst_com_z_inst_n390), .Z(
        round_inst_S_2__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U10 ( .A1(round_inst_sin_w[9]), 
        .A2(round_inst_sin_y[11]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n390) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U9 ( .A1(round_inst_n61), .A2(
        round_inst_sin_w[11]), .ZN(round_inst_S_2__sbox_inst_com_z_inst_n418)
         );
  NOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U8 ( .A1(
        round_inst_S_2__sbox_inst_com_z_inst_n439), .A2(
        round_inst_S_2__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_2__sbox_inst_com_z_inst_U7 ( .A1(round_inst_sin_w[10]), 
        .A2(round_inst_sin_w[9]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n456) );
  XNOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U6 ( .A(round_inst_sin_x[11]), 
        .B(round_inst_sin_y[11]), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n439) );
  NAND3_X1 round_inst_S_2__sbox_inst_com_z_inst_U5 ( .A1(round_inst_sin_w[10]), 
        .A2(round_inst_sin_x[11]), .A3(
        round_inst_S_2__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U4 ( .A(round_inst_n61), .B(
        round_inst_sin_y[9]), .Z(round_inst_S_2__sbox_inst_com_z_inst_n475) );
  INV_X1 round_inst_S_2__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_2__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_2__sbox_inst_com_z_inst_n496) );
  INV_X1 round_inst_S_2__sbox_inst_com_z_inst_U2 ( .A(round_inst_sin_w[8]), 
        .ZN(round_inst_S_2__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_2__sbox_inst_com_z_inst_U1 ( .A(round_inst_n41), .B(
        round_inst_sin_x[6]), .Z(round_inst_S_2__sbox_inst_com_z_inst_n417) );
  INV_X1 round_inst_S_3__sbox_inst_U6 ( .A(round_inst_sin_x[13]), .ZN(
        round_inst_S_3__sbox_inst_n4) );
  INV_X1 round_inst_S_3__sbox_inst_U5 ( .A(round_inst_sin_x[14]), .ZN(
        round_inst_S_3__sbox_inst_n6) );
  INV_X1 round_inst_S_3__sbox_inst_U4 ( .A(round_inst_sin_z[13]), .ZN(
        round_inst_S_3__sbox_inst_n2) );
  INV_X2 round_inst_S_3__sbox_inst_U3 ( .A(round_inst_S_3__sbox_inst_n4), .ZN(
        round_inst_S_3__sbox_inst_n3) );
  INV_X2 round_inst_S_3__sbox_inst_U2 ( .A(round_inst_S_3__sbox_inst_n6), .ZN(
        round_inst_S_3__sbox_inst_n5) );
  INV_X2 round_inst_S_3__sbox_inst_U1 ( .A(round_inst_S_3__sbox_inst_n2), .ZN(
        round_inst_S_3__sbox_inst_n1) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n531), .ZN(round_inst_sout_w[15])
         );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U139 ( .A1(
        round_inst_sin_z[12]), .A2(round_inst_S_3__sbox_inst_com_w_inst_n528), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n526), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n524), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n526) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[14]), .A2(round_inst_S_3__sbox_inst_com_w_inst_n523), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n525) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n518), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n516), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n518) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n514), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n513), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n512), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n513) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_w_inst_U128 ( .A1(
        round_inst_S_3__sbox_inst_n5), .A2(round_inst_sin_x[12]), .A3(
        round_inst_S_3__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n511) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U127 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n509), .A2(round_inst_sin_y[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n508), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n507), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U125 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n508) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_sin_z[15]), .A2(round_inst_S_3__sbox_inst_com_w_inst_n504), 
        .A3(round_inst_sin_x[12]), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U122 ( .A(round_inst_sin_y[11]), .B(round_inst_S_3__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U121 ( .A(
        round_inst_S_3__sbox_inst_n3), .B(round_inst_sin_z[11]), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n501) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U120 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[13])
         );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[9]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[9]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U113 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[12])
         );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_3__sbox_inst_n5), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U110 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n528), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U105 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_3__sbox_inst_n5), .B(round_inst_sin_z[14]), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_3__sbox_inst_n1), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U99 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n504), .A2(round_inst_sin_x[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_3__sbox_inst_n5), .A2(round_inst_sin_y[12]), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n507) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U94 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n461), .A2(
        round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U88 ( .A1(round_inst_sin_z[12]), 
        .A2(round_inst_S_3__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_w_inst_U85 ( .A1(round_inst_sin_y[13]), .A2(round_inst_sin_y[12]), .A3(round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_w_inst_U84 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_3__sbox_inst_n3), .A3(round_inst_sin_y[12]), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n528) );
  OR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_3__sbox_inst_n5), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U80 ( .A(round_inst_n42), .B(
        round_inst_sin_z[8]), .Z(round_inst_S_3__sbox_inst_com_w_inst_n484) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U79 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[15])
         );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U73 ( .A1(round_inst_sin_z[15]), .A2(round_inst_S_3__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U71 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_3__sbox_inst_n5), .A2(round_inst_sin_y[13]), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U69 ( .A1(
        round_inst_S_3__sbox_inst_n1), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_3__sbox_inst_n5), .A2(round_inst_S_3__sbox_inst_n1), .A3(
        round_inst_S_3__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n439), .A2(
        round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n505), .A2(
        round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U63 ( .A(round_inst_sin_z[15]), 
        .B(round_inst_S_3__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n505) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U62 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U61 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U60 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U58 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U57 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U56 ( .A(round_inst_sin_y[13]), 
        .B(round_inst_S_3__sbox_inst_n1), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U55 ( .A1(round_inst_sin_z[15]), .A2(round_inst_S_3__sbox_inst_n1), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U54 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_w_inst_U52 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n506), .A3(
        round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U51 ( .A(round_inst_sin_y[13]), 
        .B(round_inst_S_3__sbox_inst_n3), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_w_inst_U50 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n506), .A2(round_inst_sin_y[13]), 
        .A3(round_inst_S_3__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U49 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n504), .B(round_inst_sin_z[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n465) );
  INV_X1 round_inst_S_3__sbox_inst_com_w_inst_U48 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n436), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n504) );
  INV_X1 round_inst_S_3__sbox_inst_com_w_inst_U47 ( .A(round_inst_sin_y[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U45 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n520) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U44 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n421), .A2(round_inst_sin_z[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U43 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U42 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n419), .A2(
        round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U40 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_3__sbox_inst_n1), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U38 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n521) );
  INV_X1 round_inst_S_3__sbox_inst_com_w_inst_U37 ( .A(round_inst_sin_x[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n489) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U36 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U33 ( .A(round_inst_sin_x[12]), 
        .B(round_inst_sin_z[12]), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U32 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n498), .A2(
        round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U31 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U30 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U29 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U28 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U27 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U26 ( .A1(
        round_inst_S_3__sbox_inst_n3), .A2(round_inst_sin_z[12]), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n522), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U24 ( .A(
        round_inst_S_3__sbox_inst_n3), .B(round_inst_S_3__sbox_inst_n1), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_3__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U22 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U21 ( .A1(round_inst_sin_x[12]), .A2(round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U20 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[13]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U19 ( .A(round_inst_sin_y[12]), 
        .B(round_inst_sin_z[12]), .Z(round_inst_S_3__sbox_inst_com_w_inst_n418) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U17 ( .A(round_inst_sin_x[12]), 
        .B(round_inst_S_3__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U15 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n398), .A2(round_inst_sin_x[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U13 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n498), .B(
        round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_3__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_3__sbox_inst_com_w_inst_U11 ( .A(round_inst_sin_y[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_3__sbox_inst_n1), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U9 ( .A(round_inst_sin_z[15]), 
        .B(round_inst_S_3__sbox_inst_com_w_inst_n506), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n510) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U8 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U7 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_3__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_3__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U6 ( .A1(
        round_inst_S_3__sbox_inst_n3), .A2(round_inst_sin_y[12]), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U5 ( .A1(round_inst_sin_x[12]), 
        .A2(round_inst_sin_y[13]), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n477) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_w_inst_U4 ( .A1(
        round_inst_S_3__sbox_inst_com_w_inst_n506), .A2(round_inst_sin_y[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n522) );
  INV_X1 round_inst_S_3__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_3__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_3__sbox_inst_com_w_inst_n506) );
  INV_X1 round_inst_S_3__sbox_inst_com_w_inst_U2 ( .A(round_inst_sin_x[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_w_inst_n486) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_w_inst_U1 ( .A(round_inst_n43), .B(
        round_inst_sin_z[10]), .Z(round_inst_S_3__sbox_inst_com_w_inst_n402)
         );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U144 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n520), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n519), .Z(round_inst_sout_x[12])
         );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U143 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n518), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n517), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n519) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U142 ( .A(round_inst_sin_y[14]), .B(round_inst_sin_y[15]), .ZN(round_inst_S_3__sbox_inst_com_x_inst_n517) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U141 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n516), .B(round_inst_sin_z[8]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n518) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U140 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n515), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n514), .ZN(
        round_inst_srout2_x[14]) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U139 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n513), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n512), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n514) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U138 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n511), .A2(round_inst_sin_z[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n512) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U137 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n510), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n509), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n511) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U136 ( .A1(
        round_inst_sin_y[14]), .A2(round_inst_S_3__sbox_inst_com_x_inst_n508), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n507), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n506), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n513) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U133 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n510), .A2(round_inst_sin_w[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n504) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U132 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n503), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n502), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n501), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n500), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n502) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_x_inst_U130 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n499), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n498), .A3(round_inst_sin_y[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U129 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n496), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n501) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_x_inst_U128 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n495), .A2(round_inst_sin_y[12]), 
        .A3(round_inst_sin_y[14]), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U127 ( .A(round_inst_sin_y[15]), 
        .B(round_inst_sin_z[15]), .Z(round_inst_S_3__sbox_inst_com_x_inst_n495) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U126 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n494), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n410), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n497) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_x_inst_U125 ( .A1(
        round_inst_sin_y[14]), .A2(round_inst_sin_z[12]), .A3(
        round_inst_sin_z[15]), .ZN(round_inst_S_3__sbox_inst_com_x_inst_n503)
         );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U124 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n507) );
  OR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U123 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n494), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U122 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n489), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U121 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n488), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n487), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n489) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n486), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n485), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n487) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n484), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n485) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U118 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n508), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n483) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U117 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n481), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n484) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U116 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n478), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n480) );
  AND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U115 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n482), .A2(round_inst_sin_z[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n478) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U114 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .B(round_inst_sin_z[11]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n479) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_x_inst_U113 ( .A1(
        round_inst_sin_y[14]), .A2(round_inst_sin_w[12]), .A3(
        round_inst_sin_z[15]), .ZN(round_inst_S_3__sbox_inst_com_x_inst_n481)
         );
  NAND3_X1 round_inst_S_3__sbox_inst_com_x_inst_U112 ( .A1(
        round_inst_sin_y[14]), .A2(round_inst_sin_y[12]), .A3(
        round_inst_S_3__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n486) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U111 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n494), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n488) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_y[14]), .A2(round_inst_sin_z[12]), .A3(
        round_inst_sin_y[15]), .ZN(round_inst_S_3__sbox_inst_com_x_inst_n490)
         );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n520), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n475), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n515) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U108 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n474), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n473), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n520) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n472), .A2(round_inst_sin_y[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n473) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U106 ( .A(round_inst_sin_z[15]), .B(round_inst_S_3__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n472) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U105 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n470), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n510), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n474) );
  AND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U104 ( .A1(round_inst_sin_z[14]), .A2(round_inst_sin_y[15]), .ZN(round_inst_S_3__sbox_inst_com_x_inst_n510) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n468), .ZN(
        round_inst_srout2_x[12]) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n467), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n468) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U101 ( .A1(
        round_inst_sin_y[12]), .A2(round_inst_sin_z[14]), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U100 ( .A1(
        round_inst_sin_y[14]), .A2(round_inst_S_3__sbox_inst_com_x_inst_n499), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n467) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U99 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n469) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n464), .B(round_inst_sin_z[9]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n465) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n470), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n464) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U96 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n463), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n482) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U95 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n461), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n470) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U94 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n459), .A2(round_inst_sin_y[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n460) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n458), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n457), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n459) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_3__sbox_inst_n1), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n456), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n455), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n461) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U90 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n454), .A2(round_inst_sin_w[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n455) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n453), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n452), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n454) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U88 ( .A1(round_inst_sin_y[14]), .A2(round_inst_S_3__sbox_inst_n1), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n453) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n451), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n450), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n456) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U86 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n449), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n448), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U85 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n447), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n446), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n448) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n444), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n446) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n498), .B(round_inst_sin_z[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n444) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U82 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n443), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n445) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n442), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n441), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n449) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U80 ( .A1(round_inst_sin_y[14]), .A2(round_inst_sin_z[12]), .ZN(round_inst_S_3__sbox_inst_com_x_inst_n442) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_x_inst_U79 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n499), .A3(
        round_inst_S_3__sbox_inst_com_x_inst_n440), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n451) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U78 ( .A(round_inst_sin_z[14]), 
        .B(round_inst_S_3__sbox_inst_com_x_inst_n498), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n440) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U77 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n516), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_srout2_x[15]) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U76 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n438), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n439) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U75 ( .A(round_inst_sin_y[12]), 
        .B(round_inst_S_3__sbox_inst_com_x_inst_n475), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n437) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U74 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n436), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n435), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n475) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n434), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n433), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n435) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U72 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n432), .A2(round_inst_sin_w[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n433) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U71 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n431), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n430), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n432) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U70 ( .A1(
        round_inst_S_3__sbox_inst_n1), .A2(round_inst_sin_y[15]), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n430) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U69 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_z[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n431) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n429), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n428), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n434) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U67 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n427), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n428) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n425), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n424), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n426) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n423), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n422), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n424) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U64 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n508), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n457), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n422) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U63 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n441), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .B(round_inst_sin_w[13]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n441) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U61 ( .A1(round_inst_sin_z[15]), .A2(round_inst_S_3__sbox_inst_com_x_inst_n443), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n423) );
  AND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U60 ( .A1(round_inst_sin_y[12]), 
        .A2(round_inst_S_3__sbox_inst_com_x_inst_n421), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n443) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_x_inst_U59 ( .A1(round_inst_sin_w[13]), .A2(round_inst_S_3__sbox_inst_com_x_inst_n499), .A3(round_inst_sin_y[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U58 ( .A(round_inst_sin_z[12]), 
        .B(round_inst_sin_y[12]), .Z(round_inst_S_3__sbox_inst_com_x_inst_n499) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U57 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n420), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n419), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n427) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_3__sbox_inst_n1), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n417), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n416), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n418) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n417) );
  MUX2_X1 round_inst_S_3__sbox_inst_com_x_inst_U53 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n420), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n415), .S(
        round_inst_S_3__sbox_inst_com_x_inst_n414), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n436) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U52 ( .A1(round_inst_sin_y[15]), .A2(round_inst_S_3__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n414) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_y[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n413) );
  MUX2_X1 round_inst_S_3__sbox_inst_com_x_inst_U50 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n412), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n411), .S(
        round_inst_S_3__sbox_inst_com_x_inst_n410), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n415) );
  NOR3_X1 round_inst_S_3__sbox_inst_com_x_inst_U49 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n411), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n463), .A3(
        round_inst_S_3__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n412) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n420), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n411) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U47 ( .A(round_inst_sin_z[10]), 
        .B(round_inst_S_3__sbox_inst_com_x_inst_n466), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n407), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U45 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n406), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n407) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n405), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n406) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U43 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n419), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n405) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U42 ( .A(round_inst_sin_z[15]), 
        .B(round_inst_S_3__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n419) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U41 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n408) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_x_inst_U40 ( .A1(round_inst_sin_z[14]), .A2(round_inst_sin_y[15]), .A3(round_inst_S_3__sbox_inst_com_x_inst_n402), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n403) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U39 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n409), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n421), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n402) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U38 ( .A(
        round_inst_S_3__sbox_inst_n1), .B(round_inst_sin_w[13]), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n421) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U37 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n401), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n400), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n404) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U36 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n447), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n400) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U35 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n508), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n471) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n399), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n401) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U33 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n452), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U32 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n399) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U31 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n395), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n394), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n396) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U30 ( .A1(round_inst_sin_y[15]), .A2(round_inst_S_3__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n394) );
  MUX2_X1 round_inst_S_3__sbox_inst_com_x_inst_U29 ( .A(
        round_inst_S_3__sbox_inst_n1), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .S(
        round_inst_S_3__sbox_inst_com_x_inst_n498), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_3__sbox_inst_com_x_inst_U28 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n498) );
  INV_X1 round_inst_S_3__sbox_inst_com_x_inst_U27 ( .A(round_inst_sin_w[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n462) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n392), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n410), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n391), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n392) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U24 ( .A1(round_inst_sin_y[14]), .A2(round_inst_sin_w[13]), .ZN(round_inst_S_3__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U23 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_z[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n452) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U22 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n410), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n390), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n397) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U21 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n447), .Z(
        round_inst_S_3__sbox_inst_com_x_inst_n390) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U20 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n389), .A2(round_inst_sin_y[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n447) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_3__sbox_inst_n1), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n389) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n388), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n387), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n516) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U17 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n420), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n387) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U16 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_z[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n420) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U15 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n385), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n386) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U14 ( .A(round_inst_sin_w[13]), 
        .B(round_inst_S_3__sbox_inst_com_x_inst_n384), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n385) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_3__sbox_inst_n1), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n410), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n384) );
  INV_X1 round_inst_S_3__sbox_inst_com_x_inst_U12 ( .A(round_inst_sin_z[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n410) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n383), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n416), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n388) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_x_inst_U10 ( .A1(round_inst_sin_z[12]), .A2(round_inst_sin_y[15]), .ZN(round_inst_S_3__sbox_inst_com_x_inst_n416) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U9 ( .A1(
        round_inst_S_3__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_3__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_3__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_y[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U7 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n381), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n382) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_x_inst_U6 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_3__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_3__sbox_inst_com_x_inst_U5 ( .A(round_inst_sin_y[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n476) );
  INV_X1 round_inst_S_3__sbox_inst_com_x_inst_U4 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n477) );
  INV_X1 round_inst_S_3__sbox_inst_com_x_inst_U3 ( .A(round_inst_sin_y[13]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n409) );
  INV_X1 round_inst_S_3__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_3__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_3__sbox_inst_com_x_inst_n508) );
  INV_X1 round_inst_S_3__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_w[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_x_inst_n491) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n516), .Z(round_inst_sout_y[12])
         );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n515), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U134 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n513), .B(round_inst_sin_z[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n514) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U133 ( .A(round_inst_sin_x[8]), 
        .B(round_inst_S_3__sbox_inst_com_y_inst_n512), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n515) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n511), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_srout2_y[14]) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n507), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n517) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U129 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n506), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n505), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n507) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n505) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U127 ( .A1(
        round_inst_sin_w[14]), .A2(round_inst_sin_z[15]), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n506) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U125 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_3__sbox_inst_com_y_inst_U124 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_3__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U123 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_sin_x[15]), .A2(round_inst_S_3__sbox_inst_com_y_inst_n493), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U121 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n492), .A2(round_inst_sin_z[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U120 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U119 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U118 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U117 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n486), .A2(round_inst_sin_z[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U116 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_sin_w[14]), .A2(round_inst_sin_w[12]), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U114 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n513), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U112 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U111 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_3__sbox_inst_n1), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U109 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[11]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_y_inst_U108 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n513), .A2(round_inst_sin_z[15]), 
        .A3(round_inst_sin_x[12]), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U107 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_sin_w[12]), .A2(round_inst_sin_w[15]), .A3(
        round_inst_S_3__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_3__sbox_inst_com_y_inst_U105 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_3__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U104 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[12]) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U103 ( .A1(
        round_inst_S_3__sbox_inst_n5), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n508) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U98 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U97 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_3__sbox_inst_n1), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_3__sbox_inst_com_y_inst_U95 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U94 ( .A1(round_inst_sin_x[12]), .A2(round_inst_sin_w[14]), .ZN(round_inst_S_3__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_y_inst_U93 ( .A1(round_inst_sin_w[12]), .A2(round_inst_S_3__sbox_inst_n3), .A3(
        round_inst_S_3__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U92 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U91 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U88 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U87 ( .A1(
        round_inst_S_3__sbox_inst_n1), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_3__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_3__sbox_inst_n5), .B(round_inst_sin_w[14]), .S(
        round_inst_S_3__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U84 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U80 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_3__sbox_inst_n1), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U78 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n478), .B(round_inst_n61), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U77 ( .A1(round_inst_sin_w[14]), .A2(round_inst_S_3__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U76 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n513), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n438), .Z(round_inst_srout2_y[15]) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U71 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U70 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U69 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n483), .A2(
        round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_3__sbox_inst_n1), .A2(round_inst_sin_w[12]), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_y_inst_U66 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[15]), 
        .A3(round_inst_S_3__sbox_inst_n1), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U65 ( .A(round_inst_sin_w[12]), 
        .B(round_inst_sin_x[12]), .Z(round_inst_S_3__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U63 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U61 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U59 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U58 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U57 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[13]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U55 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_3__sbox_inst_com_y_inst_U54 ( .A(round_inst_sin_x[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U53 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n418), .A2(round_inst_sin_z[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U51 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U50 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U49 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n414), .B(
        round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U48 ( .A(round_inst_sin_w[13]), 
        .B(round_inst_S_3__sbox_inst_n1), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_3__sbox_inst_n1), .A2(round_inst_sin_x[12]), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U46 ( .A1(
        round_inst_S_3__sbox_inst_n1), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U45 ( .A(round_inst_sin_x[10]), 
        .B(round_inst_S_3__sbox_inst_com_y_inst_n512), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U44 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n512) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U43 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U42 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U41 ( .A(round_inst_sin_w[13]), 
        .B(round_inst_sin_x[15]), .Z(round_inst_S_3__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U40 ( .A(
        round_inst_S_3__sbox_inst_n3), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_3__sbox_inst_com_y_inst_U39 ( .A(round_inst_sin_w[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U38 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[12]), 
        .Z(round_inst_S_3__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_3__sbox_inst_com_y_inst_U36 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_3__sbox_inst_com_y_inst_U35 ( .A(round_inst_sin_z[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_3__sbox_inst_n1), .B(round_inst_sin_z[15]), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U30 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U29 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_3__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U27 ( .A(
        round_inst_S_3__sbox_inst_n5), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U26 ( .A1(round_inst_sin_w[13]), .A2(round_inst_sin_z[15]), .ZN(round_inst_S_3__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n513), .A2(round_inst_sin_w[13]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_3__sbox_inst_n1), .A2(round_inst_sin_w[15]), .A3(
        round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U22 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_3__sbox_inst_n1), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U21 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U20 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n397) );
  INV_X1 round_inst_S_3__sbox_inst_com_y_inst_U19 ( .A(round_inst_sin_w[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n396) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n503), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U17 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_z[15]), 
        .B(round_inst_sin_w[15]), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U15 ( .A(round_inst_sin_z[15]), 
        .B(round_inst_S_3__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n503) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U14 ( .A(round_inst_sin_w[15]), 
        .B(round_inst_sin_x[15]), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U13 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U12 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_y_inst_U11 ( .A1(
        round_inst_S_3__sbox_inst_n3), .A2(round_inst_sin_w[15]), .A3(
        round_inst_S_3__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_y_inst_U10 ( .A1(round_inst_sin_z[15]), .A2(round_inst_S_3__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_3__sbox_inst_com_y_inst_U9 ( .A(round_inst_sin_w[13]), 
        .B(round_inst_S_3__sbox_inst_n3), .S(round_inst_sin_w[14]), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_3__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_3__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_3__sbox_inst_n3), .A2(
        round_inst_S_3__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_3__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U6 ( .A(round_inst_sin_z[15]), 
        .B(round_inst_sin_x[15]), .Z(round_inst_S_3__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_y_inst_U5 ( .A1(
        round_inst_S_3__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_3__sbox_inst_n1), .A3(round_inst_sin_x[15]), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_3__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_y_inst_U3 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n513), .B(round_inst_sin_w[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_3__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_3__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_3__sbox_inst_com_y_inst_n513) );
  INV_X1 round_inst_S_3__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U137 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n523), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n522), .ZN(round_inst_sout_z[12])
         );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U136 ( .A(round_inst_sin_w[15]), .B(round_inst_S_3__sbox_inst_com_z_inst_n521), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n522) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U135 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n520), .B(round_inst_sin_w[14]), 
        .Z(round_inst_S_3__sbox_inst_com_z_inst_n523) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U134 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n519), .B(round_inst_sin_x[8]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n520) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U133 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n518), .B(round_inst_n42), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n519) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U132 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n517), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n516), .Z(round_inst_srout2_z[14]) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n515), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n514), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n516) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n512), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n514) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U129 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n511), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n510), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n512) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U128 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n509), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n508), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n518), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n507), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n511) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n506), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n505), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U125 ( .A(round_inst_sin_w[13]), .B(round_inst_sin_x[11]), .ZN(round_inst_S_3__sbox_inst_com_z_inst_n505) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U124 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n504), .B(round_inst_sin_y[11]), 
        .Z(round_inst_S_3__sbox_inst_com_z_inst_n506) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U123 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n503), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n502), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n504) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U122 ( .A1(
        round_inst_sin_y[12]), .A2(round_inst_S_3__sbox_inst_com_z_inst_n501), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n502) );
  INV_X1 round_inst_S_3__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n500), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n501) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U120 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n499), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n498), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n503) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_z_inst_U119 ( .A1(
        round_inst_sin_x[12]), .A2(round_inst_sin_w[15]), .A3(
        round_inst_S_3__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n498) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U118 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n496), .B(
        round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n497) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U117 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n495), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n494), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n499) );
  INV_X1 round_inst_S_3__sbox_inst_com_z_inst_U116 ( .A(round_inst_sin_x[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n494) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U115 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n500), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n518) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U114 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n491), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n493) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U113 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n508), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n490), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n491) );
  INV_X1 round_inst_S_3__sbox_inst_com_z_inst_U112 ( .A(round_inst_sin_w[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n490) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U111 ( .A1(
        round_inst_sin_w[14]), .A2(round_inst_S_3__sbox_inst_com_z_inst_n489), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n513) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U110 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n488), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n508), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n488) );
  INV_X1 round_inst_S_3__sbox_inst_com_z_inst_U108 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n486) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U107 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n484), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U106 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n482), .ZN(
        round_inst_srout2_z[12]) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n481), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n482) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U104 ( .A1(
        round_inst_sin_w[12]), .A2(round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n495) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n509), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n479), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n478), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n480) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U101 ( .A1(
        round_inst_sin_w[14]), .A2(round_inst_S_3__sbox_inst_com_z_inst_n485), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n478) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U100 ( .A(round_inst_sin_y[9]), 
        .B(round_inst_n61), .Z(round_inst_S_3__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U99 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n492), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n483) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U98 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n476), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n492) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U97 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n474), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n475) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U96 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n472), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n471), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U95 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n470), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n471) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U94 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n468), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n469) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n467), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n466), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n470) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n465), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n464), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n466) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U91 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n463), .A2(round_inst_sin_w[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n464) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U90 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n462), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U89 ( .A1(
        round_inst_S_3__sbox_inst_n3), .A2(round_inst_sin_y[12]), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n462) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U88 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n461), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n460), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U87 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n459), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n458), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n460) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n458) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U85 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n455), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n459) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U84 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n453), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n509), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U83 ( .A1(round_inst_sin_w[12]), .A2(round_inst_sin_y[14]), .ZN(round_inst_S_3__sbox_inst_com_z_inst_n509) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U82 ( .A1(round_inst_sin_w[14]), .A2(round_inst_sin_x[12]), .ZN(round_inst_S_3__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U81 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n452), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n461) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U80 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n450), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U79 ( .A(
        round_inst_S_3__sbox_inst_n5), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n449) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U78 ( .A(round_inst_sin_y[14]), 
        .B(round_inst_sin_w[14]), .Z(round_inst_S_3__sbox_inst_com_z_inst_n448) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n452), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U76 ( .A(round_inst_sin_w[14]), 
        .B(round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n452) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U75 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n446), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_srout2_z[15]) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n445) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U73 ( .A(round_inst_sin_w[12]), 
        .B(round_inst_S_3__sbox_inst_com_z_inst_n477), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U72 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n477) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U71 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n440), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n441) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U70 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n457), .A2(round_inst_sin_w[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n439) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U69 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n474), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n457) );
  AND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U68 ( .A1(round_inst_sin_w[13]), 
        .A2(round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n474) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n437), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n436), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U66 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n435), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n434), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n436) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U65 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n456), .A2(round_inst_sin_y[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n434) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U64 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n433), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n432), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n456) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U63 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n431), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n430), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U62 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n429), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n428), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n430) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_z_inst_U61 ( .A1(
        round_inst_S_3__sbox_inst_n3), .A2(round_inst_sin_w[15]), .A3(
        round_inst_S_3__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n428) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U60 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n427), .A2(round_inst_sin_w[13]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n429) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U59 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n426), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n425), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n427) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U58 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n424), .A2(
        round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U57 ( .A(round_inst_sin_x[15]), 
        .B(round_inst_sin_y[15]), .Z(round_inst_S_3__sbox_inst_com_z_inst_n424) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U56 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n422), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U55 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U54 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n419), .A2(round_inst_sin_w[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n420) );
  INV_X1 round_inst_S_3__sbox_inst_com_z_inst_U53 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n419) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U52 ( .A1(round_inst_sin_y[15]), .A2(round_inst_S_3__sbox_inst_com_z_inst_n438), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n421) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U51 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n418), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n500), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n423) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U50 ( .A1(round_inst_sin_w[15]), .A2(round_inst_S_3__sbox_inst_n5), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n500) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U49 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n417), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n432), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n437) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U48 ( .A1(round_inst_sin_w[13]), .A2(round_inst_sin_w[14]), .ZN(round_inst_S_3__sbox_inst_com_z_inst_n432) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U47 ( .A(round_inst_sin_x[15]), 
        .B(round_inst_sin_w[15]), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n417) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U46 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n416), .A2(round_inst_sin_x[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n442) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U45 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U44 ( .A(round_inst_sin_w[13]), 
        .B(round_inst_S_3__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n414) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U43 ( .A1(
        round_inst_S_3__sbox_inst_n3), .A2(round_inst_sin_w[14]), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n433) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n413), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n415) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U41 ( .A1(round_inst_sin_y[13]), .A2(round_inst_sin_w[14]), .ZN(round_inst_S_3__sbox_inst_com_z_inst_n413) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U40 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n412), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n438) );
  INV_X1 round_inst_S_3__sbox_inst_com_z_inst_U39 ( .A(round_inst_sin_y[14]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n496) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U38 ( .A(round_inst_n43), .B(
        round_inst_sin_x[10]), .Z(round_inst_S_3__sbox_inst_com_z_inst_n444)
         );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n521), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n517), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n411), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n410), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n517) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U35 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n409), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n408), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n410) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U34 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n407), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n406), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n408) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n405), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n406) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U32 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n403), .A2(round_inst_sin_y[15]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n404) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n402), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n401), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n405) );
  MUX2_X1 round_inst_S_3__sbox_inst_com_z_inst_U30 ( .A(round_inst_sin_x[15]), 
        .B(round_inst_sin_w[15]), .S(round_inst_S_3__sbox_inst_com_z_inst_n400), .Z(round_inst_S_3__sbox_inst_com_z_inst_n401) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U29 ( .A1(round_inst_sin_w[13]), .A2(round_inst_S_3__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n400) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U28 ( .A(round_inst_sin_w[12]), 
        .B(round_inst_sin_x[12]), .Z(round_inst_S_3__sbox_inst_com_z_inst_n485) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_z_inst_U27 ( .A1(round_inst_sin_w[15]), .A2(round_inst_S_3__sbox_inst_n3), .A3(
        round_inst_S_3__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n402) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U26 ( .A(round_inst_sin_w[12]), 
        .B(round_inst_sin_y[12]), .Z(round_inst_S_3__sbox_inst_com_z_inst_n473) );
  NAND3_X1 round_inst_S_3__sbox_inst_com_z_inst_U25 ( .A1(round_inst_sin_w[12]), .A2(round_inst_sin_x[15]), .A3(round_inst_S_3__sbox_inst_com_z_inst_n454), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n407) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U24 ( .A(
        round_inst_S_3__sbox_inst_n3), .B(round_inst_sin_y[13]), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n454) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U23 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n484), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n409) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U22 ( .A1(round_inst_sin_w[12]), .A2(round_inst_sin_y[13]), .ZN(round_inst_S_3__sbox_inst_com_z_inst_n447) );
  INV_X1 round_inst_S_3__sbox_inst_com_z_inst_U21 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n425), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n484) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U20 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n399), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n398), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n411) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U19 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n418), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n398) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U18 ( .A(round_inst_sin_y[13]), 
        .B(round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n418) );
  NOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U17 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_3__sbox_inst_com_z_inst_n412), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n399) );
  INV_X1 round_inst_S_3__sbox_inst_com_z_inst_U16 ( .A(round_inst_sin_w[13]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n412) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U15 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n395), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U14 ( .A1(round_inst_sin_x[15]), .A2(round_inst_sin_y[12]), .ZN(round_inst_S_3__sbox_inst_com_z_inst_n487) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U13 ( .A1(round_inst_sin_y[15]), .A2(round_inst_sin_x[12]), .ZN(round_inst_S_3__sbox_inst_com_z_inst_n395) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U12 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n394), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n393), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n521) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U11 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n392), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U10 ( .A1(round_inst_sin_x[12]), .A2(round_inst_sin_w[13]), .ZN(round_inst_S_3__sbox_inst_com_z_inst_n450) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U9 ( .A1(
        round_inst_S_3__sbox_inst_com_z_inst_n391), .A2(round_inst_sin_w[12]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n392) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U8 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n508), .B(round_inst_sin_y[13]), 
        .ZN(round_inst_S_3__sbox_inst_com_z_inst_n391) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U7 ( .A(round_inst_sin_x[15]), 
        .B(round_inst_S_3__sbox_inst_com_z_inst_n425), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n508) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U6 ( .A(round_inst_sin_w[15]), 
        .B(round_inst_sin_y[15]), .Z(round_inst_S_3__sbox_inst_com_z_inst_n425) );
  XNOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U5 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n394) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U4 ( .A1(round_inst_sin_w[15]), 
        .A2(round_inst_sin_x[12]), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n397) );
  XOR2_X1 round_inst_S_3__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_3__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_3__sbox_inst_com_z_inst_n451), .Z(
        round_inst_S_3__sbox_inst_com_z_inst_n403) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U2 ( .A1(round_inst_sin_w[12]), 
        .A2(round_inst_S_3__sbox_inst_n3), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n451) );
  NAND2_X1 round_inst_S_3__sbox_inst_com_z_inst_U1 ( .A1(round_inst_sin_w[12]), 
        .A2(round_inst_sin_w[13]), .ZN(
        round_inst_S_3__sbox_inst_com_z_inst_n468) );
  INV_X1 round_inst_S_4__sbox_inst_U6 ( .A(round_inst_sin_x[18]), .ZN(
        round_inst_S_4__sbox_inst_n6) );
  INV_X1 round_inst_S_4__sbox_inst_U5 ( .A(round_inst_sin_z[17]), .ZN(
        round_inst_S_4__sbox_inst_n2) );
  INV_X1 round_inst_S_4__sbox_inst_U4 ( .A(round_inst_sin_z[19]), .ZN(
        round_inst_S_4__sbox_inst_n4) );
  INV_X2 round_inst_S_4__sbox_inst_U3 ( .A(round_inst_S_4__sbox_inst_n2), .ZN(
        round_inst_S_4__sbox_inst_n1) );
  INV_X2 round_inst_S_4__sbox_inst_U2 ( .A(round_inst_S_4__sbox_inst_n4), .ZN(
        round_inst_S_4__sbox_inst_n3) );
  INV_X2 round_inst_S_4__sbox_inst_U1 ( .A(round_inst_S_4__sbox_inst_n6), .ZN(
        round_inst_S_4__sbox_inst_n5) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n531), .ZN(round_inst_sout_w[19])
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U139 ( .A1(
        round_inst_sin_z[16]), .A2(round_inst_S_4__sbox_inst_com_w_inst_n528), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n526), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n524), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n526) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[18]), .A2(round_inst_S_4__sbox_inst_com_w_inst_n523), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n525) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n518), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n516), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n518) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n514), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n513), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n512), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n513) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_w_inst_U128 ( .A1(
        round_inst_S_4__sbox_inst_n5), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n510), .A3(
        round_inst_S_4__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n511) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U127 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n508), .A2(round_inst_n44), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n507), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U125 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n507) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_4__sbox_inst_n3), .A2(round_inst_n45), .A3(
        round_inst_S_4__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U122 ( .A(round_inst_sin_y[15]), .B(round_inst_S_4__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U121 ( .A(round_inst_n62), .B(
        round_inst_sin_z[15]), .Z(round_inst_S_4__sbox_inst_com_w_inst_n501)
         );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U120 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[17])
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[13]), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[13]), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U113 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[16])
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_4__sbox_inst_n5), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U110 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n528), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U105 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_4__sbox_inst_n5), .B(round_inst_sin_z[18]), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_4__sbox_inst_n1), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U99 ( .A1(round_inst_n45), 
        .A2(round_inst_S_4__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_4__sbox_inst_n5), .A2(round_inst_n44), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n506) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U94 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[18]), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n461), .A2(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[18]), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U88 ( .A1(round_inst_sin_z[16]), 
        .A2(round_inst_S_4__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_w_inst_U85 ( .A1(round_inst_sin_y[17]), .A2(round_inst_n44), .A3(round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_w_inst_U84 ( .A1(round_inst_n45), 
        .A2(round_inst_n62), .A3(round_inst_n44), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n528) );
  OR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_4__sbox_inst_n5), .B(round_inst_n45), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U80 ( .A(round_inst_sin_y[12]), 
        .B(round_inst_sin_z[12]), .Z(round_inst_S_4__sbox_inst_com_w_inst_n484) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U79 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[19])
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U73 ( .A1(
        round_inst_S_4__sbox_inst_n3), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U71 ( .A1(round_inst_n45), 
        .A2(round_inst_n62), .ZN(round_inst_S_4__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_4__sbox_inst_n5), .A2(round_inst_sin_y[17]), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U69 ( .A1(
        round_inst_S_4__sbox_inst_n1), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n508), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_4__sbox_inst_n5), .A2(round_inst_S_4__sbox_inst_n1), .A3(
        round_inst_S_4__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n439), .A2(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n508), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_4__sbox_inst_n3), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n504) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U62 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n508) );
  INV_X1 round_inst_S_4__sbox_inst_com_w_inst_U61 ( .A(round_inst_n45), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U60 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U58 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U57 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U56 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U55 ( .A(round_inst_sin_y[17]), 
        .B(round_inst_S_4__sbox_inst_n1), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U54 ( .A1(
        round_inst_S_4__sbox_inst_n3), .A2(round_inst_S_4__sbox_inst_n1), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U52 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_w_inst_U51 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n505), .A3(
        round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U50 ( .A(round_inst_sin_y[17]), 
        .B(round_inst_n62), .Z(round_inst_S_4__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_w_inst_U49 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n505), .A2(round_inst_sin_y[17]), 
        .A3(round_inst_S_4__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U48 ( .A(round_inst_n45), .B(
        round_inst_sin_z[18]), .ZN(round_inst_S_4__sbox_inst_com_w_inst_n465)
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U47 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n520) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U45 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n421), .A2(
        round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U44 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U43 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n419), .A2(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U42 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U40 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_4__sbox_inst_n1), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n521) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U38 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U37 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U36 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n510), .B(round_inst_sin_z[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n498), .A2(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U33 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U32 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U31 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U30 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U29 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U28 ( .A1(round_inst_n62), 
        .A2(round_inst_sin_z[16]), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U27 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n522), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U26 ( .A(round_inst_n62), .B(
        round_inst_S_4__sbox_inst_n1), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U24 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n510), .A2(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U22 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[17]), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U21 ( .A(round_inst_n44), .B(
        round_inst_sin_z[16]), .Z(round_inst_S_4__sbox_inst_com_w_inst_n418)
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U20 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U19 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U17 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n398), .A2(
        round_inst_S_4__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U15 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n498), .B(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_4__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_4__sbox_inst_com_w_inst_U13 ( .A(round_inst_sin_y[19]), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_4__sbox_inst_n1), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U11 ( .A(
        round_inst_S_4__sbox_inst_n3), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n505), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U9 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_4__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_4__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U8 ( .A1(round_inst_n62), .A2(
        round_inst_n44), .ZN(round_inst_S_4__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U7 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n510), .A2(round_inst_sin_y[17]), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n477) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_w_inst_U6 ( .A1(
        round_inst_S_4__sbox_inst_com_w_inst_n505), .A2(round_inst_n44), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n522) );
  INV_X1 round_inst_S_4__sbox_inst_com_w_inst_U5 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n505) );
  INV_X1 round_inst_S_4__sbox_inst_com_w_inst_U4 ( .A(round_inst_sin_x[19]), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n486) );
  INV_X1 round_inst_S_4__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_4__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_4__sbox_inst_com_w_inst_n510) );
  INV_X1 round_inst_S_4__sbox_inst_com_w_inst_U2 ( .A(round_inst_sin_x[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_w_inst_n489) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_w_inst_U1 ( .A(round_inst_sin_y[14]), 
        .B(round_inst_sin_z[14]), .Z(round_inst_S_4__sbox_inst_com_w_inst_n402) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n510), .ZN(round_inst_sout_x[16])
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n509), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n510) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U133 ( .A(round_inst_n45), .B(
        round_inst_sin_y[19]), .ZN(round_inst_S_4__sbox_inst_com_x_inst_n508)
         );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U132 ( .A(round_inst_sin_z[12]), 
        .B(round_inst_S_4__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n506), .Z(round_inst_srout2_x[34]) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U130 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U129 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n503), .A2(round_inst_sin_z[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U127 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U126 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U125 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U124 ( .A1(round_inst_n45), 
        .A2(round_inst_sin_w[16]), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U122 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U121 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U118 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_sin_y[19]), .A2(round_inst_S_4__sbox_inst_com_x_inst_n490), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U115 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n487) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_x_inst_U114 ( .A1(
        round_inst_sin_z[18]), .A2(round_inst_sin_w[16]), .A3(
        round_inst_sin_y[19]), .ZN(round_inst_S_4__sbox_inst_com_x_inst_n489)
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n478), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n476), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n478) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n475), .B(round_inst_sin_z[15]), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n476) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_w[18]), .A2(round_inst_sin_y[19]), .A3(
        round_inst_sin_z[16]), .ZN(round_inst_S_4__sbox_inst_com_x_inst_n475)
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n474), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n473), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n473) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n470), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n469), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n511) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n468), .A2(round_inst_n45), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n469) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n468) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n467), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n464), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_srout2_x[32]) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U100 ( .A1(round_inst_n44), 
        .A2(round_inst_sin_z[18]), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[13]), 
        .B(round_inst_S_4__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n464) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n462), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n460), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n467), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n461) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n458), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n467) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_4__sbox_inst_n1), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n457), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n459) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n455), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n454), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n456) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n453), .A2(round_inst_sin_w[18]), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n454) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n451), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n455) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n450), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n449), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n451) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n448), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n447), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n449) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n446), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_4__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n445), .B(round_inst_n45), .S(
        round_inst_n44), .Z(round_inst_S_4__sbox_inst_com_x_inst_n446) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n444), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n448) );
  MUX2_X1 round_inst_S_4__sbox_inst_com_x_inst_U85 ( .A(round_inst_n45), .B(
        round_inst_sin_z[18]), .S(round_inst_sin_z[16]), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n443), .A2(round_inst_sin_w[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n442), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n441), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n452) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[16]), 
        .A3(round_inst_sin_z[18]), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n441) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n440), .A2(round_inst_sin_w[17]), 
        .A3(round_inst_n45), .ZN(round_inst_S_4__sbox_inst_com_x_inst_n442) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U80 ( .A(round_inst_n44), .B(
        round_inst_sin_z[16]), .Z(round_inst_S_4__sbox_inst_com_x_inst_n440)
         );
  NAND3_X1 round_inst_S_4__sbox_inst_com_x_inst_U79 ( .A1(round_inst_n44), 
        .A2(round_inst_S_4__sbox_inst_com_x_inst_n445), .A3(
        round_inst_S_4__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n460) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U77 ( .A1(round_inst_n44), 
        .A2(round_inst_n45), .ZN(round_inst_S_4__sbox_inst_com_x_inst_n482) );
  AND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U76 ( .A1(round_inst_n45), .A2(
        round_inst_sin_z[16]), .ZN(round_inst_S_4__sbox_inst_com_x_inst_n490)
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n462) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U74 ( .A1(round_inst_n44), 
        .A2(round_inst_sin_w[18]), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n497) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_srout2_x[35]) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n436), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n435), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U71 ( .A(round_inst_n44), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n435) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n434), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n433), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U69 ( .A1(round_inst_sin_z[16]), .A2(round_inst_sin_y[19]), .ZN(round_inst_S_4__sbox_inst_com_x_inst_n433) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n432), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n431), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n434) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n430), .A2(round_inst_n44), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n431) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n429), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n428), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_4__sbox_inst_n1), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n453), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n432) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[14]), 
        .B(round_inst_S_4__sbox_inst_com_x_inst_n438), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n436) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n425), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n424), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n423), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n422), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n421), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n420), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n422) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n419), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n420) );
  NOR3_X1 round_inst_S_4__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n471), .A3(
        round_inst_S_4__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n418) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n416), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n419) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n414), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U53 ( .A1(round_inst_n45), 
        .A2(round_inst_S_4__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n413) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U52 ( .A(round_inst_sin_y[19]), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n414) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n443), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n416) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U50 ( .A1(
        round_inst_S_4__sbox_inst_n1), .A2(round_inst_n45), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n443) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_x_inst_U49 ( .A1(round_inst_n45), 
        .A2(round_inst_S_4__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_4__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n421) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n411), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n423) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U47 ( .A1(round_inst_n45), 
        .A2(round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n465) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n411) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n410), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n407), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U43 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n406), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n405), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n407) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U42 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n466), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n405) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U41 ( .A(round_inst_sin_w[17]), 
        .B(round_inst_S_4__sbox_inst_n1), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n439) );
  AND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U40 ( .A1(round_inst_sin_z[18]), 
        .A2(round_inst_sin_y[19]), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_4__sbox_inst_n3), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n406) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_x_inst_U38 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U37 ( .A(round_inst_sin_z[18]), 
        .B(round_inst_sin_w[18]), .Z(round_inst_S_4__sbox_inst_com_x_inst_n445) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U36 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n404), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n410) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U35 ( .A(round_inst_sin_w[18]), 
        .B(round_inst_n45), .Z(round_inst_S_4__sbox_inst_com_x_inst_n403) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n402), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n401), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U33 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n400), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n399), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n401) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U32 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n399) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U31 ( .A1(round_inst_sin_z[16]), .A2(round_inst_S_4__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n426) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n427), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n400) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U28 ( .A(round_inst_sin_y[19]), 
        .B(round_inst_S_4__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n471) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n402) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_4__sbox_inst_n1), .A3(round_inst_n44), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n396) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n398), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n481) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U23 ( .A(round_inst_sin_y[19]), 
        .B(round_inst_S_4__sbox_inst_n3), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U21 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n392), .A2(round_inst_sin_w[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n404), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_x_inst_U17 ( .A1(round_inst_sin_z[16]), .A2(round_inst_sin_y[19]), .A3(round_inst_sin_w[17]), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n388) );
  MUX2_X1 round_inst_S_4__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n412), .B(round_inst_sin_y[19]), 
        .S(round_inst_S_4__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U15 ( .A1(round_inst_n44), 
        .A2(round_inst_S_4__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U14 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n491), .B(
        round_inst_S_4__sbox_inst_n3), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n412) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n384), .A2(round_inst_sin_z[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U10 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_4__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U9 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_w[19]), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U7 ( .A1(
        round_inst_S_4__sbox_inst_n1), .A2(round_inst_sin_y[19]), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n404) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_4__sbox_inst_com_x_inst_n427), .Z(
        round_inst_S_4__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U4 ( .A1(round_inst_n44), .A2(
        round_inst_sin_w[17]), .ZN(round_inst_S_4__sbox_inst_com_x_inst_n427)
         );
  NAND2_X1 round_inst_S_4__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_4__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_4__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_4__sbox_inst_com_x_inst_n477) );
  INV_X1 round_inst_S_4__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_y[17]), 
        .ZN(round_inst_S_4__sbox_inst_com_x_inst_n417) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n517), .Z(round_inst_sout_y[16])
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n516), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n515) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U134 ( .A(round_inst_sin_x[12]), 
        .B(round_inst_S_4__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n512), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_srout2_y[34]) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n508), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n518) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n507), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n506), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n508) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n506) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n507) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_4__sbox_inst_com_y_inst_U125 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_4__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U124 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U123 ( .A1(
        round_inst_sin_x[19]), .A2(round_inst_S_4__sbox_inst_com_y_inst_n493), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n492), .A2(
        round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U121 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U120 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U119 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U118 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n486), .A2(
        round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U117 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n503), .A2(round_inst_sin_w[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U112 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_4__sbox_inst_n1), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[15]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_y_inst_U109 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_4__sbox_inst_n3), .A3(round_inst_sin_x[16]), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U108 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_y_inst_U107 ( .A1(
        round_inst_sin_w[16]), .A2(round_inst_sin_w[19]), .A3(
        round_inst_S_4__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_4__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_4__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U105 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[32]) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U104 ( .A1(
        round_inst_S_4__sbox_inst_n5), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U98 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_4__sbox_inst_n1), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U95 ( .A1(round_inst_sin_x[16]), .A2(round_inst_S_4__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_y_inst_U94 ( .A1(round_inst_sin_w[16]), .A2(round_inst_n62), .A3(round_inst_S_4__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U93 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U92 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U88 ( .A1(
        round_inst_S_4__sbox_inst_n1), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_4__sbox_inst_com_y_inst_U87 ( .A(
        round_inst_S_4__sbox_inst_n5), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n503), .S(
        round_inst_S_4__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_4__sbox_inst_n1), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n478), .B(round_inst_sin_x[13]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n438), .Z(round_inst_srout2_y[35]) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U71 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[19]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U70 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n483), .A2(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_4__sbox_inst_n1), .A2(round_inst_sin_w[16]), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[19]), 
        .A3(round_inst_S_4__sbox_inst_n1), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U66 ( .A(round_inst_sin_w[16]), 
        .B(round_inst_sin_x[16]), .Z(round_inst_S_4__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U59 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[19]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U58 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[17]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U55 ( .A(round_inst_sin_x[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U54 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n418), .A2(
        round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U53 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U51 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U50 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n414), .B(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U49 ( .A(round_inst_sin_w[17]), 
        .B(round_inst_S_4__sbox_inst_n1), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U48 ( .A1(
        round_inst_S_4__sbox_inst_n1), .A2(round_inst_sin_x[16]), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_4__sbox_inst_n1), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U46 ( .A(round_inst_sin_x[14]), 
        .B(round_inst_S_4__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n513) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[17]), 
        .B(round_inst_sin_x[19]), .Z(round_inst_S_4__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U41 ( .A(round_inst_n62), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[19]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[16]), 
        .Z(round_inst_S_4__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U36 ( .A(round_inst_sin_z[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_4__sbox_inst_n1), .B(round_inst_S_4__sbox_inst_n3), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_4__sbox_inst_n5), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U27 ( .A1(round_inst_sin_w[17]), .A2(round_inst_S_4__sbox_inst_n3), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n514), .A2(round_inst_sin_w[17]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_4__sbox_inst_n1), .A2(round_inst_sin_w[19]), .A3(
        round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_4__sbox_inst_n1), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n504), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_4__sbox_inst_n3), .B(round_inst_sin_w[19]), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U17 ( .A(
        round_inst_S_4__sbox_inst_n3), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[19]), 
        .B(round_inst_sin_x[19]), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_y_inst_U13 ( .A1(round_inst_n62), 
        .A2(round_inst_sin_w[19]), .A3(
        round_inst_S_4__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_y_inst_U12 ( .A1(
        round_inst_S_4__sbox_inst_n3), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_4__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[17]), 
        .B(round_inst_n62), .S(round_inst_S_4__sbox_inst_com_y_inst_n503), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_y_inst_U9 ( .A1(round_inst_n62), .A2(
        round_inst_S_4__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_4__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_4__sbox_inst_n3), .B(round_inst_sin_x[19]), .Z(
        round_inst_S_4__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_4__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_4__sbox_inst_n1), .A3(round_inst_sin_x[19]), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_4__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n503) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[18]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_4__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_4__sbox_inst_com_y_inst_n514) );
  INV_X1 round_inst_S_4__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[18]), 
        .ZN(round_inst_S_4__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n516), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n515), .ZN(round_inst_sout_z[16])
         );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n514), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n513), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_w[18]), .B(round_inst_sin_w[19]), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n513) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U128 ( .A(round_inst_sin_x[12]), 
        .B(round_inst_sin_y[12]), .Z(round_inst_S_4__sbox_inst_com_z_inst_n514) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n510), .ZN(
        round_inst_srout2_z[34]) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n509), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n508), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U124 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n507), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n506), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n508) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U123 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n505), .A2(round_inst_n44), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n506) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n504), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n503), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n502), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n501), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n503) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U120 ( .A(round_inst_sin_w[17]), .B(round_inst_sin_x[15]), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n501) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U119 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n500), .B(round_inst_sin_y[15]), 
        .Z(round_inst_S_4__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U118 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n499), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n498), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n500) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U117 ( .A1(round_inst_n45), 
        .A2(round_inst_S_4__sbox_inst_com_z_inst_n497), .A3(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n498) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U116 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n495), .A2(round_inst_sin_x[16]), 
        .A3(round_inst_sin_w[19]), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n499) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U115 ( .A(
        round_inst_S_4__sbox_inst_n5), .B(round_inst_n45), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n495) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U114 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_4__sbox_inst_n5), .A3(round_inst_sin_x[19]), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n509) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n491), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n493) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U111 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n490), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n489), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n491) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n488), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n486), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n490) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U108 ( .A1(
        round_inst_sin_w[18]), .A2(round_inst_sin_x[19]), .A3(round_inst_n44), 
        .ZN(round_inst_S_4__sbox_inst_com_z_inst_n492) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U107 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n484), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U106 ( .A1(
        round_inst_sin_w[18]), .A2(round_inst_S_4__sbox_inst_com_z_inst_n497), 
        .ZN(round_inst_S_4__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n505), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n484) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n482), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n481), .Z(round_inst_srout2_z[32]) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n479), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n478), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n483), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U101 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n483) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U100 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n475), .A2(round_inst_sin_x[16]), 
        .A3(round_inst_sin_w[18]), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U99 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n474), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n477) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U98 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n472), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .A3(round_inst_n45), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n473) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U97 ( .A(round_inst_sin_w[17]), 
        .B(round_inst_sin_y[17]), .Z(round_inst_S_4__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U96 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n471), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n474) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U95 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n469), .A2(
        round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n470) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n467), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n471) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n466), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n465), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n464), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n463), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U91 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n462), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n461), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U90 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n460), .A2(round_inst_n45), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n461) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U89 ( .A1(round_inst_n62), 
        .A2(round_inst_S_4__sbox_inst_n5), .A3(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n462) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n459), .A2(round_inst_n44), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U87 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_w[18]), 
        .ZN(round_inst_S_4__sbox_inst_com_z_inst_n466) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U85 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U84 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n453), .A2(round_inst_n45), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n454) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U83 ( .A(round_inst_sin_w[17]), 
        .B(round_inst_S_4__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n451), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U81 ( .A1(round_inst_sin_w[18]), .A2(round_inst_sin_x[16]), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n478) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U79 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n487), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n448) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U78 ( .A(round_inst_sin_y[13]), 
        .B(round_inst_sin_x[13]), .Z(round_inst_S_4__sbox_inst_com_z_inst_n447) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n487) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U76 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n446), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U75 ( .A(round_inst_sin_w[18]), 
        .B(round_inst_n45), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_srout2_z[35]) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n511), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U72 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n511) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U71 ( .A1(round_inst_sin_x[16]), .A2(round_inst_sin_w[19]), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n441) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U70 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n458), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n440), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n442) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U69 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U68 ( .A(round_inst_sin_w[19]), 
        .B(round_inst_S_4__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n497) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n494) );
  MUX2_X1 round_inst_S_4__sbox_inst_com_z_inst_U66 ( .A(round_inst_sin_x[19]), 
        .B(round_inst_sin_w[19]), .S(round_inst_S_4__sbox_inst_com_z_inst_n436), .Z(round_inst_S_4__sbox_inst_com_z_inst_n437) );
  OR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U65 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n436) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U64 ( .A(round_inst_sin_x[16]), 
        .B(round_inst_S_4__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n486) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U63 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n438) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U62 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_x[19]), 
        .A3(round_inst_S_4__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n430), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U59 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n429) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U58 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n426), .A2(round_inst_sin_w[19]), 
        .ZN(round_inst_S_4__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U56 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n422), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n424) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U55 ( .A1(round_inst_sin_x[16]), .A2(round_inst_n62), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U54 ( .A1(round_inst_sin_y[17]), .A2(round_inst_sin_x[16]), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n425) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U53 ( .A1(round_inst_n44), 
        .A2(round_inst_sin_x[19]), .A3(round_inst_sin_w[17]), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n428) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U52 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_y[19]), 
        .ZN(round_inst_S_4__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U50 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n460), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n423), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n469) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U49 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_y[17]), 
        .ZN(round_inst_S_4__sbox_inst_com_z_inst_n423) );
  AND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U48 ( .A1(round_inst_sin_w[17]), 
        .A2(round_inst_sin_x[16]), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n460) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U47 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n421) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U46 ( .A1(round_inst_sin_w[17]), .A2(round_inst_S_4__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .A2(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U44 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n419), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n418), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n432) );
  INV_X1 round_inst_S_4__sbox_inst_com_z_inst_U43 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .B(round_inst_n44), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n451) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U41 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n417), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n496), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U39 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n449) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U38 ( .A1(round_inst_sin_w[19]), .A2(round_inst_S_4__sbox_inst_com_z_inst_n413), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n414) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n415) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U35 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U34 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n505), .A2(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n409) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U32 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n407) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n405) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U30 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n404) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n505), .A2(round_inst_sin_y[17]), 
        .ZN(round_inst_S_4__sbox_inst_com_z_inst_n402) );
  AND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_S_4__sbox_inst_n5), .A2(round_inst_sin_w[19]), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n505) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U27 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n401), .A2(round_inst_n45), .A3(
        round_inst_sin_w[17]), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n403)
         );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U26 ( .A(round_inst_sin_w[19]), 
        .B(round_inst_sin_x[19]), .Z(round_inst_S_4__sbox_inst_com_z_inst_n401) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U25 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n399), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n406) );
  MUX2_X1 round_inst_S_4__sbox_inst_com_z_inst_U24 ( .A(round_inst_sin_y[19]), 
        .B(round_inst_S_4__sbox_inst_com_z_inst_n398), .S(
        round_inst_S_4__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U23 ( .A1(round_inst_sin_w[17]), .A2(round_inst_S_4__sbox_inst_n5), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n398) );
  INV_X1 round_inst_S_4__sbox_inst_com_z_inst_U21 ( .A(round_inst_sin_x[19]), 
        .ZN(round_inst_S_4__sbox_inst_com_z_inst_n397) );
  NOR3_X1 round_inst_S_4__sbox_inst_com_z_inst_U20 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n488), .A3(
        round_inst_S_4__sbox_inst_com_z_inst_n395), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U19 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n394), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n395) );
  INV_X1 round_inst_S_4__sbox_inst_com_z_inst_U18 ( .A(round_inst_n62), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n394) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U17 ( .A(round_inst_sin_w[19]), 
        .B(round_inst_sin_y[19]), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n488) );
  AND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U16 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n459), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U15 ( .A1(round_inst_sin_w[18]), .A2(round_inst_n62), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n459) );
  INV_X1 round_inst_S_4__sbox_inst_com_z_inst_U14 ( .A(round_inst_sin_w[17]), 
        .ZN(round_inst_S_4__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U13 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n393), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U12 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n391), .A2(round_inst_n45), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U11 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_4__sbox_inst_com_z_inst_n390), .Z(
        round_inst_S_4__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U10 ( .A1(round_inst_sin_w[17]), .A2(round_inst_sin_y[19]), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n390) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U9 ( .A1(round_inst_n62), .A2(
        round_inst_sin_w[19]), .ZN(round_inst_S_4__sbox_inst_com_z_inst_n418)
         );
  NOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U8 ( .A1(
        round_inst_S_4__sbox_inst_com_z_inst_n439), .A2(
        round_inst_S_4__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_4__sbox_inst_com_z_inst_U7 ( .A1(round_inst_sin_w[18]), 
        .A2(round_inst_sin_w[17]), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n456) );
  XNOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U6 ( .A(round_inst_sin_x[19]), 
        .B(round_inst_sin_y[19]), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n439) );
  NAND3_X1 round_inst_S_4__sbox_inst_com_z_inst_U5 ( .A1(round_inst_sin_w[18]), 
        .A2(round_inst_sin_x[19]), .A3(
        round_inst_S_4__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U4 ( .A(round_inst_n62), .B(
        round_inst_sin_y[17]), .Z(round_inst_S_4__sbox_inst_com_z_inst_n475)
         );
  INV_X1 round_inst_S_4__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_4__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_4__sbox_inst_com_z_inst_n496) );
  INV_X1 round_inst_S_4__sbox_inst_com_z_inst_U2 ( .A(round_inst_sin_w[16]), 
        .ZN(round_inst_S_4__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_4__sbox_inst_com_z_inst_U1 ( .A(round_inst_sin_y[14]), 
        .B(round_inst_sin_x[14]), .Z(round_inst_S_4__sbox_inst_com_z_inst_n417) );
  INV_X1 round_inst_S_5__sbox_inst_U6 ( .A(round_inst_sin_x[22]), .ZN(
        round_inst_S_5__sbox_inst_n6) );
  INV_X1 round_inst_S_5__sbox_inst_U5 ( .A(round_inst_sin_z[21]), .ZN(
        round_inst_S_5__sbox_inst_n2) );
  INV_X1 round_inst_S_5__sbox_inst_U4 ( .A(round_inst_sin_z[23]), .ZN(
        round_inst_S_5__sbox_inst_n4) );
  INV_X2 round_inst_S_5__sbox_inst_U3 ( .A(round_inst_S_5__sbox_inst_n4), .ZN(
        round_inst_S_5__sbox_inst_n3) );
  INV_X2 round_inst_S_5__sbox_inst_U2 ( .A(round_inst_S_5__sbox_inst_n2), .ZN(
        round_inst_S_5__sbox_inst_n1) );
  INV_X2 round_inst_S_5__sbox_inst_U1 ( .A(round_inst_S_5__sbox_inst_n6), .ZN(
        round_inst_S_5__sbox_inst_n5) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n531), .ZN(round_inst_sout_w[23])
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U139 ( .A1(
        round_inst_sin_z[20]), .A2(round_inst_S_5__sbox_inst_com_w_inst_n528), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n526), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n524), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n526) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[22]), .A2(round_inst_S_5__sbox_inst_com_w_inst_n523), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n525) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n518), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n516), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n518) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n514), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n513), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n512), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n513) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_w_inst_U128 ( .A1(
        round_inst_S_5__sbox_inst_n5), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n510), .A3(
        round_inst_S_5__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n511) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U127 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n508), .A2(round_inst_n46), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n507), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U125 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n507) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_5__sbox_inst_n3), .A2(round_inst_n47), .A3(
        round_inst_S_5__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U122 ( .A(round_inst_sin_y[19]), .B(round_inst_S_5__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U121 ( .A(round_inst_n63), .B(
        round_inst_sin_z[19]), .Z(round_inst_S_5__sbox_inst_com_w_inst_n501)
         );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U120 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[21])
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[17]), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[17]), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U113 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[20])
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_5__sbox_inst_n5), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U110 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n528), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U105 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_5__sbox_inst_n5), .B(round_inst_sin_z[22]), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_5__sbox_inst_n1), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U99 ( .A1(round_inst_n47), 
        .A2(round_inst_S_5__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_5__sbox_inst_n5), .A2(round_inst_n46), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n506) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U94 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[22]), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n461), .A2(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[22]), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U88 ( .A1(round_inst_sin_z[20]), 
        .A2(round_inst_S_5__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_w_inst_U85 ( .A1(round_inst_sin_y[21]), .A2(round_inst_n46), .A3(round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_w_inst_U84 ( .A1(round_inst_n47), 
        .A2(round_inst_n63), .A3(round_inst_n46), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n528) );
  OR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_5__sbox_inst_n5), .B(round_inst_n47), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U80 ( .A(round_inst_n44), .B(
        round_inst_sin_z[16]), .Z(round_inst_S_5__sbox_inst_com_w_inst_n484)
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U79 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[23])
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U73 ( .A1(
        round_inst_S_5__sbox_inst_n3), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U71 ( .A1(round_inst_n47), 
        .A2(round_inst_n63), .ZN(round_inst_S_5__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_5__sbox_inst_n5), .A2(round_inst_sin_y[21]), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U69 ( .A1(
        round_inst_S_5__sbox_inst_n1), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n508), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_5__sbox_inst_n5), .A2(round_inst_S_5__sbox_inst_n1), .A3(
        round_inst_S_5__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n439), .A2(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n508), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_5__sbox_inst_n3), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n504) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U62 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n508) );
  INV_X1 round_inst_S_5__sbox_inst_com_w_inst_U61 ( .A(round_inst_n47), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U60 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U58 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U57 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U56 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U55 ( .A(round_inst_sin_y[21]), 
        .B(round_inst_S_5__sbox_inst_n1), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U54 ( .A1(
        round_inst_S_5__sbox_inst_n3), .A2(round_inst_S_5__sbox_inst_n1), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U52 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_w_inst_U51 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n505), .A3(
        round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U50 ( .A(round_inst_sin_y[21]), 
        .B(round_inst_n63), .Z(round_inst_S_5__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_w_inst_U49 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n505), .A2(round_inst_sin_y[21]), 
        .A3(round_inst_S_5__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U48 ( .A(round_inst_n47), .B(
        round_inst_sin_z[22]), .ZN(round_inst_S_5__sbox_inst_com_w_inst_n465)
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U47 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n520) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U45 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n421), .A2(
        round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U44 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U43 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n419), .A2(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U42 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U40 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_5__sbox_inst_n1), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n521) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U38 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U37 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U36 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n510), .B(round_inst_sin_z[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n498), .A2(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U33 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U32 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U31 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U30 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U29 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U28 ( .A1(round_inst_n63), 
        .A2(round_inst_sin_z[20]), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U27 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n522), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U26 ( .A(round_inst_n63), .B(
        round_inst_S_5__sbox_inst_n1), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U24 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n510), .A2(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U22 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[21]), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U21 ( .A(round_inst_n46), .B(
        round_inst_sin_z[20]), .Z(round_inst_S_5__sbox_inst_com_w_inst_n418)
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U20 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U19 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U17 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n398), .A2(
        round_inst_S_5__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U15 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n498), .B(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_5__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_5__sbox_inst_com_w_inst_U13 ( .A(round_inst_sin_y[23]), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_5__sbox_inst_n1), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U11 ( .A(
        round_inst_S_5__sbox_inst_n3), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n505), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U9 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_5__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_5__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U8 ( .A1(round_inst_n63), .A2(
        round_inst_n46), .ZN(round_inst_S_5__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U7 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n510), .A2(round_inst_sin_y[21]), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n477) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_w_inst_U6 ( .A1(
        round_inst_S_5__sbox_inst_com_w_inst_n505), .A2(round_inst_n46), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n522) );
  INV_X1 round_inst_S_5__sbox_inst_com_w_inst_U5 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n505) );
  INV_X1 round_inst_S_5__sbox_inst_com_w_inst_U4 ( .A(round_inst_sin_x[23]), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n486) );
  INV_X1 round_inst_S_5__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_5__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_5__sbox_inst_com_w_inst_n510) );
  INV_X1 round_inst_S_5__sbox_inst_com_w_inst_U2 ( .A(round_inst_sin_x[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_w_inst_n489) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_w_inst_U1 ( .A(round_inst_n45), .B(
        round_inst_sin_z[18]), .Z(round_inst_S_5__sbox_inst_com_w_inst_n402)
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n510), .ZN(round_inst_sout_x[20])
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n509), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n510) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U133 ( .A(round_inst_n47), .B(
        round_inst_sin_y[23]), .ZN(round_inst_S_5__sbox_inst_com_x_inst_n508)
         );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U132 ( .A(round_inst_sin_z[16]), 
        .B(round_inst_S_5__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n506), .Z(round_inst_srout2_x[54]) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U130 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U129 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n503), .A2(round_inst_sin_z[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U127 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U126 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U125 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U124 ( .A1(round_inst_n47), 
        .A2(round_inst_sin_w[20]), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U122 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U121 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U118 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_sin_y[23]), .A2(round_inst_S_5__sbox_inst_com_x_inst_n490), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U115 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n487) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_x_inst_U114 ( .A1(
        round_inst_sin_z[22]), .A2(round_inst_sin_w[20]), .A3(
        round_inst_sin_y[23]), .ZN(round_inst_S_5__sbox_inst_com_x_inst_n489)
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n478), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n476), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n478) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n475), .B(round_inst_sin_z[19]), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n476) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_w[22]), .A2(round_inst_sin_y[23]), .A3(
        round_inst_sin_z[20]), .ZN(round_inst_S_5__sbox_inst_com_x_inst_n475)
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n474), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n473), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n473) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n470), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n469), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n511) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n468), .A2(round_inst_n47), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n469) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n468) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n467), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n464), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_srout2_x[52]) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U100 ( .A1(round_inst_n46), 
        .A2(round_inst_sin_z[22]), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[17]), 
        .B(round_inst_S_5__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n464) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n462), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n460), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n467), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n461) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n458), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n467) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_5__sbox_inst_n1), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n457), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n459) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n455), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n454), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n456) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n453), .A2(round_inst_sin_w[22]), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n454) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n451), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n455) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n450), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n449), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n451) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n448), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n447), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n449) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n446), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_5__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n445), .B(round_inst_n47), .S(
        round_inst_n46), .Z(round_inst_S_5__sbox_inst_com_x_inst_n446) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n444), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n448) );
  MUX2_X1 round_inst_S_5__sbox_inst_com_x_inst_U85 ( .A(round_inst_n47), .B(
        round_inst_sin_z[22]), .S(round_inst_sin_z[20]), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n443), .A2(round_inst_sin_w[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n442), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n441), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n452) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[20]), 
        .A3(round_inst_sin_z[22]), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n441) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n440), .A2(round_inst_sin_w[21]), 
        .A3(round_inst_n47), .ZN(round_inst_S_5__sbox_inst_com_x_inst_n442) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U80 ( .A(round_inst_n46), .B(
        round_inst_sin_z[20]), .Z(round_inst_S_5__sbox_inst_com_x_inst_n440)
         );
  NAND3_X1 round_inst_S_5__sbox_inst_com_x_inst_U79 ( .A1(round_inst_n46), 
        .A2(round_inst_S_5__sbox_inst_com_x_inst_n445), .A3(
        round_inst_S_5__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n460) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U77 ( .A1(round_inst_n46), 
        .A2(round_inst_n47), .ZN(round_inst_S_5__sbox_inst_com_x_inst_n482) );
  AND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U76 ( .A1(round_inst_n47), .A2(
        round_inst_sin_z[20]), .ZN(round_inst_S_5__sbox_inst_com_x_inst_n490)
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n462) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U74 ( .A1(round_inst_n46), 
        .A2(round_inst_sin_w[22]), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n497) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_srout2_x[55]) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n436), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n435), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U71 ( .A(round_inst_n46), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n435) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n434), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n433), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U69 ( .A1(round_inst_sin_z[20]), .A2(round_inst_sin_y[23]), .ZN(round_inst_S_5__sbox_inst_com_x_inst_n433) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n432), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n431), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n434) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n430), .A2(round_inst_n46), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n431) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n429), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n428), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_5__sbox_inst_n1), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n453), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n432) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[18]), 
        .B(round_inst_S_5__sbox_inst_com_x_inst_n438), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n436) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n425), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n424), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n423), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n422), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n421), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n420), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n422) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n419), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n420) );
  NOR3_X1 round_inst_S_5__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n471), .A3(
        round_inst_S_5__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n418) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n416), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n419) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n414), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U53 ( .A1(round_inst_n47), 
        .A2(round_inst_S_5__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n413) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U52 ( .A(round_inst_sin_y[23]), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n414) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n443), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n416) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U50 ( .A1(
        round_inst_S_5__sbox_inst_n1), .A2(round_inst_n47), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n443) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_x_inst_U49 ( .A1(round_inst_n47), 
        .A2(round_inst_S_5__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_5__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n421) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n411), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n423) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U47 ( .A1(round_inst_n47), 
        .A2(round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n465) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n411) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n410), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n407), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U43 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n406), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n405), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n407) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U42 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n466), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n405) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U41 ( .A(round_inst_sin_w[21]), 
        .B(round_inst_S_5__sbox_inst_n1), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n439) );
  AND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U40 ( .A1(round_inst_sin_z[22]), 
        .A2(round_inst_sin_y[23]), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_5__sbox_inst_n3), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n406) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_x_inst_U38 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U37 ( .A(round_inst_sin_z[22]), 
        .B(round_inst_sin_w[22]), .Z(round_inst_S_5__sbox_inst_com_x_inst_n445) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U36 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n404), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n410) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U35 ( .A(round_inst_sin_w[22]), 
        .B(round_inst_n47), .Z(round_inst_S_5__sbox_inst_com_x_inst_n403) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n402), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n401), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U33 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n400), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n399), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n401) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U32 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n399) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U31 ( .A1(round_inst_sin_z[20]), .A2(round_inst_S_5__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n426) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n427), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n400) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U28 ( .A(round_inst_sin_y[23]), 
        .B(round_inst_S_5__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n471) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n402) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_5__sbox_inst_n1), .A3(round_inst_n46), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n396) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n398), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n481) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U23 ( .A(round_inst_sin_y[23]), 
        .B(round_inst_S_5__sbox_inst_n3), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U21 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n392), .A2(round_inst_sin_w[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n404), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_x_inst_U17 ( .A1(round_inst_sin_z[20]), .A2(round_inst_sin_y[23]), .A3(round_inst_sin_w[21]), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n388) );
  MUX2_X1 round_inst_S_5__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n412), .B(round_inst_sin_y[23]), 
        .S(round_inst_S_5__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U15 ( .A1(round_inst_n46), 
        .A2(round_inst_S_5__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U14 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n491), .B(
        round_inst_S_5__sbox_inst_n3), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n412) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n384), .A2(round_inst_sin_z[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U10 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_5__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U9 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_w[23]), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U7 ( .A1(
        round_inst_S_5__sbox_inst_n1), .A2(round_inst_sin_y[23]), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n404) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_5__sbox_inst_com_x_inst_n427), .Z(
        round_inst_S_5__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U4 ( .A1(round_inst_n46), .A2(
        round_inst_sin_w[21]), .ZN(round_inst_S_5__sbox_inst_com_x_inst_n427)
         );
  NAND2_X1 round_inst_S_5__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_5__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_5__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_5__sbox_inst_com_x_inst_n477) );
  INV_X1 round_inst_S_5__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_y[21]), 
        .ZN(round_inst_S_5__sbox_inst_com_x_inst_n417) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n517), .Z(round_inst_sout_y[20])
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n516), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n515) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U134 ( .A(round_inst_sin_x[16]), 
        .B(round_inst_S_5__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n512), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_srout2_y[54]) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n508), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n518) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n507), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n506), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n508) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n506) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n507) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_5__sbox_inst_com_y_inst_U125 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_5__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U124 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U123 ( .A1(
        round_inst_sin_x[23]), .A2(round_inst_S_5__sbox_inst_com_y_inst_n493), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n492), .A2(
        round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U121 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U120 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U119 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U118 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n486), .A2(
        round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U117 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n503), .A2(round_inst_sin_w[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U112 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_5__sbox_inst_n1), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[19]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_y_inst_U109 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_5__sbox_inst_n3), .A3(round_inst_sin_x[20]), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U108 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_y_inst_U107 ( .A1(
        round_inst_sin_w[20]), .A2(round_inst_sin_w[23]), .A3(
        round_inst_S_5__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_5__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_5__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U105 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[52]) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U104 ( .A1(
        round_inst_S_5__sbox_inst_n5), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U98 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_5__sbox_inst_n1), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U95 ( .A1(round_inst_sin_x[20]), .A2(round_inst_S_5__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_y_inst_U94 ( .A1(round_inst_sin_w[20]), .A2(round_inst_n63), .A3(round_inst_S_5__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U93 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U92 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U88 ( .A1(
        round_inst_S_5__sbox_inst_n1), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_5__sbox_inst_com_y_inst_U87 ( .A(
        round_inst_S_5__sbox_inst_n5), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n503), .S(
        round_inst_S_5__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_5__sbox_inst_n1), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n478), .B(round_inst_n62), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n438), .Z(round_inst_srout2_y[55]) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U71 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[23]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U70 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n483), .A2(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_5__sbox_inst_n1), .A2(round_inst_sin_w[20]), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[23]), 
        .A3(round_inst_S_5__sbox_inst_n1), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U66 ( .A(round_inst_sin_w[20]), 
        .B(round_inst_sin_x[20]), .Z(round_inst_S_5__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U59 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[23]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U58 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[21]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U55 ( .A(round_inst_sin_x[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U54 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n418), .A2(
        round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U53 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U51 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U50 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n414), .B(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U49 ( .A(round_inst_sin_w[21]), 
        .B(round_inst_S_5__sbox_inst_n1), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U48 ( .A1(
        round_inst_S_5__sbox_inst_n1), .A2(round_inst_sin_x[20]), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_5__sbox_inst_n1), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U46 ( .A(round_inst_sin_x[18]), 
        .B(round_inst_S_5__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n513) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[21]), 
        .B(round_inst_sin_x[23]), .Z(round_inst_S_5__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U41 ( .A(round_inst_n63), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[23]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[20]), 
        .Z(round_inst_S_5__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U36 ( .A(round_inst_sin_z[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_5__sbox_inst_n1), .B(round_inst_S_5__sbox_inst_n3), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_5__sbox_inst_n5), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U27 ( .A1(round_inst_sin_w[21]), .A2(round_inst_S_5__sbox_inst_n3), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n514), .A2(round_inst_sin_w[21]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_5__sbox_inst_n1), .A2(round_inst_sin_w[23]), .A3(
        round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_5__sbox_inst_n1), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n504), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_5__sbox_inst_n3), .B(round_inst_sin_w[23]), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U17 ( .A(
        round_inst_S_5__sbox_inst_n3), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[23]), 
        .B(round_inst_sin_x[23]), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_y_inst_U13 ( .A1(round_inst_n63), 
        .A2(round_inst_sin_w[23]), .A3(
        round_inst_S_5__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_y_inst_U12 ( .A1(
        round_inst_S_5__sbox_inst_n3), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_5__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[21]), 
        .B(round_inst_n63), .S(round_inst_S_5__sbox_inst_com_y_inst_n503), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_y_inst_U9 ( .A1(round_inst_n63), .A2(
        round_inst_S_5__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_5__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_5__sbox_inst_n3), .B(round_inst_sin_x[23]), .Z(
        round_inst_S_5__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_5__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_5__sbox_inst_n1), .A3(round_inst_sin_x[23]), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_5__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n503) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[22]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_5__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_5__sbox_inst_com_y_inst_n514) );
  INV_X1 round_inst_S_5__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[22]), 
        .ZN(round_inst_S_5__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n516), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n515), .ZN(round_inst_sout_z[20])
         );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n514), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n513), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_w[22]), .B(round_inst_sin_w[23]), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n513) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U128 ( .A(round_inst_sin_x[16]), 
        .B(round_inst_n44), .Z(round_inst_S_5__sbox_inst_com_z_inst_n514) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n510), .ZN(
        round_inst_srout2_z[54]) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n509), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n508), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U124 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n507), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n506), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n508) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U123 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n505), .A2(round_inst_n46), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n506) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n504), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n503), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n502), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n501), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n503) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U120 ( .A(round_inst_sin_w[21]), .B(round_inst_sin_x[19]), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n501) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U119 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n500), .B(round_inst_sin_y[19]), 
        .Z(round_inst_S_5__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U118 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n499), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n498), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n500) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U117 ( .A1(round_inst_n47), 
        .A2(round_inst_S_5__sbox_inst_com_z_inst_n497), .A3(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n498) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U116 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n495), .A2(round_inst_sin_x[20]), 
        .A3(round_inst_sin_w[23]), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n499) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U115 ( .A(
        round_inst_S_5__sbox_inst_n5), .B(round_inst_n47), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n495) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U114 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_5__sbox_inst_n5), .A3(round_inst_sin_x[23]), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n509) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n491), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n493) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U111 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n490), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n489), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n491) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n488), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n486), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n490) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U108 ( .A1(
        round_inst_sin_w[22]), .A2(round_inst_sin_x[23]), .A3(round_inst_n46), 
        .ZN(round_inst_S_5__sbox_inst_com_z_inst_n492) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U107 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n484), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U106 ( .A1(
        round_inst_sin_w[22]), .A2(round_inst_S_5__sbox_inst_com_z_inst_n497), 
        .ZN(round_inst_S_5__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n505), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n484) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n482), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n481), .Z(round_inst_srout2_z[52]) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n479), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n478), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n483), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U101 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n483) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U100 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n475), .A2(round_inst_sin_x[20]), 
        .A3(round_inst_sin_w[22]), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U99 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n474), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n477) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U98 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n472), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .A3(round_inst_n47), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n473) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U97 ( .A(round_inst_sin_w[21]), 
        .B(round_inst_sin_y[21]), .Z(round_inst_S_5__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U96 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n471), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n474) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U95 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n469), .A2(
        round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n470) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n467), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n471) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n466), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n465), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n464), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n463), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U91 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n462), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n461), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U90 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n460), .A2(round_inst_n47), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n461) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U89 ( .A1(round_inst_n63), 
        .A2(round_inst_S_5__sbox_inst_n5), .A3(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n462) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n459), .A2(round_inst_n46), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U87 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_w[22]), 
        .ZN(round_inst_S_5__sbox_inst_com_z_inst_n466) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U85 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U84 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n453), .A2(round_inst_n47), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n454) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U83 ( .A(round_inst_sin_w[21]), 
        .B(round_inst_S_5__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n451), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U81 ( .A1(round_inst_sin_w[22]), .A2(round_inst_sin_x[20]), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n478) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U79 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n487), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n448) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U78 ( .A(round_inst_sin_y[17]), 
        .B(round_inst_n62), .Z(round_inst_S_5__sbox_inst_com_z_inst_n447) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n487) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U76 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n446), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U75 ( .A(round_inst_sin_w[22]), 
        .B(round_inst_n47), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_srout2_z[55]) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n511), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U72 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n511) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U71 ( .A1(round_inst_sin_x[20]), .A2(round_inst_sin_w[23]), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n441) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U70 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n458), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n440), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n442) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U69 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U68 ( .A(round_inst_sin_w[23]), 
        .B(round_inst_S_5__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n497) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n494) );
  MUX2_X1 round_inst_S_5__sbox_inst_com_z_inst_U66 ( .A(round_inst_sin_x[23]), 
        .B(round_inst_sin_w[23]), .S(round_inst_S_5__sbox_inst_com_z_inst_n436), .Z(round_inst_S_5__sbox_inst_com_z_inst_n437) );
  OR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U65 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n436) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U64 ( .A(round_inst_sin_x[20]), 
        .B(round_inst_S_5__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n486) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U63 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n438) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U62 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_x[23]), 
        .A3(round_inst_S_5__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n430), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U59 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n429) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U58 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n426), .A2(round_inst_sin_w[23]), 
        .ZN(round_inst_S_5__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U56 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n422), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n424) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U55 ( .A1(round_inst_sin_x[20]), .A2(round_inst_n63), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U54 ( .A1(round_inst_sin_y[21]), .A2(round_inst_sin_x[20]), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n425) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U53 ( .A1(round_inst_n46), 
        .A2(round_inst_sin_x[23]), .A3(round_inst_sin_w[21]), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n428) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U52 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_y[23]), 
        .ZN(round_inst_S_5__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U50 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n460), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n423), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n469) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U49 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_y[21]), 
        .ZN(round_inst_S_5__sbox_inst_com_z_inst_n423) );
  AND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U48 ( .A1(round_inst_sin_w[21]), 
        .A2(round_inst_sin_x[20]), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n460) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U47 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n421) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U46 ( .A1(round_inst_sin_w[21]), .A2(round_inst_S_5__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .A2(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U44 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n419), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n418), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n432) );
  INV_X1 round_inst_S_5__sbox_inst_com_z_inst_U43 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .B(round_inst_n46), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n451) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U41 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n417), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n496), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U39 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n449) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U38 ( .A1(round_inst_sin_w[23]), .A2(round_inst_S_5__sbox_inst_com_z_inst_n413), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n414) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n415) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U35 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U34 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n505), .A2(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n409) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U32 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n407) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n405) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U30 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n404) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n505), .A2(round_inst_sin_y[21]), 
        .ZN(round_inst_S_5__sbox_inst_com_z_inst_n402) );
  AND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_S_5__sbox_inst_n5), .A2(round_inst_sin_w[23]), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n505) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U27 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n401), .A2(round_inst_n47), .A3(
        round_inst_sin_w[21]), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n403)
         );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U26 ( .A(round_inst_sin_w[23]), 
        .B(round_inst_sin_x[23]), .Z(round_inst_S_5__sbox_inst_com_z_inst_n401) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U25 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n399), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n406) );
  MUX2_X1 round_inst_S_5__sbox_inst_com_z_inst_U24 ( .A(round_inst_sin_y[23]), 
        .B(round_inst_S_5__sbox_inst_com_z_inst_n398), .S(
        round_inst_S_5__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U23 ( .A1(round_inst_sin_w[21]), .A2(round_inst_S_5__sbox_inst_n5), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n398) );
  INV_X1 round_inst_S_5__sbox_inst_com_z_inst_U21 ( .A(round_inst_sin_x[23]), 
        .ZN(round_inst_S_5__sbox_inst_com_z_inst_n397) );
  NOR3_X1 round_inst_S_5__sbox_inst_com_z_inst_U20 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n488), .A3(
        round_inst_S_5__sbox_inst_com_z_inst_n395), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U19 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n394), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n395) );
  INV_X1 round_inst_S_5__sbox_inst_com_z_inst_U18 ( .A(round_inst_n63), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n394) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U17 ( .A(round_inst_sin_w[23]), 
        .B(round_inst_sin_y[23]), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n488) );
  AND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U16 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n459), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U15 ( .A1(round_inst_sin_w[22]), .A2(round_inst_n63), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n459) );
  INV_X1 round_inst_S_5__sbox_inst_com_z_inst_U14 ( .A(round_inst_sin_w[21]), 
        .ZN(round_inst_S_5__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U13 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n393), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U12 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n391), .A2(round_inst_n47), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U11 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_5__sbox_inst_com_z_inst_n390), .Z(
        round_inst_S_5__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U10 ( .A1(round_inst_sin_w[21]), .A2(round_inst_sin_y[23]), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n390) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U9 ( .A1(round_inst_n63), .A2(
        round_inst_sin_w[23]), .ZN(round_inst_S_5__sbox_inst_com_z_inst_n418)
         );
  NOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U8 ( .A1(
        round_inst_S_5__sbox_inst_com_z_inst_n439), .A2(
        round_inst_S_5__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_5__sbox_inst_com_z_inst_U7 ( .A1(round_inst_sin_w[22]), 
        .A2(round_inst_sin_w[21]), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n456) );
  XNOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U6 ( .A(round_inst_sin_x[23]), 
        .B(round_inst_sin_y[23]), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n439) );
  NAND3_X1 round_inst_S_5__sbox_inst_com_z_inst_U5 ( .A1(round_inst_sin_w[22]), 
        .A2(round_inst_sin_x[23]), .A3(
        round_inst_S_5__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U4 ( .A(round_inst_n63), .B(
        round_inst_sin_y[21]), .Z(round_inst_S_5__sbox_inst_com_z_inst_n475)
         );
  INV_X1 round_inst_S_5__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_5__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_5__sbox_inst_com_z_inst_n496) );
  INV_X1 round_inst_S_5__sbox_inst_com_z_inst_U2 ( .A(round_inst_sin_w[20]), 
        .ZN(round_inst_S_5__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_5__sbox_inst_com_z_inst_U1 ( .A(round_inst_n45), .B(
        round_inst_sin_x[18]), .Z(round_inst_S_5__sbox_inst_com_z_inst_n417)
         );
  INV_X1 round_inst_S_6__sbox_inst_U6 ( .A(round_inst_sin_x[26]), .ZN(
        round_inst_S_6__sbox_inst_n6) );
  INV_X1 round_inst_S_6__sbox_inst_U5 ( .A(round_inst_sin_z[25]), .ZN(
        round_inst_S_6__sbox_inst_n2) );
  INV_X1 round_inst_S_6__sbox_inst_U4 ( .A(round_inst_sin_z[27]), .ZN(
        round_inst_S_6__sbox_inst_n4) );
  INV_X2 round_inst_S_6__sbox_inst_U3 ( .A(round_inst_S_6__sbox_inst_n4), .ZN(
        round_inst_S_6__sbox_inst_n3) );
  INV_X2 round_inst_S_6__sbox_inst_U2 ( .A(round_inst_S_6__sbox_inst_n2), .ZN(
        round_inst_S_6__sbox_inst_n1) );
  INV_X2 round_inst_S_6__sbox_inst_U1 ( .A(round_inst_S_6__sbox_inst_n6), .ZN(
        round_inst_S_6__sbox_inst_n5) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n531), .ZN(round_inst_sout_w[27])
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U139 ( .A1(
        round_inst_sin_z[24]), .A2(round_inst_S_6__sbox_inst_com_w_inst_n528), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n526), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n524), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n526) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[26]), .A2(round_inst_S_6__sbox_inst_com_w_inst_n523), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n525) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n518), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n516), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n518) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n514), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n513), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n512), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n513) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_w_inst_U128 ( .A1(
        round_inst_S_6__sbox_inst_n5), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n510), .A3(
        round_inst_S_6__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n511) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U127 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n508), .A2(round_inst_n48), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n507), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U125 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n507) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_6__sbox_inst_n3), .A2(round_inst_n49), .A3(
        round_inst_S_6__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U122 ( .A(round_inst_sin_y[23]), .B(round_inst_S_6__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U121 ( .A(round_inst_n64), .B(
        round_inst_sin_z[23]), .Z(round_inst_S_6__sbox_inst_com_w_inst_n501)
         );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U120 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[25])
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[21]), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[21]), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U113 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[24])
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_6__sbox_inst_n5), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U110 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n528), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U105 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_6__sbox_inst_n5), .B(round_inst_sin_z[26]), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_6__sbox_inst_n1), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U99 ( .A1(round_inst_n49), 
        .A2(round_inst_S_6__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_6__sbox_inst_n5), .A2(round_inst_n48), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n506) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U94 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[26]), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n461), .A2(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[26]), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U88 ( .A1(round_inst_sin_z[24]), 
        .A2(round_inst_S_6__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_w_inst_U85 ( .A1(round_inst_sin_y[25]), .A2(round_inst_n48), .A3(round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_w_inst_U84 ( .A1(round_inst_n49), 
        .A2(round_inst_n64), .A3(round_inst_n48), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n528) );
  OR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_6__sbox_inst_n5), .B(round_inst_n49), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U80 ( .A(round_inst_n46), .B(
        round_inst_sin_z[20]), .Z(round_inst_S_6__sbox_inst_com_w_inst_n484)
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U79 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[27])
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U73 ( .A1(
        round_inst_S_6__sbox_inst_n3), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U71 ( .A1(round_inst_n49), 
        .A2(round_inst_n64), .ZN(round_inst_S_6__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_6__sbox_inst_n5), .A2(round_inst_sin_y[25]), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U69 ( .A1(
        round_inst_S_6__sbox_inst_n1), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n508), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_6__sbox_inst_n5), .A2(round_inst_S_6__sbox_inst_n1), .A3(
        round_inst_S_6__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n439), .A2(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n508), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_6__sbox_inst_n3), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n504) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U62 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n508) );
  INV_X1 round_inst_S_6__sbox_inst_com_w_inst_U61 ( .A(round_inst_n49), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U60 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U58 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U57 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U56 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U55 ( .A(round_inst_sin_y[25]), 
        .B(round_inst_S_6__sbox_inst_n1), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U54 ( .A1(
        round_inst_S_6__sbox_inst_n3), .A2(round_inst_S_6__sbox_inst_n1), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U52 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_w_inst_U51 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n505), .A3(
        round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U50 ( .A(round_inst_sin_y[25]), 
        .B(round_inst_n64), .Z(round_inst_S_6__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_w_inst_U49 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n505), .A2(round_inst_sin_y[25]), 
        .A3(round_inst_S_6__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U48 ( .A(round_inst_n49), .B(
        round_inst_sin_z[26]), .ZN(round_inst_S_6__sbox_inst_com_w_inst_n465)
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U47 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n520) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U45 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n421), .A2(
        round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U44 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U43 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n419), .A2(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U42 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U40 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_6__sbox_inst_n1), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n521) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U38 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U37 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U36 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n510), .B(round_inst_sin_z[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n498), .A2(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U33 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U32 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U31 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U30 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U29 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U28 ( .A1(round_inst_n64), 
        .A2(round_inst_sin_z[24]), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U27 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n522), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U26 ( .A(round_inst_n64), .B(
        round_inst_S_6__sbox_inst_n1), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U24 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n510), .A2(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U22 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[25]), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U21 ( .A(round_inst_n48), .B(
        round_inst_sin_z[24]), .Z(round_inst_S_6__sbox_inst_com_w_inst_n418)
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U20 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U19 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U17 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n398), .A2(
        round_inst_S_6__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U15 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n498), .B(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_6__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_6__sbox_inst_com_w_inst_U13 ( .A(round_inst_sin_y[27]), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_6__sbox_inst_n1), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U11 ( .A(
        round_inst_S_6__sbox_inst_n3), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n505), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U9 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_6__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_6__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U8 ( .A1(round_inst_n64), .A2(
        round_inst_n48), .ZN(round_inst_S_6__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U7 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n510), .A2(round_inst_sin_y[25]), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n477) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_w_inst_U6 ( .A1(
        round_inst_S_6__sbox_inst_com_w_inst_n505), .A2(round_inst_n48), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n522) );
  INV_X1 round_inst_S_6__sbox_inst_com_w_inst_U5 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n505) );
  INV_X1 round_inst_S_6__sbox_inst_com_w_inst_U4 ( .A(round_inst_sin_x[27]), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n486) );
  INV_X1 round_inst_S_6__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_6__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_6__sbox_inst_com_w_inst_n510) );
  INV_X1 round_inst_S_6__sbox_inst_com_w_inst_U2 ( .A(round_inst_sin_x[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_w_inst_n489) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_w_inst_U1 ( .A(round_inst_n47), .B(
        round_inst_sin_z[22]), .Z(round_inst_S_6__sbox_inst_com_w_inst_n402)
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n510), .ZN(round_inst_sout_x[24])
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n509), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n510) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U133 ( .A(round_inst_n49), .B(
        round_inst_sin_y[27]), .ZN(round_inst_S_6__sbox_inst_com_x_inst_n508)
         );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U132 ( .A(round_inst_sin_z[20]), 
        .B(round_inst_S_6__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n506), .Z(round_inst_srout2_x[10]) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U130 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U129 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n503), .A2(round_inst_sin_z[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U127 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U126 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U125 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U124 ( .A1(round_inst_n49), 
        .A2(round_inst_sin_w[24]), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U122 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U121 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U118 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_sin_y[27]), .A2(round_inst_S_6__sbox_inst_com_x_inst_n490), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U115 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n487) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_x_inst_U114 ( .A1(
        round_inst_sin_z[26]), .A2(round_inst_sin_w[24]), .A3(
        round_inst_sin_y[27]), .ZN(round_inst_S_6__sbox_inst_com_x_inst_n489)
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n478), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n476), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n478) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n475), .B(round_inst_sin_z[23]), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n476) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_w[26]), .A2(round_inst_sin_y[27]), .A3(
        round_inst_sin_z[24]), .ZN(round_inst_S_6__sbox_inst_com_x_inst_n475)
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n474), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n473), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n473) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n470), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n469), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n511) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n468), .A2(round_inst_n49), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n469) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n468) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n467), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n464), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n480), .ZN(round_inst_srout2_x[8]) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U100 ( .A1(round_inst_n48), 
        .A2(round_inst_sin_z[26]), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[21]), 
        .B(round_inst_S_6__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n464) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n462), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n460), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n467), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n461) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n458), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n467) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_6__sbox_inst_n1), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n457), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n459) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n455), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n454), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n456) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n453), .A2(round_inst_sin_w[26]), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n454) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n451), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n455) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n450), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n449), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n451) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n448), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n447), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n449) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n446), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_6__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n445), .B(round_inst_n49), .S(
        round_inst_n48), .Z(round_inst_S_6__sbox_inst_com_x_inst_n446) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n444), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n448) );
  MUX2_X1 round_inst_S_6__sbox_inst_com_x_inst_U85 ( .A(round_inst_n49), .B(
        round_inst_sin_z[26]), .S(round_inst_sin_z[24]), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n443), .A2(round_inst_sin_w[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n442), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n441), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n452) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[24]), 
        .A3(round_inst_sin_z[26]), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n441) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n440), .A2(round_inst_sin_w[25]), 
        .A3(round_inst_n49), .ZN(round_inst_S_6__sbox_inst_com_x_inst_n442) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U80 ( .A(round_inst_n48), .B(
        round_inst_sin_z[24]), .Z(round_inst_S_6__sbox_inst_com_x_inst_n440)
         );
  NAND3_X1 round_inst_S_6__sbox_inst_com_x_inst_U79 ( .A1(round_inst_n48), 
        .A2(round_inst_S_6__sbox_inst_com_x_inst_n445), .A3(
        round_inst_S_6__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n460) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U77 ( .A1(round_inst_n48), 
        .A2(round_inst_n49), .ZN(round_inst_S_6__sbox_inst_com_x_inst_n482) );
  AND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U76 ( .A1(round_inst_n49), .A2(
        round_inst_sin_z[24]), .ZN(round_inst_S_6__sbox_inst_com_x_inst_n490)
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n462) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U74 ( .A1(round_inst_n48), 
        .A2(round_inst_sin_w[26]), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n497) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_srout2_x[11]) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n436), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n435), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U71 ( .A(round_inst_n48), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n435) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n434), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n433), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U69 ( .A1(round_inst_sin_z[24]), .A2(round_inst_sin_y[27]), .ZN(round_inst_S_6__sbox_inst_com_x_inst_n433) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n432), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n431), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n434) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n430), .A2(round_inst_n48), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n431) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n429), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n428), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_6__sbox_inst_n1), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n453), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n432) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[22]), 
        .B(round_inst_S_6__sbox_inst_com_x_inst_n438), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n436) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n425), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n424), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n423), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n422), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n421), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n420), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n422) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n419), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n420) );
  NOR3_X1 round_inst_S_6__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n471), .A3(
        round_inst_S_6__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n418) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n416), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n419) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n414), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U53 ( .A1(round_inst_n49), 
        .A2(round_inst_S_6__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n413) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U52 ( .A(round_inst_sin_y[27]), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n414) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n443), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n416) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U50 ( .A1(
        round_inst_S_6__sbox_inst_n1), .A2(round_inst_n49), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n443) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_x_inst_U49 ( .A1(round_inst_n49), 
        .A2(round_inst_S_6__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_6__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n421) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n411), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n423) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U47 ( .A1(round_inst_n49), 
        .A2(round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n465) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n411) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n410), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n407), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U43 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n406), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n405), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n407) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U42 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n466), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n405) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U41 ( .A(round_inst_sin_w[25]), 
        .B(round_inst_S_6__sbox_inst_n1), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n439) );
  AND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U40 ( .A1(round_inst_sin_z[26]), 
        .A2(round_inst_sin_y[27]), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_6__sbox_inst_n3), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n406) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_x_inst_U38 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U37 ( .A(round_inst_sin_z[26]), 
        .B(round_inst_sin_w[26]), .Z(round_inst_S_6__sbox_inst_com_x_inst_n445) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U36 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n404), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n410) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U35 ( .A(round_inst_sin_w[26]), 
        .B(round_inst_n49), .Z(round_inst_S_6__sbox_inst_com_x_inst_n403) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n402), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n401), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U33 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n400), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n399), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n401) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U32 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n399) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U31 ( .A1(round_inst_sin_z[24]), .A2(round_inst_S_6__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n426) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n427), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n400) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U28 ( .A(round_inst_sin_y[27]), 
        .B(round_inst_S_6__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n471) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n402) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_6__sbox_inst_n1), .A3(round_inst_n48), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n396) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n398), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n481) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U23 ( .A(round_inst_sin_y[27]), 
        .B(round_inst_S_6__sbox_inst_n3), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U21 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n392), .A2(round_inst_sin_w[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n404), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_x_inst_U17 ( .A1(round_inst_sin_z[24]), .A2(round_inst_sin_y[27]), .A3(round_inst_sin_w[25]), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n388) );
  MUX2_X1 round_inst_S_6__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n412), .B(round_inst_sin_y[27]), 
        .S(round_inst_S_6__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U15 ( .A1(round_inst_n48), 
        .A2(round_inst_S_6__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U14 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n491), .B(
        round_inst_S_6__sbox_inst_n3), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n412) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n384), .A2(round_inst_sin_z[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U10 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_6__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U9 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_w[27]), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U7 ( .A1(
        round_inst_S_6__sbox_inst_n1), .A2(round_inst_sin_y[27]), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n404) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_6__sbox_inst_com_x_inst_n427), .Z(
        round_inst_S_6__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U4 ( .A1(round_inst_n48), .A2(
        round_inst_sin_w[25]), .ZN(round_inst_S_6__sbox_inst_com_x_inst_n427)
         );
  NAND2_X1 round_inst_S_6__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_6__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_6__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_6__sbox_inst_com_x_inst_n477) );
  INV_X1 round_inst_S_6__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_y[25]), 
        .ZN(round_inst_S_6__sbox_inst_com_x_inst_n417) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n517), .Z(round_inst_sout_y[24])
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n516), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n515) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U134 ( .A(round_inst_sin_x[20]), 
        .B(round_inst_S_6__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n512), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_srout2_y[10]) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n508), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n518) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n507), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n506), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n508) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n506) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n507) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_6__sbox_inst_com_y_inst_U125 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_6__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U124 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U123 ( .A1(
        round_inst_sin_x[27]), .A2(round_inst_S_6__sbox_inst_com_y_inst_n493), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n492), .A2(
        round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U121 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U120 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U119 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U118 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n486), .A2(
        round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U117 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n503), .A2(round_inst_sin_w[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U112 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_6__sbox_inst_n1), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[23]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_y_inst_U109 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_6__sbox_inst_n3), .A3(round_inst_sin_x[24]), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U108 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_y_inst_U107 ( .A1(
        round_inst_sin_w[24]), .A2(round_inst_sin_w[27]), .A3(
        round_inst_S_6__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_6__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_6__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U105 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n470), .ZN(round_inst_srout2_y[8]) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U104 ( .A1(
        round_inst_S_6__sbox_inst_n5), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U98 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_6__sbox_inst_n1), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U95 ( .A1(round_inst_sin_x[24]), .A2(round_inst_S_6__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_y_inst_U94 ( .A1(round_inst_sin_w[24]), .A2(round_inst_n64), .A3(round_inst_S_6__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U93 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U92 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U88 ( .A1(
        round_inst_S_6__sbox_inst_n1), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_6__sbox_inst_com_y_inst_U87 ( .A(
        round_inst_S_6__sbox_inst_n5), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n503), .S(
        round_inst_S_6__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_6__sbox_inst_n1), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n478), .B(round_inst_n63), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n438), .Z(round_inst_srout2_y[11]) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U71 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[27]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U70 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n483), .A2(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_6__sbox_inst_n1), .A2(round_inst_sin_w[24]), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[27]), 
        .A3(round_inst_S_6__sbox_inst_n1), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U66 ( .A(round_inst_sin_w[24]), 
        .B(round_inst_sin_x[24]), .Z(round_inst_S_6__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U59 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[27]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U58 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[25]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U55 ( .A(round_inst_sin_x[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U54 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n418), .A2(
        round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U53 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U51 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U50 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n414), .B(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U49 ( .A(round_inst_sin_w[25]), 
        .B(round_inst_S_6__sbox_inst_n1), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U48 ( .A1(
        round_inst_S_6__sbox_inst_n1), .A2(round_inst_sin_x[24]), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_6__sbox_inst_n1), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U46 ( .A(round_inst_sin_x[22]), 
        .B(round_inst_S_6__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n513) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[25]), 
        .B(round_inst_sin_x[27]), .Z(round_inst_S_6__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U41 ( .A(round_inst_n64), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[27]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[24]), 
        .Z(round_inst_S_6__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U36 ( .A(round_inst_sin_z[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_6__sbox_inst_n1), .B(round_inst_S_6__sbox_inst_n3), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_6__sbox_inst_n5), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U27 ( .A1(round_inst_sin_w[25]), .A2(round_inst_S_6__sbox_inst_n3), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n514), .A2(round_inst_sin_w[25]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_6__sbox_inst_n1), .A2(round_inst_sin_w[27]), .A3(
        round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_6__sbox_inst_n1), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n504), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_6__sbox_inst_n3), .B(round_inst_sin_w[27]), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U17 ( .A(
        round_inst_S_6__sbox_inst_n3), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[27]), 
        .B(round_inst_sin_x[27]), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_y_inst_U13 ( .A1(round_inst_n64), 
        .A2(round_inst_sin_w[27]), .A3(
        round_inst_S_6__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_y_inst_U12 ( .A1(
        round_inst_S_6__sbox_inst_n3), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_6__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[25]), 
        .B(round_inst_n64), .S(round_inst_S_6__sbox_inst_com_y_inst_n503), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_y_inst_U9 ( .A1(round_inst_n64), .A2(
        round_inst_S_6__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_6__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_6__sbox_inst_n3), .B(round_inst_sin_x[27]), .Z(
        round_inst_S_6__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_6__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_6__sbox_inst_n1), .A3(round_inst_sin_x[27]), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_6__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n503) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[26]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_6__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_6__sbox_inst_com_y_inst_n514) );
  INV_X1 round_inst_S_6__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[26]), 
        .ZN(round_inst_S_6__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n516), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n515), .ZN(round_inst_sout_z[24])
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n514), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n513), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_w[26]), .B(round_inst_sin_w[27]), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n513) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U128 ( .A(round_inst_sin_x[20]), 
        .B(round_inst_n46), .Z(round_inst_S_6__sbox_inst_com_z_inst_n514) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n510), .ZN(
        round_inst_srout2_z[10]) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n509), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n508), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U124 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n507), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n506), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n508) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U123 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n505), .A2(round_inst_n48), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n506) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n504), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n503), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n502), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n501), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n503) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U120 ( .A(round_inst_sin_w[25]), .B(round_inst_sin_x[23]), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n501) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U119 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n500), .B(round_inst_sin_y[23]), 
        .Z(round_inst_S_6__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U118 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n499), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n498), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n500) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U117 ( .A1(round_inst_n49), 
        .A2(round_inst_S_6__sbox_inst_com_z_inst_n497), .A3(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n498) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U116 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n495), .A2(round_inst_sin_x[24]), 
        .A3(round_inst_sin_w[27]), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n499) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U115 ( .A(
        round_inst_S_6__sbox_inst_n5), .B(round_inst_n49), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n495) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U114 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_6__sbox_inst_n5), .A3(round_inst_sin_x[27]), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n509) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n491), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n493) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U111 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n490), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n489), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n491) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n488), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n486), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n490) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U108 ( .A1(
        round_inst_sin_w[26]), .A2(round_inst_sin_x[27]), .A3(round_inst_n48), 
        .ZN(round_inst_S_6__sbox_inst_com_z_inst_n492) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U107 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n484), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U106 ( .A1(
        round_inst_sin_w[26]), .A2(round_inst_S_6__sbox_inst_com_z_inst_n497), 
        .ZN(round_inst_S_6__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n505), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n484) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n482), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n481), .Z(round_inst_srout2_z[8])
         );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n479), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n478), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n483), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U101 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n483) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U100 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n475), .A2(round_inst_sin_x[24]), 
        .A3(round_inst_sin_w[26]), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U99 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n474), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n477) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U98 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n472), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .A3(round_inst_n49), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n473) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U97 ( .A(round_inst_sin_w[25]), 
        .B(round_inst_sin_y[25]), .Z(round_inst_S_6__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U96 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n471), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n474) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U95 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n469), .A2(
        round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n470) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n467), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n471) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n466), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n465), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n464), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n463), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U91 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n462), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n461), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U90 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n460), .A2(round_inst_n49), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n461) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U89 ( .A1(round_inst_n64), 
        .A2(round_inst_S_6__sbox_inst_n5), .A3(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n462) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n459), .A2(round_inst_n48), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U87 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_w[26]), 
        .ZN(round_inst_S_6__sbox_inst_com_z_inst_n466) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U85 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U84 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n453), .A2(round_inst_n49), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n454) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U83 ( .A(round_inst_sin_w[25]), 
        .B(round_inst_S_6__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n451), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U81 ( .A1(round_inst_sin_w[26]), .A2(round_inst_sin_x[24]), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n478) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U79 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n487), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n448) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U78 ( .A(round_inst_sin_y[21]), 
        .B(round_inst_n63), .Z(round_inst_S_6__sbox_inst_com_z_inst_n447) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n487) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U76 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n446), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U75 ( .A(round_inst_sin_w[26]), 
        .B(round_inst_n49), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_srout2_z[11]) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n511), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U72 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n511) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U71 ( .A1(round_inst_sin_x[24]), .A2(round_inst_sin_w[27]), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n441) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U70 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n458), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n440), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n442) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U69 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U68 ( .A(round_inst_sin_w[27]), 
        .B(round_inst_S_6__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n497) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n494) );
  MUX2_X1 round_inst_S_6__sbox_inst_com_z_inst_U66 ( .A(round_inst_sin_x[27]), 
        .B(round_inst_sin_w[27]), .S(round_inst_S_6__sbox_inst_com_z_inst_n436), .Z(round_inst_S_6__sbox_inst_com_z_inst_n437) );
  OR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U65 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n436) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U64 ( .A(round_inst_sin_x[24]), 
        .B(round_inst_S_6__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n486) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U63 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n438) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U62 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_x[27]), 
        .A3(round_inst_S_6__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n430), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U59 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n429) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U58 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n426), .A2(round_inst_sin_w[27]), 
        .ZN(round_inst_S_6__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U56 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n422), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n424) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U55 ( .A1(round_inst_sin_x[24]), .A2(round_inst_n64), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U54 ( .A1(round_inst_sin_y[25]), .A2(round_inst_sin_x[24]), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n425) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U53 ( .A1(round_inst_n48), 
        .A2(round_inst_sin_x[27]), .A3(round_inst_sin_w[25]), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n428) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U52 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_y[27]), 
        .ZN(round_inst_S_6__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U50 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n460), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n423), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n469) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U49 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_y[25]), 
        .ZN(round_inst_S_6__sbox_inst_com_z_inst_n423) );
  AND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U48 ( .A1(round_inst_sin_w[25]), 
        .A2(round_inst_sin_x[24]), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n460) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U47 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n421) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U46 ( .A1(round_inst_sin_w[25]), .A2(round_inst_S_6__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .A2(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U44 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n419), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n418), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n432) );
  INV_X1 round_inst_S_6__sbox_inst_com_z_inst_U43 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .B(round_inst_n48), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n451) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U41 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n417), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n496), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U39 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n449) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U38 ( .A1(round_inst_sin_w[27]), .A2(round_inst_S_6__sbox_inst_com_z_inst_n413), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n414) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n415) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U35 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U34 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n505), .A2(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n409) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U32 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n407) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n405) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U30 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n404) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n505), .A2(round_inst_sin_y[25]), 
        .ZN(round_inst_S_6__sbox_inst_com_z_inst_n402) );
  AND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_S_6__sbox_inst_n5), .A2(round_inst_sin_w[27]), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n505) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U27 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n401), .A2(round_inst_n49), .A3(
        round_inst_sin_w[25]), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n403)
         );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U26 ( .A(round_inst_sin_w[27]), 
        .B(round_inst_sin_x[27]), .Z(round_inst_S_6__sbox_inst_com_z_inst_n401) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U25 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n399), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n406) );
  MUX2_X1 round_inst_S_6__sbox_inst_com_z_inst_U24 ( .A(round_inst_sin_y[27]), 
        .B(round_inst_S_6__sbox_inst_com_z_inst_n398), .S(
        round_inst_S_6__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U23 ( .A1(round_inst_sin_w[25]), .A2(round_inst_S_6__sbox_inst_n5), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n398) );
  INV_X1 round_inst_S_6__sbox_inst_com_z_inst_U21 ( .A(round_inst_sin_x[27]), 
        .ZN(round_inst_S_6__sbox_inst_com_z_inst_n397) );
  NOR3_X1 round_inst_S_6__sbox_inst_com_z_inst_U20 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n488), .A3(
        round_inst_S_6__sbox_inst_com_z_inst_n395), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U19 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n394), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n395) );
  INV_X1 round_inst_S_6__sbox_inst_com_z_inst_U18 ( .A(round_inst_n64), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n394) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U17 ( .A(round_inst_sin_w[27]), 
        .B(round_inst_sin_y[27]), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n488) );
  AND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U16 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n459), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U15 ( .A1(round_inst_sin_w[26]), .A2(round_inst_n64), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n459) );
  INV_X1 round_inst_S_6__sbox_inst_com_z_inst_U14 ( .A(round_inst_sin_w[25]), 
        .ZN(round_inst_S_6__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U13 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n393), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U12 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n391), .A2(round_inst_n49), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U11 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_6__sbox_inst_com_z_inst_n390), .Z(
        round_inst_S_6__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U10 ( .A1(round_inst_sin_w[25]), .A2(round_inst_sin_y[27]), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n390) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U9 ( .A1(round_inst_n64), .A2(
        round_inst_sin_w[27]), .ZN(round_inst_S_6__sbox_inst_com_z_inst_n418)
         );
  NOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U8 ( .A1(
        round_inst_S_6__sbox_inst_com_z_inst_n439), .A2(
        round_inst_S_6__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_6__sbox_inst_com_z_inst_U7 ( .A1(round_inst_sin_w[26]), 
        .A2(round_inst_sin_w[25]), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n456) );
  XNOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U6 ( .A(round_inst_sin_x[27]), 
        .B(round_inst_sin_y[27]), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n439) );
  NAND3_X1 round_inst_S_6__sbox_inst_com_z_inst_U5 ( .A1(round_inst_sin_w[26]), 
        .A2(round_inst_sin_x[27]), .A3(
        round_inst_S_6__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U4 ( .A(round_inst_n64), .B(
        round_inst_sin_y[25]), .Z(round_inst_S_6__sbox_inst_com_z_inst_n475)
         );
  INV_X1 round_inst_S_6__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_6__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_6__sbox_inst_com_z_inst_n496) );
  INV_X1 round_inst_S_6__sbox_inst_com_z_inst_U2 ( .A(round_inst_sin_w[24]), 
        .ZN(round_inst_S_6__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_6__sbox_inst_com_z_inst_U1 ( .A(round_inst_n47), .B(
        round_inst_sin_x[22]), .Z(round_inst_S_6__sbox_inst_com_z_inst_n417)
         );
  INV_X1 round_inst_S_7__sbox_inst_U6 ( .A(round_inst_sin_x[30]), .ZN(
        round_inst_S_7__sbox_inst_n6) );
  INV_X1 round_inst_S_7__sbox_inst_U5 ( .A(round_inst_sin_z[29]), .ZN(
        round_inst_S_7__sbox_inst_n2) );
  INV_X1 round_inst_S_7__sbox_inst_U4 ( .A(round_inst_sin_z[31]), .ZN(
        round_inst_S_7__sbox_inst_n4) );
  INV_X2 round_inst_S_7__sbox_inst_U3 ( .A(round_inst_S_7__sbox_inst_n4), .ZN(
        round_inst_S_7__sbox_inst_n3) );
  INV_X2 round_inst_S_7__sbox_inst_U2 ( .A(round_inst_S_7__sbox_inst_n2), .ZN(
        round_inst_S_7__sbox_inst_n1) );
  INV_X2 round_inst_S_7__sbox_inst_U1 ( .A(round_inst_S_7__sbox_inst_n6), .ZN(
        round_inst_S_7__sbox_inst_n5) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n531), .ZN(round_inst_sout_w[31])
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U139 ( .A1(
        round_inst_sin_z[28]), .A2(round_inst_S_7__sbox_inst_com_w_inst_n528), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n526), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n524), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n526) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[30]), .A2(round_inst_S_7__sbox_inst_com_w_inst_n523), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n525) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n518), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n516), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n518) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n514), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n513), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n512), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n513) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_w_inst_U128 ( .A1(
        round_inst_S_7__sbox_inst_n5), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n510), .A3(
        round_inst_S_7__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n511) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U127 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n508), .A2(round_inst_n50), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n507), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U125 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n507) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_7__sbox_inst_n3), .A2(round_inst_n51), .A3(
        round_inst_S_7__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U122 ( .A(round_inst_sin_y[27]), .B(round_inst_S_7__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U121 ( .A(round_inst_n65), .B(
        round_inst_sin_z[27]), .Z(round_inst_S_7__sbox_inst_com_w_inst_n501)
         );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U120 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[29])
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[25]), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[25]), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U113 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[28])
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_7__sbox_inst_n5), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U110 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n528), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U105 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_7__sbox_inst_n5), .B(round_inst_sin_z[30]), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_7__sbox_inst_n1), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U99 ( .A1(round_inst_n51), 
        .A2(round_inst_S_7__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_7__sbox_inst_n5), .A2(round_inst_n50), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n506) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U94 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[30]), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n461), .A2(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[30]), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U88 ( .A1(round_inst_sin_z[28]), 
        .A2(round_inst_S_7__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_w_inst_U85 ( .A1(round_inst_sin_y[29]), .A2(round_inst_n50), .A3(round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_w_inst_U84 ( .A1(round_inst_n51), 
        .A2(round_inst_n65), .A3(round_inst_n50), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n528) );
  OR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_7__sbox_inst_n5), .B(round_inst_n51), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U80 ( .A(round_inst_n48), .B(
        round_inst_sin_z[24]), .Z(round_inst_S_7__sbox_inst_com_w_inst_n484)
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U79 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[31])
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U73 ( .A1(
        round_inst_S_7__sbox_inst_n3), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U71 ( .A1(round_inst_n51), 
        .A2(round_inst_n65), .ZN(round_inst_S_7__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_7__sbox_inst_n5), .A2(round_inst_sin_y[29]), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U69 ( .A1(
        round_inst_S_7__sbox_inst_n1), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n508), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_7__sbox_inst_n5), .A2(round_inst_S_7__sbox_inst_n1), .A3(
        round_inst_S_7__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n439), .A2(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n508), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_7__sbox_inst_n3), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n504) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U62 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n508) );
  INV_X1 round_inst_S_7__sbox_inst_com_w_inst_U61 ( .A(round_inst_n51), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U60 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U58 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U57 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U56 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U55 ( .A(round_inst_sin_y[29]), 
        .B(round_inst_S_7__sbox_inst_n1), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U54 ( .A1(
        round_inst_S_7__sbox_inst_n3), .A2(round_inst_S_7__sbox_inst_n1), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U52 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_w_inst_U51 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n505), .A3(
        round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U50 ( .A(round_inst_sin_y[29]), 
        .B(round_inst_n65), .Z(round_inst_S_7__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_w_inst_U49 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n505), .A2(round_inst_sin_y[29]), 
        .A3(round_inst_S_7__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U48 ( .A(round_inst_n51), .B(
        round_inst_sin_z[30]), .ZN(round_inst_S_7__sbox_inst_com_w_inst_n465)
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U47 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n520) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U45 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n421), .A2(
        round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U44 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U43 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n419), .A2(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U42 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U40 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_7__sbox_inst_n1), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n521) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U38 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U37 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U36 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n510), .B(round_inst_sin_z[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n498), .A2(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U33 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U32 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U31 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U30 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U29 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U28 ( .A1(round_inst_n65), 
        .A2(round_inst_sin_z[28]), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U27 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n522), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U26 ( .A(round_inst_n65), .B(
        round_inst_S_7__sbox_inst_n1), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U24 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n510), .A2(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U22 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[29]), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U21 ( .A(round_inst_n50), .B(
        round_inst_sin_z[28]), .Z(round_inst_S_7__sbox_inst_com_w_inst_n418)
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U20 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U19 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U17 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n398), .A2(
        round_inst_S_7__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U15 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n498), .B(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_7__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_7__sbox_inst_com_w_inst_U13 ( .A(round_inst_sin_y[31]), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_7__sbox_inst_n1), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U11 ( .A(
        round_inst_S_7__sbox_inst_n3), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n505), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U9 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_7__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_7__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U8 ( .A1(round_inst_n65), .A2(
        round_inst_n50), .ZN(round_inst_S_7__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U7 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n510), .A2(round_inst_sin_y[29]), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n477) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_w_inst_U6 ( .A1(
        round_inst_S_7__sbox_inst_com_w_inst_n505), .A2(round_inst_n50), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n522) );
  INV_X1 round_inst_S_7__sbox_inst_com_w_inst_U5 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n505) );
  INV_X1 round_inst_S_7__sbox_inst_com_w_inst_U4 ( .A(round_inst_sin_x[31]), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n486) );
  INV_X1 round_inst_S_7__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_7__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_7__sbox_inst_com_w_inst_n510) );
  INV_X1 round_inst_S_7__sbox_inst_com_w_inst_U2 ( .A(round_inst_sin_x[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_w_inst_n489) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_w_inst_U1 ( .A(round_inst_n49), .B(
        round_inst_sin_z[26]), .Z(round_inst_S_7__sbox_inst_com_w_inst_n402)
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n510), .ZN(round_inst_sout_x[28])
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n509), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n510) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U133 ( .A(round_inst_n51), .B(
        round_inst_sin_y[31]), .ZN(round_inst_S_7__sbox_inst_com_x_inst_n508)
         );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U132 ( .A(round_inst_sin_z[24]), 
        .B(round_inst_S_7__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n506), .Z(round_inst_srout2_x[30]) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U130 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U129 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n503), .A2(round_inst_sin_z[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U127 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U126 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U125 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U124 ( .A1(round_inst_n51), 
        .A2(round_inst_sin_w[28]), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U122 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U121 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U118 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_sin_y[31]), .A2(round_inst_S_7__sbox_inst_com_x_inst_n490), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U115 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n487) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_x_inst_U114 ( .A1(
        round_inst_sin_z[30]), .A2(round_inst_sin_w[28]), .A3(
        round_inst_sin_y[31]), .ZN(round_inst_S_7__sbox_inst_com_x_inst_n489)
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n478), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n476), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n478) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n475), .B(round_inst_sin_z[27]), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n476) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_w[30]), .A2(round_inst_sin_y[31]), .A3(
        round_inst_sin_z[28]), .ZN(round_inst_S_7__sbox_inst_com_x_inst_n475)
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n474), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n473), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n473) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n470), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n469), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n511) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n468), .A2(round_inst_n51), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n469) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n468) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n467), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n464), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_srout2_x[28]) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U100 ( .A1(round_inst_n50), 
        .A2(round_inst_sin_z[30]), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[25]), 
        .B(round_inst_S_7__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n464) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n462), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n460), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n467), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n461) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n458), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n467) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_7__sbox_inst_n1), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n457), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n459) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n455), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n454), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n456) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n453), .A2(round_inst_sin_w[30]), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n454) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n451), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n455) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n450), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n449), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n451) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n448), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n447), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n449) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n446), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_7__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n445), .B(round_inst_n51), .S(
        round_inst_n50), .Z(round_inst_S_7__sbox_inst_com_x_inst_n446) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n444), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n448) );
  MUX2_X1 round_inst_S_7__sbox_inst_com_x_inst_U85 ( .A(round_inst_n51), .B(
        round_inst_sin_z[30]), .S(round_inst_sin_z[28]), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n443), .A2(round_inst_sin_w[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n442), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n441), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n452) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[28]), 
        .A3(round_inst_sin_z[30]), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n441) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n440), .A2(round_inst_sin_w[29]), 
        .A3(round_inst_n51), .ZN(round_inst_S_7__sbox_inst_com_x_inst_n442) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U80 ( .A(round_inst_n50), .B(
        round_inst_sin_z[28]), .Z(round_inst_S_7__sbox_inst_com_x_inst_n440)
         );
  NAND3_X1 round_inst_S_7__sbox_inst_com_x_inst_U79 ( .A1(round_inst_n50), 
        .A2(round_inst_S_7__sbox_inst_com_x_inst_n445), .A3(
        round_inst_S_7__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n460) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U77 ( .A1(round_inst_n50), 
        .A2(round_inst_n51), .ZN(round_inst_S_7__sbox_inst_com_x_inst_n482) );
  AND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U76 ( .A1(round_inst_n51), .A2(
        round_inst_sin_z[28]), .ZN(round_inst_S_7__sbox_inst_com_x_inst_n490)
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n462) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U74 ( .A1(round_inst_n50), 
        .A2(round_inst_sin_w[30]), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n497) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_srout2_x[31]) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n436), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n435), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U71 ( .A(round_inst_n50), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n435) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n434), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n433), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U69 ( .A1(round_inst_sin_z[28]), .A2(round_inst_sin_y[31]), .ZN(round_inst_S_7__sbox_inst_com_x_inst_n433) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n432), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n431), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n434) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n430), .A2(round_inst_n50), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n431) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n429), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n428), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_7__sbox_inst_n1), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n453), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n432) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[26]), 
        .B(round_inst_S_7__sbox_inst_com_x_inst_n438), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n436) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n425), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n424), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n423), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n422), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n421), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n420), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n422) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n419), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n420) );
  NOR3_X1 round_inst_S_7__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n471), .A3(
        round_inst_S_7__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n418) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n416), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n419) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n414), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U53 ( .A1(round_inst_n51), 
        .A2(round_inst_S_7__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n413) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U52 ( .A(round_inst_sin_y[31]), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n414) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n443), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n416) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U50 ( .A1(
        round_inst_S_7__sbox_inst_n1), .A2(round_inst_n51), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n443) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_x_inst_U49 ( .A1(round_inst_n51), 
        .A2(round_inst_S_7__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_7__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n421) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n411), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n423) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U47 ( .A1(round_inst_n51), 
        .A2(round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n465) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n411) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n410), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n407), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U43 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n406), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n405), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n407) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U42 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n466), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n405) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U41 ( .A(round_inst_sin_w[29]), 
        .B(round_inst_S_7__sbox_inst_n1), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n439) );
  AND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U40 ( .A1(round_inst_sin_z[30]), 
        .A2(round_inst_sin_y[31]), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_7__sbox_inst_n3), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n406) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_x_inst_U38 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U37 ( .A(round_inst_sin_z[30]), 
        .B(round_inst_sin_w[30]), .Z(round_inst_S_7__sbox_inst_com_x_inst_n445) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U36 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n404), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n410) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U35 ( .A(round_inst_sin_w[30]), 
        .B(round_inst_n51), .Z(round_inst_S_7__sbox_inst_com_x_inst_n403) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n402), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n401), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U33 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n400), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n399), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n401) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U32 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n399) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U31 ( .A1(round_inst_sin_z[28]), .A2(round_inst_S_7__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n426) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n427), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n400) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U28 ( .A(round_inst_sin_y[31]), 
        .B(round_inst_S_7__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n471) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n402) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_7__sbox_inst_n1), .A3(round_inst_n50), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n396) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n398), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n481) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U23 ( .A(round_inst_sin_y[31]), 
        .B(round_inst_S_7__sbox_inst_n3), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U21 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n392), .A2(round_inst_sin_w[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n404), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_x_inst_U17 ( .A1(round_inst_sin_z[28]), .A2(round_inst_sin_y[31]), .A3(round_inst_sin_w[29]), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n388) );
  MUX2_X1 round_inst_S_7__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n412), .B(round_inst_sin_y[31]), 
        .S(round_inst_S_7__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U15 ( .A1(round_inst_n50), 
        .A2(round_inst_S_7__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U14 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n491), .B(
        round_inst_S_7__sbox_inst_n3), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n412) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n384), .A2(round_inst_sin_z[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U10 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_7__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U9 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_w[31]), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U7 ( .A1(
        round_inst_S_7__sbox_inst_n1), .A2(round_inst_sin_y[31]), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n404) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_7__sbox_inst_com_x_inst_n427), .Z(
        round_inst_S_7__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U4 ( .A1(round_inst_n50), .A2(
        round_inst_sin_w[29]), .ZN(round_inst_S_7__sbox_inst_com_x_inst_n427)
         );
  NAND2_X1 round_inst_S_7__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_7__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_7__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_7__sbox_inst_com_x_inst_n477) );
  INV_X1 round_inst_S_7__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_y[29]), 
        .ZN(round_inst_S_7__sbox_inst_com_x_inst_n417) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n517), .Z(round_inst_sout_y[28])
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n516), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n515) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U134 ( .A(round_inst_sin_x[24]), 
        .B(round_inst_S_7__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n512), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_srout2_y[30]) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n508), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n518) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n507), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n506), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n508) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n506) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n507) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_7__sbox_inst_com_y_inst_U125 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_7__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U124 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U123 ( .A1(
        round_inst_sin_x[31]), .A2(round_inst_S_7__sbox_inst_com_y_inst_n493), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n492), .A2(
        round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U121 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U120 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U119 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U118 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n486), .A2(
        round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U117 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n503), .A2(round_inst_sin_w[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U112 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_7__sbox_inst_n1), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[27]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_y_inst_U109 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_7__sbox_inst_n3), .A3(round_inst_sin_x[28]), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U108 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_y_inst_U107 ( .A1(
        round_inst_sin_w[28]), .A2(round_inst_sin_w[31]), .A3(
        round_inst_S_7__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_7__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_7__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U105 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[28]) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U104 ( .A1(
        round_inst_S_7__sbox_inst_n5), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U98 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_7__sbox_inst_n1), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U95 ( .A1(round_inst_sin_x[28]), .A2(round_inst_S_7__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_y_inst_U94 ( .A1(round_inst_sin_w[28]), .A2(round_inst_n65), .A3(round_inst_S_7__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U93 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U92 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U88 ( .A1(
        round_inst_S_7__sbox_inst_n1), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_7__sbox_inst_com_y_inst_U87 ( .A(
        round_inst_S_7__sbox_inst_n5), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n503), .S(
        round_inst_S_7__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_7__sbox_inst_n1), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n478), .B(round_inst_n64), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n438), .Z(round_inst_srout2_y[31]) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U71 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[31]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U70 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n483), .A2(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_7__sbox_inst_n1), .A2(round_inst_sin_w[28]), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[31]), 
        .A3(round_inst_S_7__sbox_inst_n1), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U66 ( .A(round_inst_sin_w[28]), 
        .B(round_inst_sin_x[28]), .Z(round_inst_S_7__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U59 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[31]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U58 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[29]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U55 ( .A(round_inst_sin_x[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U54 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n418), .A2(
        round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U53 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U51 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U50 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n414), .B(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U49 ( .A(round_inst_sin_w[29]), 
        .B(round_inst_S_7__sbox_inst_n1), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U48 ( .A1(
        round_inst_S_7__sbox_inst_n1), .A2(round_inst_sin_x[28]), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_7__sbox_inst_n1), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U46 ( .A(round_inst_sin_x[26]), 
        .B(round_inst_S_7__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n513) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[29]), 
        .B(round_inst_sin_x[31]), .Z(round_inst_S_7__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U41 ( .A(round_inst_n65), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[31]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[28]), 
        .Z(round_inst_S_7__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U36 ( .A(round_inst_sin_z[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_7__sbox_inst_n1), .B(round_inst_S_7__sbox_inst_n3), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_7__sbox_inst_n5), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U27 ( .A1(round_inst_sin_w[29]), .A2(round_inst_S_7__sbox_inst_n3), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n514), .A2(round_inst_sin_w[29]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_7__sbox_inst_n1), .A2(round_inst_sin_w[31]), .A3(
        round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_7__sbox_inst_n1), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n504), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_7__sbox_inst_n3), .B(round_inst_sin_w[31]), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U17 ( .A(
        round_inst_S_7__sbox_inst_n3), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[31]), 
        .B(round_inst_sin_x[31]), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_y_inst_U13 ( .A1(round_inst_n65), 
        .A2(round_inst_sin_w[31]), .A3(
        round_inst_S_7__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_y_inst_U12 ( .A1(
        round_inst_S_7__sbox_inst_n3), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_7__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[29]), 
        .B(round_inst_n65), .S(round_inst_S_7__sbox_inst_com_y_inst_n503), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_y_inst_U9 ( .A1(round_inst_n65), .A2(
        round_inst_S_7__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_7__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_7__sbox_inst_n3), .B(round_inst_sin_x[31]), .Z(
        round_inst_S_7__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_7__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_7__sbox_inst_n1), .A3(round_inst_sin_x[31]), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_7__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n503) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[30]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_7__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_7__sbox_inst_com_y_inst_n514) );
  INV_X1 round_inst_S_7__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[30]), 
        .ZN(round_inst_S_7__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n516), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n515), .ZN(round_inst_sout_z[28])
         );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n514), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n513), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_w[30]), .B(round_inst_sin_w[31]), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n513) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U128 ( .A(round_inst_sin_x[24]), 
        .B(round_inst_n48), .Z(round_inst_S_7__sbox_inst_com_z_inst_n514) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n510), .ZN(
        round_inst_srout2_z[30]) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n509), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n508), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U124 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n507), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n506), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n508) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U123 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n505), .A2(round_inst_n50), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n506) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n504), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n503), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n502), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n501), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n503) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U120 ( .A(round_inst_sin_w[29]), .B(round_inst_sin_x[27]), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n501) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U119 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n500), .B(round_inst_sin_y[27]), 
        .Z(round_inst_S_7__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U118 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n499), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n498), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n500) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U117 ( .A1(round_inst_n51), 
        .A2(round_inst_S_7__sbox_inst_com_z_inst_n497), .A3(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n498) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U116 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n495), .A2(round_inst_sin_x[28]), 
        .A3(round_inst_sin_w[31]), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n499) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U115 ( .A(
        round_inst_S_7__sbox_inst_n5), .B(round_inst_n51), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n495) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U114 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_7__sbox_inst_n5), .A3(round_inst_sin_x[31]), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n509) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n491), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n493) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U111 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n490), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n489), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n491) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n488), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n486), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n490) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U108 ( .A1(
        round_inst_sin_w[30]), .A2(round_inst_sin_x[31]), .A3(round_inst_n50), 
        .ZN(round_inst_S_7__sbox_inst_com_z_inst_n492) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U107 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n484), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U106 ( .A1(
        round_inst_sin_w[30]), .A2(round_inst_S_7__sbox_inst_com_z_inst_n497), 
        .ZN(round_inst_S_7__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n505), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n484) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n482), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n481), .Z(round_inst_srout2_z[28]) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n479), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n478), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n483), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U101 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n483) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U100 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n475), .A2(round_inst_sin_x[28]), 
        .A3(round_inst_sin_w[30]), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U99 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n474), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n477) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U98 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n472), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .A3(round_inst_n51), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n473) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U97 ( .A(round_inst_sin_w[29]), 
        .B(round_inst_sin_y[29]), .Z(round_inst_S_7__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U96 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n471), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n474) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U95 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n469), .A2(
        round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n470) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n467), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n471) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n466), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n465), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n464), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n463), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U91 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n462), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n461), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U90 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n460), .A2(round_inst_n51), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n461) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U89 ( .A1(round_inst_n65), 
        .A2(round_inst_S_7__sbox_inst_n5), .A3(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n462) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n459), .A2(round_inst_n50), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U87 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_w[30]), 
        .ZN(round_inst_S_7__sbox_inst_com_z_inst_n466) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U85 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U84 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n453), .A2(round_inst_n51), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n454) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U83 ( .A(round_inst_sin_w[29]), 
        .B(round_inst_S_7__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n451), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U81 ( .A1(round_inst_sin_w[30]), .A2(round_inst_sin_x[28]), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n478) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U79 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n487), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n448) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U78 ( .A(round_inst_sin_y[25]), 
        .B(round_inst_n64), .Z(round_inst_S_7__sbox_inst_com_z_inst_n447) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n487) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U76 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n446), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U75 ( .A(round_inst_sin_w[30]), 
        .B(round_inst_n51), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_srout2_z[31]) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n511), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U72 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n511) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U71 ( .A1(round_inst_sin_x[28]), .A2(round_inst_sin_w[31]), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n441) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U70 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n458), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n440), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n442) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U69 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U68 ( .A(round_inst_sin_w[31]), 
        .B(round_inst_S_7__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n497) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n494) );
  MUX2_X1 round_inst_S_7__sbox_inst_com_z_inst_U66 ( .A(round_inst_sin_x[31]), 
        .B(round_inst_sin_w[31]), .S(round_inst_S_7__sbox_inst_com_z_inst_n436), .Z(round_inst_S_7__sbox_inst_com_z_inst_n437) );
  OR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U65 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n436) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U64 ( .A(round_inst_sin_x[28]), 
        .B(round_inst_S_7__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n486) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U63 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n438) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U62 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_x[31]), 
        .A3(round_inst_S_7__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n430), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U59 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n429) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U58 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n426), .A2(round_inst_sin_w[31]), 
        .ZN(round_inst_S_7__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U56 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n422), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n424) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U55 ( .A1(round_inst_sin_x[28]), .A2(round_inst_n65), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U54 ( .A1(round_inst_sin_y[29]), .A2(round_inst_sin_x[28]), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n425) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U53 ( .A1(round_inst_n50), 
        .A2(round_inst_sin_x[31]), .A3(round_inst_sin_w[29]), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n428) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U52 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_y[31]), 
        .ZN(round_inst_S_7__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U50 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n460), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n423), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n469) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U49 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_y[29]), 
        .ZN(round_inst_S_7__sbox_inst_com_z_inst_n423) );
  AND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U48 ( .A1(round_inst_sin_w[29]), 
        .A2(round_inst_sin_x[28]), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n460) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U47 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n421) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U46 ( .A1(round_inst_sin_w[29]), .A2(round_inst_S_7__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .A2(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U44 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n419), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n418), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n432) );
  INV_X1 round_inst_S_7__sbox_inst_com_z_inst_U43 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .B(round_inst_n50), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n451) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U41 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n417), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n496), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U39 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n449) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U38 ( .A1(round_inst_sin_w[31]), .A2(round_inst_S_7__sbox_inst_com_z_inst_n413), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n414) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n415) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U35 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U34 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n505), .A2(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n409) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U32 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n407) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n405) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U30 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n404) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n505), .A2(round_inst_sin_y[29]), 
        .ZN(round_inst_S_7__sbox_inst_com_z_inst_n402) );
  AND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_S_7__sbox_inst_n5), .A2(round_inst_sin_w[31]), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n505) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U27 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n401), .A2(round_inst_n51), .A3(
        round_inst_sin_w[29]), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n403)
         );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U26 ( .A(round_inst_sin_w[31]), 
        .B(round_inst_sin_x[31]), .Z(round_inst_S_7__sbox_inst_com_z_inst_n401) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U25 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n399), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n406) );
  MUX2_X1 round_inst_S_7__sbox_inst_com_z_inst_U24 ( .A(round_inst_sin_y[31]), 
        .B(round_inst_S_7__sbox_inst_com_z_inst_n398), .S(
        round_inst_S_7__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U23 ( .A1(round_inst_sin_w[29]), .A2(round_inst_S_7__sbox_inst_n5), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n398) );
  INV_X1 round_inst_S_7__sbox_inst_com_z_inst_U21 ( .A(round_inst_sin_x[31]), 
        .ZN(round_inst_S_7__sbox_inst_com_z_inst_n397) );
  NOR3_X1 round_inst_S_7__sbox_inst_com_z_inst_U20 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n488), .A3(
        round_inst_S_7__sbox_inst_com_z_inst_n395), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U19 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n394), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n395) );
  INV_X1 round_inst_S_7__sbox_inst_com_z_inst_U18 ( .A(round_inst_n65), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n394) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U17 ( .A(round_inst_sin_w[31]), 
        .B(round_inst_sin_y[31]), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n488) );
  AND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U16 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n459), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U15 ( .A1(round_inst_sin_w[30]), .A2(round_inst_n65), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n459) );
  INV_X1 round_inst_S_7__sbox_inst_com_z_inst_U14 ( .A(round_inst_sin_w[29]), 
        .ZN(round_inst_S_7__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U13 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n393), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U12 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n391), .A2(round_inst_n51), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U11 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_7__sbox_inst_com_z_inst_n390), .Z(
        round_inst_S_7__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U10 ( .A1(round_inst_sin_w[29]), .A2(round_inst_sin_y[31]), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n390) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U9 ( .A1(round_inst_n65), .A2(
        round_inst_sin_w[31]), .ZN(round_inst_S_7__sbox_inst_com_z_inst_n418)
         );
  NOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U8 ( .A1(
        round_inst_S_7__sbox_inst_com_z_inst_n439), .A2(
        round_inst_S_7__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_7__sbox_inst_com_z_inst_U7 ( .A1(round_inst_sin_w[30]), 
        .A2(round_inst_sin_w[29]), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n456) );
  XNOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U6 ( .A(round_inst_sin_x[31]), 
        .B(round_inst_sin_y[31]), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n439) );
  NAND3_X1 round_inst_S_7__sbox_inst_com_z_inst_U5 ( .A1(round_inst_sin_w[30]), 
        .A2(round_inst_sin_x[31]), .A3(
        round_inst_S_7__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U4 ( .A(round_inst_n65), .B(
        round_inst_sin_y[29]), .Z(round_inst_S_7__sbox_inst_com_z_inst_n475)
         );
  INV_X1 round_inst_S_7__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_7__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_7__sbox_inst_com_z_inst_n496) );
  INV_X1 round_inst_S_7__sbox_inst_com_z_inst_U2 ( .A(round_inst_sin_w[28]), 
        .ZN(round_inst_S_7__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_7__sbox_inst_com_z_inst_U1 ( .A(round_inst_n49), .B(
        round_inst_sin_x[26]), .Z(round_inst_S_7__sbox_inst_com_z_inst_n417)
         );
  INV_X1 round_inst_S_8__sbox_inst_U6 ( .A(round_inst_sin_x[34]), .ZN(
        round_inst_S_8__sbox_inst_n6) );
  INV_X1 round_inst_S_8__sbox_inst_U5 ( .A(round_inst_sin_z[33]), .ZN(
        round_inst_S_8__sbox_inst_n2) );
  INV_X1 round_inst_S_8__sbox_inst_U4 ( .A(round_inst_sin_z[35]), .ZN(
        round_inst_S_8__sbox_inst_n4) );
  INV_X2 round_inst_S_8__sbox_inst_U3 ( .A(round_inst_S_8__sbox_inst_n4), .ZN(
        round_inst_S_8__sbox_inst_n3) );
  INV_X2 round_inst_S_8__sbox_inst_U2 ( .A(round_inst_S_8__sbox_inst_n2), .ZN(
        round_inst_S_8__sbox_inst_n1) );
  INV_X2 round_inst_S_8__sbox_inst_U1 ( .A(round_inst_S_8__sbox_inst_n6), .ZN(
        round_inst_S_8__sbox_inst_n5) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n529), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n528), .ZN(round_inst_sout_w[35])
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n526), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n528) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[32]), .A2(round_inst_S_8__sbox_inst_com_w_inst_n525), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n526) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n524), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n523), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n523) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U133 ( .A1(
        round_inst_sin_z[34]), .A2(round_inst_S_8__sbox_inst_com_w_inst_n520), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n521) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U132 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n519), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n518), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n520) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n517), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n516), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n522) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n515), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n514), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n516) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U129 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n518), .A2(
        round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U128 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n513), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n512), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U127 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n511), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n512) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U126 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n508), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n510) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_w_inst_U125 ( .A1(
        round_inst_S_8__sbox_inst_n5), .A2(round_inst_sin_x[32]), .A3(
        round_inst_S_8__sbox_inst_com_w_inst_n507), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n508) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n506), .A2(round_inst_n52), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n509) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U123 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n505), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n511) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U122 ( .A(round_inst_sin_x[35]), .B(round_inst_S_8__sbox_inst_com_w_inst_n503), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n505) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_w_inst_U121 ( .A1(
        round_inst_S_8__sbox_inst_n3), .A2(round_inst_n53), .A3(
        round_inst_sin_x[32]), .ZN(round_inst_S_8__sbox_inst_com_w_inst_n513)
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U120 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n502), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U119 ( .A(round_inst_sin_y[31]), .B(round_inst_S_8__sbox_inst_com_w_inst_n500), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n501) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U118 ( .A(round_inst_n66), .B(
        round_inst_sin_z[31]), .Z(round_inst_S_8__sbox_inst_com_w_inst_n500)
         );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U117 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n499), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n502) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U116 ( .A(round_inst_sin_x[35]), .B(round_inst_sin_y[35]), .ZN(round_inst_S_8__sbox_inst_com_w_inst_n499) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[33])
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U113 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[29]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[29]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U110 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[32])
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_8__sbox_inst_n5), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n529), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U105 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n529) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U104 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U102 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_8__sbox_inst_n5), .B(round_inst_sin_z[34]), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U99 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_8__sbox_inst_n1), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n504), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U96 ( .A1(round_inst_n53), 
        .A2(round_inst_sin_x[32]), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n498) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U95 ( .A1(
        round_inst_S_8__sbox_inst_n5), .A2(round_inst_n52), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n504) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U94 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U93 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[34]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U90 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U89 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U88 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n461), .A2(round_inst_n66), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[34]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U86 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U85 ( .A1(round_inst_sin_z[32]), 
        .A2(round_inst_S_8__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U84 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_w_inst_U82 ( .A1(round_inst_sin_y[33]), .A2(round_inst_n52), .A3(round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_w_inst_U81 ( .A1(round_inst_n53), 
        .A2(round_inst_n66), .A3(round_inst_n52), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U80 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n525) );
  OR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U79 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_8__sbox_inst_n5), .B(round_inst_n53), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U77 ( .A(round_inst_n50), .B(
        round_inst_sin_z[28]), .Z(round_inst_S_8__sbox_inst_com_w_inst_n484)
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[35])
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U73 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U71 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_8__sbox_inst_n3), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U69 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U68 ( .A1(round_inst_n53), 
        .A2(round_inst_n66), .ZN(round_inst_S_8__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_8__sbox_inst_n5), .A2(round_inst_sin_y[33]), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U66 ( .A1(
        round_inst_S_8__sbox_inst_n1), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_w_inst_U65 ( .A1(
        round_inst_S_8__sbox_inst_n5), .A2(round_inst_S_8__sbox_inst_n1), .A3(
        round_inst_sin_x[35]), .ZN(round_inst_S_8__sbox_inst_com_w_inst_n444)
         );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n439), .A2(round_inst_n66), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U62 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U61 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n503), .A2(
        round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U60 ( .A(
        round_inst_S_8__sbox_inst_n3), .B(round_inst_sin_y[35]), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n503) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n506) );
  INV_X1 round_inst_S_8__sbox_inst_com_w_inst_U58 ( .A(round_inst_sin_x[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n486) );
  INV_X1 round_inst_S_8__sbox_inst_com_w_inst_U57 ( .A(round_inst_n53), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U56 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U55 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U54 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U52 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U51 ( .A(round_inst_sin_y[33]), 
        .B(round_inst_S_8__sbox_inst_n1), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U50 ( .A1(
        round_inst_S_8__sbox_inst_n3), .A2(round_inst_S_8__sbox_inst_n1), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U49 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U48 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_w_inst_U47 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n425), .A2(round_inst_sin_x[35]), 
        .A3(round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U46 ( .A(round_inst_sin_y[33]), 
        .B(round_inst_n66), .Z(round_inst_S_8__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_w_inst_U45 ( .A1(round_inst_sin_x[35]), .A2(round_inst_sin_y[33]), .A3(round_inst_S_8__sbox_inst_com_w_inst_n465), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U44 ( .A(round_inst_n53), .B(
        round_inst_sin_z[34]), .ZN(round_inst_S_8__sbox_inst_com_w_inst_n465)
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U43 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U42 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n517) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U41 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n421), .A2(
        round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U40 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n419), .A2(round_inst_n66), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U38 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U37 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U36 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n518), .A2(
        round_inst_S_8__sbox_inst_n1), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U35 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n518) );
  INV_X1 round_inst_S_8__sbox_inst_com_w_inst_U34 ( .A(round_inst_sin_x[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n489) );
  INV_X1 round_inst_S_8__sbox_inst_com_w_inst_U33 ( .A(round_inst_sin_y[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n434) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U32 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U31 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U30 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U29 ( .A(round_inst_sin_x[32]), 
        .B(round_inst_sin_z[32]), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U28 ( .A1(round_inst_sin_y[35]), .A2(round_inst_n66), .ZN(round_inst_S_8__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U27 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U26 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n407), .A2(round_inst_sin_y[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U24 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_x[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U23 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U22 ( .A1(round_inst_n66), 
        .A2(round_inst_sin_z[32]), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U21 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_8__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U20 ( .A(round_inst_n66), .B(
        round_inst_S_8__sbox_inst_n1), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U19 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n404), .A2(round_inst_sin_x[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U17 ( .A1(round_inst_sin_x[32]), .A2(round_inst_n66), .ZN(round_inst_S_8__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U16 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[33]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U15 ( .A(round_inst_n52), .B(
        round_inst_sin_z[32]), .Z(round_inst_S_8__sbox_inst_com_w_inst_n418)
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U13 ( .A(round_inst_sin_x[32]), 
        .B(round_inst_S_8__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U11 ( .A1(
        round_inst_S_8__sbox_inst_com_w_inst_n398), .A2(round_inst_sin_x[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U9 ( .A(round_inst_sin_y[35]), 
        .B(round_inst_n66), .ZN(round_inst_S_8__sbox_inst_com_w_inst_n396) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U8 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_8__sbox_inst_n1), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U7 ( .A(
        round_inst_S_8__sbox_inst_n3), .B(round_inst_sin_x[35]), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n507) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U6 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n519), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U5 ( .A(
        round_inst_S_8__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_8__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_8__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U4 ( .A1(round_inst_n66), .A2(
        round_inst_n52), .ZN(round_inst_S_8__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U3 ( .A1(round_inst_sin_x[32]), 
        .A2(round_inst_sin_y[33]), .ZN(
        round_inst_S_8__sbox_inst_com_w_inst_n477) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_w_inst_U2 ( .A1(round_inst_sin_x[35]), 
        .A2(round_inst_n52), .ZN(round_inst_S_8__sbox_inst_com_w_inst_n519) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_w_inst_U1 ( .A(round_inst_n51), .B(
        round_inst_sin_z[30]), .Z(round_inst_S_8__sbox_inst_com_w_inst_n402)
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U136 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n512), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n511), .ZN(round_inst_sout_x[32])
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n510), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n509), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n511) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U134 ( .A(round_inst_n53), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U133 ( .A(round_inst_sin_z[28]), 
        .B(round_inst_S_8__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n510) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U132 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n512), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n506), .Z(round_inst_srout2_x[50]) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U130 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n503), .A2(round_inst_sin_z[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U129 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U127 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U126 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U125 ( .A1(round_inst_n53), 
        .A2(round_inst_sin_w[32]), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U124 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U122 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U121 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U118 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n508), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n487) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U115 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n481) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_x_inst_U114 ( .A1(
        round_inst_sin_z[34]), .A2(round_inst_sin_w[32]), .A3(
        round_inst_S_8__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n489) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n478), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n475), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n477) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n474), .B(round_inst_sin_z[31]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n475) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_w[34]), .A2(round_inst_S_8__sbox_inst_com_x_inst_n508), 
        .A3(round_inst_sin_z[32]), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n473), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n478) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n470), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n473) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n468), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n512) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n467), .A2(round_inst_n53), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n468) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n467) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n469) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n465), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n463), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_srout2_x[48]) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U100 ( .A1(round_inst_n52), 
        .A2(round_inst_sin_z[34]), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[29]), 
        .B(round_inst_S_8__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n461), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n462) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n466), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n460) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n458), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n457), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_8__sbox_inst_n1), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n459), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n456), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n455), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n454), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n453), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n455) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n452), .A2(round_inst_sin_w[34]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n451), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n450), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n454) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n449), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n448), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n447), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n446), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n448) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n445), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n446) );
  MUX2_X1 round_inst_S_8__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n444), .B(round_inst_n53), .S(
        round_inst_n52), .Z(round_inst_S_8__sbox_inst_com_x_inst_n445) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n443), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_8__sbox_inst_com_x_inst_U85 ( .A(round_inst_n53), .B(
        round_inst_sin_z[34]), .S(round_inst_sin_z[32]), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n443) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n442), .A2(round_inst_sin_w[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n449) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n441), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n440), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n451) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_w[32]), 
        .A3(round_inst_sin_z[34]), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n440) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n439), .A2(round_inst_sin_w[33]), 
        .A3(round_inst_n53), .ZN(round_inst_S_8__sbox_inst_com_x_inst_n441) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U80 ( .A(round_inst_n52), .B(
        round_inst_sin_z[32]), .Z(round_inst_S_8__sbox_inst_com_x_inst_n439)
         );
  NAND3_X1 round_inst_S_8__sbox_inst_com_x_inst_U79 ( .A1(round_inst_n52), 
        .A2(round_inst_S_8__sbox_inst_com_x_inst_n444), .A3(
        round_inst_S_8__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n456) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n459) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U77 ( .A1(round_inst_n52), 
        .A2(round_inst_n53), .ZN(round_inst_S_8__sbox_inst_com_x_inst_n482) );
  AND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U76 ( .A1(round_inst_n53), .A2(
        round_inst_sin_z[32]), .ZN(round_inst_S_8__sbox_inst_com_x_inst_n490)
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n461) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U74 ( .A1(round_inst_n52), 
        .A2(round_inst_sin_w[34]), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n497) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n436), .ZN(
        round_inst_srout2_x[51]) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n435), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n434), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n436) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U71 ( .A(round_inst_n52), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n434) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n433), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n432), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U69 ( .A1(round_inst_sin_z[32]), .A2(round_inst_S_8__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n432) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n431), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n430), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n433) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n429), .A2(round_inst_n52), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n428), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n427) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_8__sbox_inst_n1), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n431) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n452) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[30]), 
        .B(round_inst_S_8__sbox_inst_com_x_inst_n437), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n435) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n424), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n423), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n422), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n421), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n423) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n420), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n419), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n421) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n418), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n419) );
  NOR3_X1 round_inst_S_8__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n470), .A3(
        round_inst_S_8__sbox_inst_com_x_inst_n416), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n417) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n415), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n414), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n418) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n413), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n414) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U53 ( .A1(round_inst_n53), 
        .A2(round_inst_S_8__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n412) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U52 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n442), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_8__sbox_inst_n1), .A2(round_inst_n53), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n442) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_x_inst_U50 ( .A1(round_inst_n53), 
        .A2(round_inst_S_8__sbox_inst_com_x_inst_n476), .A3(
        round_inst_S_8__sbox_inst_com_x_inst_n411), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n420) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U49 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n410), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n422) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U48 ( .A1(round_inst_n53), 
        .A2(round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n464) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U47 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n410) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n409), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n407), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n406), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n405), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n404), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n406) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U43 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n465), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n404) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U42 ( .A(round_inst_sin_w[33]), 
        .B(round_inst_S_8__sbox_inst_n1), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n438) );
  AND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U41 ( .A1(round_inst_sin_z[34]), 
        .A2(round_inst_S_8__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n465) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U40 ( .A1(
        round_inst_S_8__sbox_inst_n3), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n405) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n476), .A3(
        round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n407) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U38 ( .A(round_inst_sin_z[34]), 
        .B(round_inst_sin_w[34]), .Z(round_inst_S_8__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U37 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n403), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n402), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U36 ( .A(round_inst_sin_w[34]), 
        .B(round_inst_n53), .Z(round_inst_S_8__sbox_inst_com_x_inst_n402) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U35 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n401), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n400), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n399), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n400) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U33 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n398) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U32 ( .A1(round_inst_sin_z[32]), .A2(round_inst_S_8__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n425) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U31 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n479), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n471) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_8__sbox_inst_n3), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n426), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n399) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U28 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n401) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_8__sbox_inst_n1), .A3(round_inst_n52), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n396) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n411), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U23 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n392), .A2(round_inst_sin_w[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U21 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_x_inst_U19 ( .A1(round_inst_sin_z[32]), .A2(round_inst_S_8__sbox_inst_com_x_inst_n508), .A3(round_inst_sin_w[33]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n388) );
  MUX2_X1 round_inst_S_8__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n411), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n508), .S(
        round_inst_S_8__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U17 ( .A1(round_inst_n52), 
        .A2(round_inst_S_8__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n491), .B(
        round_inst_S_8__sbox_inst_n3), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n411) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U15 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U14 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n384), .A2(round_inst_sin_z[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n403), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U10 ( .A(round_inst_sin_w[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U9 ( .A1(
        round_inst_S_8__sbox_inst_n1), .A2(
        round_inst_S_8__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n403) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U8 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n508) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U7 ( .A(round_inst_sin_y[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n413) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_8__sbox_inst_com_x_inst_n426), .Z(
        round_inst_S_8__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U4 ( .A1(round_inst_n52), .A2(
        round_inst_sin_w[33]), .ZN(round_inst_S_8__sbox_inst_com_x_inst_n426)
         );
  NAND2_X1 round_inst_S_8__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_8__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_w[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_8__sbox_inst_com_x_inst_n416), .ZN(
        round_inst_S_8__sbox_inst_com_x_inst_n476) );
  INV_X1 round_inst_S_8__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_y[33]), 
        .ZN(round_inst_S_8__sbox_inst_com_x_inst_n416) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U138 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n519), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n518), .Z(round_inst_sout_y[32])
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n516), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n518) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n515), .B(
        round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n516) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U135 ( .A(round_inst_sin_x[28]), 
        .B(round_inst_S_8__sbox_inst_com_y_inst_n514), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U134 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n513), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n512), .ZN(
        round_inst_srout2_y[50]) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n519), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n510), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n519) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n507), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n509) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U130 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n506), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n507) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n508) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U128 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n503), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n502), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n513) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n501), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n500), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n502) );
  NOR3_X1 round_inst_S_8__sbox_inst_com_y_inst_U126 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n499), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n498), .A3(
        round_inst_S_8__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n500) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U125 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n496), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n495), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n501) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U124 ( .A1(
        round_inst_sin_x[35]), .A2(round_inst_S_8__sbox_inst_com_y_inst_n494), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n495) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U123 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n493), .A2(
        round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U122 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n492), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n491), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U121 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n490), .A2(round_inst_sin_w[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n492) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U120 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n489), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n488), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n503) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U119 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n487), .A2(
        round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n488) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U118 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n486), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n485), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n487) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U117 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n504), .A2(round_inst_sin_w[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n485) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n515), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n486) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U115 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n482), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n489) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n481), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n480), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n482) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U113 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n479), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U112 ( .A(
        round_inst_S_8__sbox_inst_n1), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n478), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n481) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n477), .B(round_inst_sin_x[31]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n478) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_y_inst_U110 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n515), .A2(
        round_inst_S_8__sbox_inst_n3), .A3(
        round_inst_S_8__sbox_inst_com_y_inst_n476), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n477) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U109 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n483) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_y_inst_U108 ( .A1(
        round_inst_sin_w[32]), .A2(round_inst_sin_w[35]), .A3(
        round_inst_S_8__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_8__sbox_inst_com_y_inst_U107 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n506), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_8__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U106 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[48]) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U105 ( .A1(
        round_inst_S_8__sbox_inst_n5), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U104 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n510), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U99 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_8__sbox_inst_n1), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U98 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U96 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n476), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n491) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_y_inst_U95 ( .A1(round_inst_sin_w[32]), .A2(round_inst_n66), .A3(round_inst_S_8__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U94 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U93 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U92 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U89 ( .A1(
        round_inst_S_8__sbox_inst_n1), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_8__sbox_inst_com_y_inst_U88 ( .A(
        round_inst_S_8__sbox_inst_n5), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n504), .S(
        round_inst_S_8__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U87 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U85 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U81 ( .A(
        round_inst_S_8__sbox_inst_n1), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n479), .B(round_inst_n65), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U79 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n479) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n515), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U77 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n438), .Z(round_inst_srout2_y[51]) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n484), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U72 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U71 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U70 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n484), .A2(round_inst_n66), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_8__sbox_inst_n1), .A2(round_inst_sin_w[32]), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[35]), 
        .A3(round_inst_S_8__sbox_inst_n1), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U67 ( .A(round_inst_sin_w[32]), 
        .B(round_inst_S_8__sbox_inst_com_y_inst_n476), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U66 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U64 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U62 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U60 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U59 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U58 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n484), .A2(round_inst_sin_w[33]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n422) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n418), .A2(
        round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U55 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U54 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U53 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n414), .B(round_inst_n66), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U51 ( .A(round_inst_sin_w[33]), 
        .B(round_inst_S_8__sbox_inst_n1), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U50 ( .A1(
        round_inst_S_8__sbox_inst_n1), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n476), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n444) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U49 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n473), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n476) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U48 ( .A(round_inst_sin_x[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_8__sbox_inst_n1), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U46 ( .A(round_inst_sin_x[30]), 
        .B(round_inst_S_8__sbox_inst_com_y_inst_n514), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n514) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[33]), 
        .B(round_inst_sin_x[35]), .Z(round_inst_S_8__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U41 ( .A(round_inst_n66), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n499) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n484), .B(round_inst_sin_w[32]), 
        .Z(round_inst_S_8__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n484) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U36 ( .A(round_inst_sin_z[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n497) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_8__sbox_inst_n1), .B(round_inst_S_8__sbox_inst_n3), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n490), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n498) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_8__sbox_inst_n5), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n506), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n490) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U27 ( .A1(round_inst_sin_w[33]), .A2(round_inst_S_8__sbox_inst_n3), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n515), .A2(round_inst_sin_w[33]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_8__sbox_inst_n1), .A2(round_inst_sin_w[35]), .A3(
        round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_8__sbox_inst_n1), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n505), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n506), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_8__sbox_inst_n3), .B(round_inst_sin_w[35]), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U17 ( .A(
        round_inst_S_8__sbox_inst_n3), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[35]), 
        .B(round_inst_sin_x[35]), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_y_inst_U13 ( .A1(round_inst_n66), 
        .A2(round_inst_sin_w[35]), .A3(
        round_inst_S_8__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_y_inst_U12 ( .A1(
        round_inst_S_8__sbox_inst_n3), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_8__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[33]), 
        .B(round_inst_n66), .S(round_inst_S_8__sbox_inst_com_y_inst_n504), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_y_inst_U9 ( .A1(round_inst_n66), .A2(
        round_inst_S_8__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_8__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_8__sbox_inst_n3), .B(round_inst_sin_x[35]), .Z(
        round_inst_S_8__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_8__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_8__sbox_inst_n1), .A3(round_inst_sin_x[35]), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n515), .B(
        round_inst_S_8__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n504) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[34]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_8__sbox_inst_com_y_inst_n506), .ZN(
        round_inst_S_8__sbox_inst_com_y_inst_n515) );
  INV_X1 round_inst_S_8__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[34]), 
        .ZN(round_inst_S_8__sbox_inst_com_y_inst_n506) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U132 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n517), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n516), .ZN(round_inst_sout_z[32])
         );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n515), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n514), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U130 ( .A(round_inst_sin_w[34]), .B(round_inst_sin_w[35]), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n514) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_x[28]), 
        .B(round_inst_n50), .Z(round_inst_S_8__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U128 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n512), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n517) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_srout2_z[50]) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n510), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n509), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n511) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n508), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n507), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n509) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U124 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n506), .A2(round_inst_n52), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U123 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n505), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n504), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n508) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n503), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n502), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U121 ( .A(round_inst_sin_w[33]), .B(round_inst_sin_x[31]), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U120 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n501), .B(round_inst_sin_y[31]), 
        .Z(round_inst_S_8__sbox_inst_com_z_inst_n503) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U119 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n500), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n499), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n501) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U118 ( .A1(round_inst_n53), 
        .A2(round_inst_S_8__sbox_inst_com_z_inst_n498), .A3(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n499) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U117 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_x[32]), 
        .A3(round_inst_sin_w[35]), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n500) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U116 ( .A(
        round_inst_S_8__sbox_inst_n5), .B(round_inst_n53), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n496) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U115 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_8__sbox_inst_n5), .A3(
        round_inst_S_8__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n505) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U114 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n491), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n493) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n490), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n489), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n491) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U111 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n488), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n486), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n490) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_sin_w[34]), .A2(round_inst_S_8__sbox_inst_com_z_inst_n495), 
        .A3(round_inst_n52), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n492) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U108 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n484), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n513) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U107 ( .A1(
        round_inst_sin_w[34]), .A2(round_inst_S_8__sbox_inst_com_z_inst_n498), 
        .ZN(round_inst_S_8__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U106 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n506), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n484) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n482), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n481), .Z(round_inst_srout2_z[48]) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n479), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n478), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n483), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n483) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U101 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n475), .A2(round_inst_sin_x[32]), 
        .A3(round_inst_sin_w[34]), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U100 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n474), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n477) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U99 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n472), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .A3(round_inst_n53), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n473) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U98 ( .A(round_inst_sin_w[33]), 
        .B(round_inst_sin_y[33]), .Z(round_inst_S_8__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U97 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n471), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n474) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U96 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n469), .A2(
        round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n470) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U95 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n467), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n471) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n466), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n465), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n464), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n463), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n462), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n461), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U91 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n460), .A2(round_inst_n53), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n461) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U90 ( .A1(round_inst_n66), 
        .A2(round_inst_S_8__sbox_inst_n5), .A3(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n462) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U89 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n459), .A2(round_inst_n52), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_w[34]), 
        .ZN(round_inst_S_8__sbox_inst_com_z_inst_n466) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U87 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U85 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n453), .A2(round_inst_n53), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n454) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U84 ( .A(round_inst_sin_w[33]), 
        .B(round_inst_S_8__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U83 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n451), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U82 ( .A1(round_inst_sin_w[34]), .A2(round_inst_sin_x[32]), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n478) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U81 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n487), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n448) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U79 ( .A(round_inst_sin_y[29]), 
        .B(round_inst_n65), .Z(round_inst_S_8__sbox_inst_com_z_inst_n447) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U78 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n487) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n446), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U76 ( .A(round_inst_sin_w[34]), 
        .B(round_inst_n53), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U75 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_srout2_z[51]) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n512), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U72 ( .A1(round_inst_sin_x[32]), .A2(round_inst_sin_w[35]), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n441) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U71 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n458), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n440), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n442) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U70 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n498), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U69 ( .A(round_inst_sin_w[35]), 
        .B(round_inst_S_8__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n498) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U68 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n494) );
  MUX2_X1 round_inst_S_8__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n495), .B(round_inst_sin_w[35]), 
        .S(round_inst_S_8__sbox_inst_com_z_inst_n436), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n437) );
  OR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U66 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n436) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U65 ( .A(round_inst_sin_x[32]), 
        .B(round_inst_S_8__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n486) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U64 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n438) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U63 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n495), .A3(
        round_inst_S_8__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U62 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n430), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n429) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U59 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n426), .A2(round_inst_sin_w[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U58 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n422), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n424) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U56 ( .A1(round_inst_sin_x[32]), .A2(round_inst_n66), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U55 ( .A1(round_inst_sin_y[33]), .A2(round_inst_sin_x[32]), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n425) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U54 ( .A1(round_inst_n52), 
        .A2(round_inst_S_8__sbox_inst_com_z_inst_n495), .A3(
        round_inst_sin_w[33]), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n428)
         );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U53 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_y[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U52 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n460), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n423), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n469) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U50 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .A2(round_inst_sin_y[33]), 
        .ZN(round_inst_S_8__sbox_inst_com_z_inst_n423) );
  AND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U49 ( .A1(round_inst_sin_w[33]), 
        .A2(round_inst_sin_x[32]), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n460) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U48 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n421) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U47 ( .A1(round_inst_sin_w[33]), .A2(round_inst_S_8__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U46 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .A2(round_inst_n66), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n419), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n418), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n432) );
  INV_X1 round_inst_S_8__sbox_inst_com_z_inst_U44 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U43 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .B(round_inst_n52), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n451) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n417), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U41 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n497), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n449) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U39 ( .A1(round_inst_sin_w[35]), .A2(round_inst_S_8__sbox_inst_com_z_inst_n413), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n414) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U38 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n415) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U35 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n506), .A2(round_inst_n66), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n409) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U34 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n407) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U32 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n405) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n404) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U30 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n506), .A2(round_inst_sin_y[33]), 
        .ZN(round_inst_S_8__sbox_inst_com_z_inst_n402) );
  AND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_S_8__sbox_inst_n5), .A2(round_inst_sin_w[35]), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n506) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n401), .A2(round_inst_n53), .A3(
        round_inst_sin_w[33]), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n403)
         );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U27 ( .A(round_inst_sin_w[35]), 
        .B(round_inst_S_8__sbox_inst_com_z_inst_n495), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n401) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U26 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n399), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n406) );
  MUX2_X1 round_inst_S_8__sbox_inst_com_z_inst_U25 ( .A(round_inst_sin_y[35]), 
        .B(round_inst_S_8__sbox_inst_com_z_inst_n398), .S(
        round_inst_S_8__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U24 ( .A1(round_inst_sin_w[33]), .A2(round_inst_S_8__sbox_inst_n5), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U23 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n398) );
  NOR3_X1 round_inst_S_8__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n488), .A3(
        round_inst_S_8__sbox_inst_com_z_inst_n395), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U21 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n394), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n395) );
  INV_X1 round_inst_S_8__sbox_inst_com_z_inst_U20 ( .A(round_inst_n66), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n394) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U19 ( .A(round_inst_sin_w[35]), 
        .B(round_inst_sin_y[35]), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n488) );
  AND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U18 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n459), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U17 ( .A1(round_inst_sin_w[34]), .A2(round_inst_n66), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n459) );
  INV_X1 round_inst_S_8__sbox_inst_com_z_inst_U16 ( .A(round_inst_sin_w[33]), 
        .ZN(round_inst_S_8__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U15 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n393), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U14 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n391), .A2(round_inst_n53), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U13 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_8__sbox_inst_com_z_inst_n390), .Z(
        round_inst_S_8__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U12 ( .A1(round_inst_sin_w[33]), .A2(round_inst_sin_y[35]), .ZN(round_inst_S_8__sbox_inst_com_z_inst_n390) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U11 ( .A1(round_inst_n66), 
        .A2(round_inst_sin_w[35]), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n418) );
  NOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U10 ( .A1(
        round_inst_S_8__sbox_inst_com_z_inst_n439), .A2(
        round_inst_S_8__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_8__sbox_inst_com_z_inst_U9 ( .A1(round_inst_sin_w[34]), 
        .A2(round_inst_sin_w[33]), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n456) );
  XNOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U8 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n495), .B(round_inst_sin_y[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_z_inst_n439) );
  NAND3_X1 round_inst_S_8__sbox_inst_com_z_inst_U7 ( .A1(round_inst_sin_w[34]), 
        .A2(round_inst_S_8__sbox_inst_com_z_inst_n495), .A3(
        round_inst_S_8__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U6 ( .A(round_inst_n66), .B(
        round_inst_sin_y[33]), .Z(round_inst_S_8__sbox_inst_com_z_inst_n475)
         );
  INV_X1 round_inst_S_8__sbox_inst_com_z_inst_U5 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n495) );
  INV_X1 round_inst_S_8__sbox_inst_com_z_inst_U4 ( .A(round_inst_sin_x[35]), 
        .ZN(round_inst_S_8__sbox_inst_com_z_inst_n397) );
  INV_X1 round_inst_S_8__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_8__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_8__sbox_inst_com_z_inst_n497) );
  INV_X1 round_inst_S_8__sbox_inst_com_z_inst_U2 ( .A(round_inst_sin_w[32]), 
        .ZN(round_inst_S_8__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_8__sbox_inst_com_z_inst_U1 ( .A(round_inst_n51), .B(
        round_inst_sin_x[30]), .Z(round_inst_S_8__sbox_inst_com_z_inst_n417)
         );
  INV_X1 round_inst_S_9__sbox_inst_U10 ( .A(round_inst_sin_x[38]), .ZN(
        round_inst_S_9__sbox_inst_n8) );
  INV_X1 round_inst_S_9__sbox_inst_U9 ( .A(round_inst_sin_w[36]), .ZN(
        round_inst_S_9__sbox_inst_n10) );
  INV_X1 round_inst_S_9__sbox_inst_U8 ( .A(round_inst_sin_x[37]), .ZN(
        round_inst_S_9__sbox_inst_n6) );
  INV_X1 round_inst_S_9__sbox_inst_U7 ( .A(round_inst_sin_z[37]), .ZN(
        round_inst_S_9__sbox_inst_n2) );
  INV_X1 round_inst_S_9__sbox_inst_U6 ( .A(round_inst_sin_z[39]), .ZN(
        round_inst_S_9__sbox_inst_n4) );
  INV_X2 round_inst_S_9__sbox_inst_U5 ( .A(round_inst_S_9__sbox_inst_n6), .ZN(
        round_inst_S_9__sbox_inst_n5) );
  INV_X2 round_inst_S_9__sbox_inst_U4 ( .A(round_inst_S_9__sbox_inst_n4), .ZN(
        round_inst_S_9__sbox_inst_n3) );
  INV_X2 round_inst_S_9__sbox_inst_U3 ( .A(round_inst_S_9__sbox_inst_n8), .ZN(
        round_inst_S_9__sbox_inst_n7) );
  INV_X2 round_inst_S_9__sbox_inst_U2 ( .A(round_inst_S_9__sbox_inst_n2), .ZN(
        round_inst_S_9__sbox_inst_n1) );
  INV_X2 round_inst_S_9__sbox_inst_U1 ( .A(round_inst_S_9__sbox_inst_n10), 
        .ZN(round_inst_S_9__sbox_inst_n9) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n531), .ZN(round_inst_sout_w[39])
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U139 ( .A1(
        round_inst_sin_z[36]), .A2(round_inst_S_9__sbox_inst_com_w_inst_n528), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n526), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n524), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n526) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[38]), .A2(round_inst_S_9__sbox_inst_com_w_inst_n523), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n525) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n518), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n516), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n518) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n514), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n513), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n512), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n513) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_w_inst_U128 ( .A1(
        round_inst_S_9__sbox_inst_n7), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n510), .A3(
        round_inst_S_9__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n511) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U127 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n508), .A2(round_inst_n54), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n507), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U125 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n507) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_9__sbox_inst_n3), .A2(round_inst_n55), .A3(
        round_inst_S_9__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U122 ( .A(round_inst_sin_y[35]), .B(round_inst_S_9__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U121 ( .A(
        round_inst_S_9__sbox_inst_n5), .B(round_inst_sin_z[35]), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n501) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U120 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[37])
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[33]), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[33]), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U113 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[36])
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_9__sbox_inst_n7), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U110 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n528), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U105 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_9__sbox_inst_n7), .B(round_inst_sin_z[38]), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_9__sbox_inst_n1), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U99 ( .A1(round_inst_n55), 
        .A2(round_inst_S_9__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_9__sbox_inst_n7), .A2(round_inst_n54), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n506) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U94 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[38]), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n461), .A2(
        round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[38]), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U88 ( .A1(round_inst_sin_z[36]), 
        .A2(round_inst_S_9__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_w_inst_U85 ( .A1(round_inst_sin_y[37]), .A2(round_inst_n54), .A3(round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_w_inst_U84 ( .A1(round_inst_n55), 
        .A2(round_inst_S_9__sbox_inst_n5), .A3(round_inst_n54), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n528) );
  OR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_9__sbox_inst_n7), .B(round_inst_n55), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U80 ( .A(round_inst_n52), .B(
        round_inst_sin_z[32]), .Z(round_inst_S_9__sbox_inst_com_w_inst_n484)
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U79 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[39])
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U73 ( .A1(
        round_inst_S_9__sbox_inst_n3), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U71 ( .A1(round_inst_n55), 
        .A2(round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_9__sbox_inst_n7), .A2(round_inst_sin_y[37]), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U69 ( .A1(
        round_inst_S_9__sbox_inst_n1), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n508), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_9__sbox_inst_n7), .A2(round_inst_S_9__sbox_inst_n1), .A3(
        round_inst_S_9__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n439), .A2(
        round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n508), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_9__sbox_inst_n3), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n504) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U62 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n508) );
  INV_X1 round_inst_S_9__sbox_inst_com_w_inst_U61 ( .A(round_inst_n55), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U60 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U58 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U57 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U56 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U55 ( .A(round_inst_sin_y[37]), 
        .B(round_inst_S_9__sbox_inst_n1), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U54 ( .A1(
        round_inst_S_9__sbox_inst_n3), .A2(round_inst_S_9__sbox_inst_n1), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U52 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_w_inst_U51 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n505), .A3(
        round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U50 ( .A(round_inst_sin_y[37]), 
        .B(round_inst_S_9__sbox_inst_n5), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_w_inst_U49 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n505), .A2(round_inst_sin_y[37]), 
        .A3(round_inst_S_9__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U48 ( .A(round_inst_n55), .B(
        round_inst_sin_z[38]), .ZN(round_inst_S_9__sbox_inst_com_w_inst_n465)
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U47 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n520) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U45 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n421), .A2(
        round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U44 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U43 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n419), .A2(
        round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U42 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U40 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_9__sbox_inst_n1), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n521) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U38 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U37 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U36 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n510), .B(round_inst_sin_z[36]), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n498), .A2(
        round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U33 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U32 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U31 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U30 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U29 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U28 ( .A1(
        round_inst_S_9__sbox_inst_n5), .A2(round_inst_sin_z[36]), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U27 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n522), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U26 ( .A(
        round_inst_S_9__sbox_inst_n5), .B(round_inst_S_9__sbox_inst_n1), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U24 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n510), .A2(
        round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U22 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[37]), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U21 ( .A(round_inst_n54), .B(
        round_inst_sin_z[36]), .Z(round_inst_S_9__sbox_inst_com_w_inst_n418)
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U20 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U19 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U17 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n398), .A2(
        round_inst_S_9__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U15 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n498), .B(
        round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_9__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_9__sbox_inst_com_w_inst_U13 ( .A(round_inst_sin_y[39]), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_9__sbox_inst_n1), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U11 ( .A(
        round_inst_S_9__sbox_inst_n3), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n505), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U9 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_9__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_9__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U8 ( .A1(
        round_inst_S_9__sbox_inst_n5), .A2(round_inst_n54), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U7 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n510), .A2(round_inst_sin_y[37]), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n477) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_w_inst_U6 ( .A1(
        round_inst_S_9__sbox_inst_com_w_inst_n505), .A2(round_inst_n54), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n522) );
  INV_X1 round_inst_S_9__sbox_inst_com_w_inst_U5 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n505) );
  INV_X1 round_inst_S_9__sbox_inst_com_w_inst_U4 ( .A(round_inst_sin_x[39]), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n486) );
  INV_X1 round_inst_S_9__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_9__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_9__sbox_inst_com_w_inst_n510) );
  INV_X1 round_inst_S_9__sbox_inst_com_w_inst_U2 ( .A(round_inst_sin_x[36]), 
        .ZN(round_inst_S_9__sbox_inst_com_w_inst_n489) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_w_inst_U1 ( .A(round_inst_n53), .B(
        round_inst_sin_z[34]), .Z(round_inst_S_9__sbox_inst_com_w_inst_n402)
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n510), .ZN(round_inst_sout_x[36])
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n509), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n510) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U133 ( .A(round_inst_n55), .B(
        round_inst_sin_y[39]), .ZN(round_inst_S_9__sbox_inst_com_x_inst_n508)
         );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U132 ( .A(round_inst_sin_z[32]), 
        .B(round_inst_S_9__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n506), .Z(round_inst_srout2_x[6])
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U130 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U129 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n503), .A2(round_inst_sin_z[36]), 
        .ZN(round_inst_S_9__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U127 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U126 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U125 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U124 ( .A1(round_inst_n55), 
        .A2(round_inst_S_9__sbox_inst_n9), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U122 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U121 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U118 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_sin_y[39]), .A2(round_inst_S_9__sbox_inst_com_x_inst_n490), 
        .ZN(round_inst_S_9__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U115 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n487) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_x_inst_U114 ( .A1(
        round_inst_sin_z[38]), .A2(round_inst_S_9__sbox_inst_n9), .A3(
        round_inst_sin_y[39]), .ZN(round_inst_S_9__sbox_inst_com_x_inst_n489)
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n478), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n476), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n478) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n475), .B(round_inst_sin_z[35]), 
        .ZN(round_inst_S_9__sbox_inst_com_x_inst_n476) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_w[38]), .A2(round_inst_sin_y[39]), .A3(
        round_inst_sin_z[36]), .ZN(round_inst_S_9__sbox_inst_com_x_inst_n475)
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n474), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n473), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n473) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n470), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n469), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n511) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n468), .A2(round_inst_n55), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n469) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n468) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n467), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n464), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n480), .ZN(round_inst_srout2_x[4]) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U100 ( .A1(round_inst_n54), 
        .A2(round_inst_sin_z[38]), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[33]), 
        .B(round_inst_S_9__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n464) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n462), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n460), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n467), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n461) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n458), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n467) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_9__sbox_inst_n1), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n457), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n459) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n455), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n454), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n456) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n453), .A2(round_inst_sin_w[38]), 
        .ZN(round_inst_S_9__sbox_inst_com_x_inst_n454) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n451), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n455) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n450), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n449), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n451) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n448), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n447), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n449) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n446), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_9__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n445), .B(round_inst_n55), .S(
        round_inst_n54), .Z(round_inst_S_9__sbox_inst_com_x_inst_n446) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n444), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n448) );
  MUX2_X1 round_inst_S_9__sbox_inst_com_x_inst_U85 ( .A(round_inst_n55), .B(
        round_inst_sin_z[38]), .S(round_inst_sin_z[36]), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n443), .A2(
        round_inst_S_9__sbox_inst_n9), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n442), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n441), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n452) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_9__sbox_inst_n9), .A3(round_inst_sin_z[38]), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n441) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n440), .A2(round_inst_sin_w[37]), 
        .A3(round_inst_n55), .ZN(round_inst_S_9__sbox_inst_com_x_inst_n442) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U80 ( .A(round_inst_n54), .B(
        round_inst_sin_z[36]), .Z(round_inst_S_9__sbox_inst_com_x_inst_n440)
         );
  NAND3_X1 round_inst_S_9__sbox_inst_com_x_inst_U79 ( .A1(round_inst_n54), 
        .A2(round_inst_S_9__sbox_inst_com_x_inst_n445), .A3(
        round_inst_S_9__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n460) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U77 ( .A1(round_inst_n54), 
        .A2(round_inst_n55), .ZN(round_inst_S_9__sbox_inst_com_x_inst_n482) );
  AND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U76 ( .A1(round_inst_n55), .A2(
        round_inst_sin_z[36]), .ZN(round_inst_S_9__sbox_inst_com_x_inst_n490)
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n462) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U74 ( .A1(round_inst_n54), 
        .A2(round_inst_sin_w[38]), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n497) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n437), .ZN(round_inst_srout2_x[7]) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n436), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n435), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U71 ( .A(round_inst_n54), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n435) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n434), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n433), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U69 ( .A1(round_inst_sin_z[36]), .A2(round_inst_sin_y[39]), .ZN(round_inst_S_9__sbox_inst_com_x_inst_n433) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n432), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n431), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n434) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n430), .A2(round_inst_n54), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n431) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n429), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n428), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_9__sbox_inst_n1), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n453), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n432) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[34]), 
        .B(round_inst_S_9__sbox_inst_com_x_inst_n438), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n436) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n425), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n424), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n423), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n422), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n421), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n420), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n422) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n419), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n420) );
  NOR3_X1 round_inst_S_9__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n471), .A3(
        round_inst_S_9__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n418) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n416), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n419) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n414), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U53 ( .A1(round_inst_n55), 
        .A2(round_inst_S_9__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n413) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U52 ( .A(round_inst_sin_y[39]), 
        .ZN(round_inst_S_9__sbox_inst_com_x_inst_n414) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n443), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n416) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U50 ( .A1(
        round_inst_S_9__sbox_inst_n1), .A2(round_inst_n55), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n443) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_x_inst_U49 ( .A1(round_inst_n55), 
        .A2(round_inst_S_9__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_9__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n421) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n411), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n423) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U47 ( .A1(round_inst_n55), 
        .A2(round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n465) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n411) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n410), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n407), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U43 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n406), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n405), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n407) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U42 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n466), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n405) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U41 ( .A(round_inst_sin_w[37]), 
        .B(round_inst_S_9__sbox_inst_n1), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n439) );
  AND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U40 ( .A1(round_inst_sin_z[38]), 
        .A2(round_inst_sin_y[39]), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_9__sbox_inst_n3), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n406) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_x_inst_U38 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U37 ( .A(round_inst_sin_z[38]), 
        .B(round_inst_sin_w[38]), .Z(round_inst_S_9__sbox_inst_com_x_inst_n445) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U36 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n404), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n410) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U35 ( .A(round_inst_sin_w[38]), 
        .B(round_inst_n55), .Z(round_inst_S_9__sbox_inst_com_x_inst_n403) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n402), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n401), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U33 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n400), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n399), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n401) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U32 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n399) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U31 ( .A1(round_inst_sin_z[36]), .A2(round_inst_S_9__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n426) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n427), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n400) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U28 ( .A(round_inst_sin_y[39]), 
        .B(round_inst_S_9__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n471) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n402) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_9__sbox_inst_n1), .A3(round_inst_n54), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n396) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n398), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n481) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U23 ( .A(round_inst_sin_y[39]), 
        .B(round_inst_S_9__sbox_inst_n3), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U21 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n392), .A2(
        round_inst_S_9__sbox_inst_n9), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n404), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_x_inst_U17 ( .A1(round_inst_sin_z[36]), .A2(round_inst_sin_y[39]), .A3(round_inst_sin_w[37]), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n388) );
  MUX2_X1 round_inst_S_9__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n412), .B(round_inst_sin_y[39]), 
        .S(round_inst_S_9__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U15 ( .A1(round_inst_n54), 
        .A2(round_inst_S_9__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U14 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n491), .B(
        round_inst_S_9__sbox_inst_n3), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n412) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n384), .A2(round_inst_sin_z[36]), 
        .ZN(round_inst_S_9__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U10 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_9__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U9 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_w[39]), 
        .ZN(round_inst_S_9__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U7 ( .A1(
        round_inst_S_9__sbox_inst_n1), .A2(round_inst_sin_y[39]), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n404) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_9__sbox_inst_com_x_inst_n427), .Z(
        round_inst_S_9__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U4 ( .A1(round_inst_n54), .A2(
        round_inst_sin_w[37]), .ZN(round_inst_S_9__sbox_inst_com_x_inst_n427)
         );
  NAND2_X1 round_inst_S_9__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_9__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_9__sbox_inst_n9), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_9__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_9__sbox_inst_com_x_inst_n477) );
  INV_X1 round_inst_S_9__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_y[37]), 
        .ZN(round_inst_S_9__sbox_inst_com_x_inst_n417) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n517), .Z(round_inst_sout_y[36])
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n516), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n515) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U134 ( .A(round_inst_sin_x[32]), 
        .B(round_inst_S_9__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n512), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n511), .ZN(round_inst_srout2_y[6]) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n508), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n518) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n507), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n506), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n508) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n506) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n507) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_9__sbox_inst_com_y_inst_U125 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_9__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U124 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U123 ( .A1(
        round_inst_sin_x[39]), .A2(round_inst_S_9__sbox_inst_com_y_inst_n493), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n492), .A2(
        round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U121 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U120 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n489), .A2(
        round_inst_S_9__sbox_inst_n9), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U119 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U118 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n486), .A2(
        round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U117 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_9__sbox_inst_n9), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U112 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_9__sbox_inst_n1), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[35]), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_y_inst_U109 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_9__sbox_inst_n3), .A3(round_inst_sin_x[36]), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U108 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_y_inst_U107 ( .A1(
        round_inst_S_9__sbox_inst_n9), .A2(round_inst_sin_w[39]), .A3(
        round_inst_S_9__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_9__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_9__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U105 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n470), .ZN(round_inst_srout2_y[4]) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U104 ( .A1(
        round_inst_S_9__sbox_inst_n7), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U98 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_9__sbox_inst_n1), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U95 ( .A1(round_inst_sin_x[36]), .A2(round_inst_S_9__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_y_inst_U94 ( .A1(
        round_inst_S_9__sbox_inst_n9), .A2(round_inst_S_9__sbox_inst_n5), .A3(
        round_inst_S_9__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U93 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U92 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U88 ( .A1(
        round_inst_S_9__sbox_inst_n1), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_9__sbox_inst_com_y_inst_U87 ( .A(
        round_inst_S_9__sbox_inst_n7), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n503), .S(
        round_inst_S_9__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_9__sbox_inst_n1), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n478), .B(round_inst_n66), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n438), .Z(round_inst_srout2_y[7])
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U71 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[39]), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U70 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n483), .A2(
        round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_9__sbox_inst_n1), .A2(round_inst_S_9__sbox_inst_n9), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[39]), 
        .A3(round_inst_S_9__sbox_inst_n1), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U66 ( .A(
        round_inst_S_9__sbox_inst_n9), .B(round_inst_sin_x[36]), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U59 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[39]), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U58 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[37]), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U55 ( .A(round_inst_sin_x[36]), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U54 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n418), .A2(
        round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U53 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U51 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n415), .A2(
        round_inst_S_9__sbox_inst_n9), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U50 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n414), .B(
        round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U49 ( .A(round_inst_sin_w[37]), 
        .B(round_inst_S_9__sbox_inst_n1), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U48 ( .A1(
        round_inst_S_9__sbox_inst_n1), .A2(round_inst_sin_x[36]), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_9__sbox_inst_n1), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U46 ( .A(round_inst_sin_x[34]), 
        .B(round_inst_S_9__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n513) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[37]), 
        .B(round_inst_sin_x[39]), .Z(round_inst_S_9__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U41 ( .A(
        round_inst_S_9__sbox_inst_n5), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[39]), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_9__sbox_inst_n9), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U36 ( .A(round_inst_sin_z[36]), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_9__sbox_inst_n1), .B(round_inst_S_9__sbox_inst_n3), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_9__sbox_inst_n7), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U27 ( .A1(round_inst_sin_w[37]), .A2(round_inst_S_9__sbox_inst_n3), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n514), .A2(round_inst_sin_w[37]), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_9__sbox_inst_n1), .A2(round_inst_sin_w[39]), .A3(
        round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_9__sbox_inst_n1), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n504), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_9__sbox_inst_n3), .B(round_inst_sin_w[39]), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U17 ( .A(
        round_inst_S_9__sbox_inst_n3), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[39]), 
        .B(round_inst_sin_x[39]), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_y_inst_U13 ( .A1(
        round_inst_S_9__sbox_inst_n5), .A2(round_inst_sin_w[39]), .A3(
        round_inst_S_9__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_y_inst_U12 ( .A1(
        round_inst_S_9__sbox_inst_n3), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_9__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[37]), 
        .B(round_inst_S_9__sbox_inst_n5), .S(
        round_inst_S_9__sbox_inst_com_y_inst_n503), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_y_inst_U9 ( .A1(
        round_inst_S_9__sbox_inst_n5), .A2(
        round_inst_S_9__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_9__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_9__sbox_inst_n3), .B(round_inst_sin_x[39]), .Z(
        round_inst_S_9__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_9__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_9__sbox_inst_n1), .A3(round_inst_sin_x[39]), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_9__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n503) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[38]), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_9__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_9__sbox_inst_com_y_inst_n514) );
  INV_X1 round_inst_S_9__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[38]), 
        .ZN(round_inst_S_9__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U132 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n516), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n515), .ZN(round_inst_sout_z[36])
         );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n514), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n513), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U130 ( .A(round_inst_sin_w[38]), .B(round_inst_sin_w[39]), .ZN(round_inst_S_9__sbox_inst_com_z_inst_n513) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_x[32]), 
        .B(round_inst_n52), .Z(round_inst_S_9__sbox_inst_com_z_inst_n514) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U128 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n510), .ZN(round_inst_srout2_z[6]) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n509), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n508), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n507), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n506), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n508) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U124 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n505), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n504), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n506) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U123 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n503), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n502), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U122 ( .A(round_inst_sin_w[37]), .B(round_inst_S_9__sbox_inst_com_z_inst_n501), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n500), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n499), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n501) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_z_inst_U120 ( .A1(
        round_inst_S_9__sbox_inst_n7), .A2(round_inst_sin_x[39]), .A3(
        round_inst_S_9__sbox_inst_n9), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n499) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U119 ( .A1(round_inst_n54), 
        .A2(round_inst_S_9__sbox_inst_com_z_inst_n498), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n500) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U118 ( .A(round_inst_sin_y[35]), 
        .B(round_inst_sin_x[35]), .Z(round_inst_S_9__sbox_inst_com_z_inst_n503) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_z_inst_U117 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n497), .A2(round_inst_sin_x[36]), 
        .A3(round_inst_sin_w[39]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n505) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U116 ( .A(
        round_inst_S_9__sbox_inst_n7), .B(round_inst_n55), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n497) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U115 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U114 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n509) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n491), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n493) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n490), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n489), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n491) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U111 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n488), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n486), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n490) );
  INV_X1 round_inst_S_9__sbox_inst_com_z_inst_U109 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n484), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n486) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_z_inst_U108 ( .A1(
        round_inst_sin_w[38]), .A2(round_inst_sin_x[39]), .A3(round_inst_n54), 
        .ZN(round_inst_S_9__sbox_inst_com_z_inst_n492) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U107 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U106 ( .A1(
        round_inst_sin_w[38]), .A2(round_inst_S_9__sbox_inst_com_z_inst_n482), 
        .ZN(round_inst_S_9__sbox_inst_com_z_inst_n485) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n481), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n480), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n483) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n479), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n478), .ZN(round_inst_srout2_z[4]) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n481), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n478) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n476), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U101 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n474), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n475) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U100 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n472), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n471), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n473) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_z_inst_U99 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n470), .A2(round_inst_sin_x[36]), 
        .A3(round_inst_sin_w[38]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n471) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_z_inst_U98 ( .A1(
        round_inst_S_9__sbox_inst_n9), .A2(round_inst_n55), .A3(
        round_inst_sin_w[37]), .ZN(round_inst_S_9__sbox_inst_com_z_inst_n472)
         );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U97 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n469), .A2(round_inst_sin_w[38]), 
        .ZN(round_inst_S_9__sbox_inst_com_z_inst_n474) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U96 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n467), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n476) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U95 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n466), .A2(
        round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n467) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n465), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n464), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n463), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n462), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n464) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n461), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n460), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U91 ( .A1(round_inst_sin_w[37]), .A2(round_inst_n55), .ZN(round_inst_S_9__sbox_inst_com_z_inst_n460) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U90 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n459), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n458), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n461) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U89 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n457), .A2(round_inst_n55), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n458) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n456), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n455), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n459) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U87 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n454), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n453), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n465) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n451), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n453) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U85 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n450), .A2(round_inst_n55), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n451) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U84 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n449), .A2(round_inst_n54), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U83 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n448), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n454) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_S_9__sbox_inst_n9), .A2(round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n447) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U81 ( .A(
        round_inst_S_9__sbox_inst_n7), .B(round_inst_n55), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n448) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U80 ( .A1(round_inst_sin_w[38]), .A2(round_inst_sin_x[36]), .ZN(round_inst_S_9__sbox_inst_com_z_inst_n477) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U79 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n446), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U78 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n445) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_9__sbox_inst_n9), .A2(round_inst_sin_w[38]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U76 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n487), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n442), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n444) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U75 ( .A1(
        round_inst_S_9__sbox_inst_n9), .A2(round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n487) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n496), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n446) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U73 ( .A(round_inst_sin_y[33]), 
        .B(round_inst_n66), .Z(round_inst_S_9__sbox_inst_com_z_inst_n441) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U72 ( .A1(
        round_inst_S_9__sbox_inst_n9), .A2(round_inst_n55), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n496) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U71 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n440), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n439), .ZN(round_inst_srout2_z[7]) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U70 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n511), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n439) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U69 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n511) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U68 ( .A1(round_inst_sin_x[36]), .A2(round_inst_sin_w[39]), .ZN(round_inst_S_9__sbox_inst_com_z_inst_n437) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n469), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n436), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n438) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U66 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n482), .A2(
        round_inst_S_9__sbox_inst_n9), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n436) );
  INV_X1 round_inst_S_9__sbox_inst_com_z_inst_U65 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U64 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n466), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n435), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n469) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U63 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n494) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U62 ( .A1(round_inst_sin_w[39]), .A2(round_inst_S_9__sbox_inst_com_z_inst_n432), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n433) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n431), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n430), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n432) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U60 ( .A1(round_inst_sin_x[36]), .A2(round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U59 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n429), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n428), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U58 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n427), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n426), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n428) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n426) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U56 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n422), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n424) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_z_inst_U55 ( .A1(round_inst_sin_x[36]), .A2(round_inst_sin_y[37]), .A3(round_inst_sin_w[39]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n422) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_z_inst_U54 ( .A1(round_inst_n54), 
        .A2(round_inst_sin_x[39]), .A3(round_inst_sin_w[37]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n423) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U53 ( .A1(round_inst_sin_y[39]), .A2(round_inst_S_9__sbox_inst_com_z_inst_n466), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n425) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U52 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n466) );
  INV_X1 round_inst_S_9__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n450) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U50 ( .A1(
        round_inst_S_9__sbox_inst_n9), .A2(round_inst_sin_y[37]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n431) );
  AND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U49 ( .A1(round_inst_sin_w[37]), 
        .A2(round_inst_sin_x[36]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n457) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U48 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n427) );
  MUX2_X1 round_inst_S_9__sbox_inst_com_z_inst_U47 ( .A(round_inst_sin_x[39]), 
        .B(round_inst_sin_w[39]), .S(round_inst_S_9__sbox_inst_com_z_inst_n419), .Z(round_inst_S_9__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U46 ( .A1(round_inst_sin_w[37]), .A2(round_inst_S_9__sbox_inst_com_z_inst_n484), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U45 ( .A(round_inst_sin_x[36]), 
        .B(round_inst_S_9__sbox_inst_n9), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n484) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U44 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n417), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n421) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_z_inst_U43 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n456), .A2(round_inst_sin_w[39]), 
        .A3(round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n417) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_9__sbox_inst_n9), .B(round_inst_n54), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n456) );
  OR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U41 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n418) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U40 ( .A1(
        round_inst_S_9__sbox_inst_n9), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n415), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n435) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_z_inst_U39 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n470), .A2(
        round_inst_S_9__sbox_inst_n9), .A3(round_inst_sin_x[39]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n429) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U38 ( .A(round_inst_sin_y[37]), 
        .B(round_inst_S_9__sbox_inst_n5), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n470) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n414), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n413), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_9__sbox_inst_n9), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n442), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U35 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n442) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U34 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n409), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U33 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n498), .A2(round_inst_sin_y[37]), 
        .ZN(round_inst_S_9__sbox_inst_com_z_inst_n409) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U32 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n462), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n410) );
  INV_X1 round_inst_S_9__sbox_inst_com_z_inst_U31 ( .A(round_inst_sin_y[39]), 
        .ZN(round_inst_S_9__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U30 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n412) );
  NAND3_X1 round_inst_S_9__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n406), .A2(round_inst_sin_w[38]), 
        .A3(round_inst_sin_x[39]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n407) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U28 ( .A(round_inst_sin_y[37]), 
        .B(round_inst_sin_w[37]), .Z(round_inst_S_9__sbox_inst_com_z_inst_n406) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U27 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n405), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n408) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U26 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n404) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U25 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n401), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n400), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n402) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U24 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n399), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n398), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U23 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n455), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n398) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U22 ( .A(round_inst_sin_w[39]), 
        .B(round_inst_S_9__sbox_inst_com_z_inst_n397), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n495) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U21 ( .A(round_inst_sin_y[39]), 
        .B(round_inst_sin_x[39]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n397) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U20 ( .A1(round_inst_sin_w[37]), .A2(round_inst_S_9__sbox_inst_n7), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U19 ( .A1(round_inst_sin_w[37]), .A2(round_inst_S_9__sbox_inst_com_z_inst_n396), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n399) );
  MUX2_X1 round_inst_S_9__sbox_inst_com_z_inst_U18 ( .A(round_inst_sin_x[39]), 
        .B(round_inst_sin_y[39]), .S(round_inst_n55), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n396) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U17 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n395), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n394), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n401) );
  INV_X1 round_inst_S_9__sbox_inst_com_z_inst_U16 ( .A(round_inst_sin_w[39]), 
        .ZN(round_inst_S_9__sbox_inst_com_z_inst_n394) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U15 ( .A(
        round_inst_S_9__sbox_inst_n5), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n393), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n395) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U14 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n462), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U13 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n415), .A2(round_inst_n55), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U12 ( .A(round_inst_sin_w[37]), 
        .B(round_inst_S_9__sbox_inst_n5), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n415) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U11 ( .A1(round_inst_sin_w[38]), .A2(round_inst_sin_w[37]), .ZN(round_inst_S_9__sbox_inst_com_z_inst_n462) );
  NOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U10 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n488), .A2(
        round_inst_S_9__sbox_inst_com_z_inst_n391), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n403) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U9 ( .A(round_inst_sin_w[37]), 
        .B(round_inst_S_9__sbox_inst_com_z_inst_n449), .Z(
        round_inst_S_9__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U8 ( .A1(round_inst_sin_w[38]), 
        .A2(round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n449) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U7 ( .A(round_inst_sin_w[39]), 
        .B(round_inst_sin_y[39]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n488) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U6 ( .A1(
        round_inst_S_9__sbox_inst_com_z_inst_n390), .A2(
        round_inst_S_9__sbox_inst_n5), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n405) );
  XNOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U5 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n389), .B(
        round_inst_S_9__sbox_inst_com_z_inst_n498), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n390) );
  INV_X1 round_inst_S_9__sbox_inst_com_z_inst_U4 ( .A(
        round_inst_S_9__sbox_inst_com_z_inst_n480), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n498) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U3 ( .A1(
        round_inst_S_9__sbox_inst_n7), .A2(round_inst_sin_w[39]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n480) );
  NAND2_X1 round_inst_S_9__sbox_inst_com_z_inst_U2 ( .A1(round_inst_sin_x[39]), 
        .A2(round_inst_sin_w[38]), .ZN(
        round_inst_S_9__sbox_inst_com_z_inst_n389) );
  XOR2_X1 round_inst_S_9__sbox_inst_com_z_inst_U1 ( .A(round_inst_n53), .B(
        round_inst_sin_x[34]), .Z(round_inst_S_9__sbox_inst_com_z_inst_n414)
         );
  INV_X1 round_inst_S_10__sbox_inst_U6 ( .A(round_inst_sin_x[41]), .ZN(
        round_inst_S_10__sbox_inst_n4) );
  INV_X1 round_inst_S_10__sbox_inst_U5 ( .A(round_inst_sin_x[42]), .ZN(
        round_inst_S_10__sbox_inst_n6) );
  INV_X1 round_inst_S_10__sbox_inst_U4 ( .A(round_inst_sin_z[41]), .ZN(
        round_inst_S_10__sbox_inst_n2) );
  INV_X2 round_inst_S_10__sbox_inst_U3 ( .A(round_inst_S_10__sbox_inst_n4), 
        .ZN(round_inst_S_10__sbox_inst_n3) );
  INV_X2 round_inst_S_10__sbox_inst_U2 ( .A(round_inst_S_10__sbox_inst_n6), 
        .ZN(round_inst_S_10__sbox_inst_n5) );
  INV_X2 round_inst_S_10__sbox_inst_U1 ( .A(round_inst_S_10__sbox_inst_n2), 
        .ZN(round_inst_S_10__sbox_inst_n1) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n531), .ZN(round_inst_sout_w[43]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U139 ( .A1(
        round_inst_sin_z[40]), .A2(round_inst_S_10__sbox_inst_com_w_inst_n528), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n526), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n524), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n526) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[42]), .A2(round_inst_S_10__sbox_inst_com_w_inst_n523), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n525) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n518), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n516), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n518) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n514), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n513), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n512), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n513) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_w_inst_U128 ( .A1(
        round_inst_S_10__sbox_inst_n5), .A2(round_inst_sin_x[40]), .A3(
        round_inst_S_10__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n511) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U127 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n509), .A2(round_inst_sin_y[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n508), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n507), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U125 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n508) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_sin_z[43]), .A2(round_inst_S_10__sbox_inst_com_w_inst_n504), 
        .A3(round_inst_sin_x[40]), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U122 ( .A(
        round_inst_sin_y[39]), .B(round_inst_S_10__sbox_inst_com_w_inst_n501), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U121 ( .A(
        round_inst_S_10__sbox_inst_n3), .B(round_inst_sin_z[39]), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n501) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U120 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[41]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[37]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[37]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U113 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[40]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_10__sbox_inst_n5), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U110 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n528), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U105 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_10__sbox_inst_n5), .B(round_inst_sin_z[42]), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_10__sbox_inst_n1), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U99 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n504), .A2(round_inst_sin_x[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_10__sbox_inst_n5), .A2(round_inst_sin_y[40]), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n507) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U94 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n461), .A2(
        round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U88 ( .A1(round_inst_sin_z[40]), .A2(round_inst_S_10__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_w_inst_U85 ( .A1(
        round_inst_sin_y[41]), .A2(round_inst_sin_y[40]), .A3(
        round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_w_inst_U84 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_10__sbox_inst_n3), .A3(round_inst_sin_y[40]), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n528) );
  OR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_10__sbox_inst_n5), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U80 ( .A(round_inst_n54), .B(
        round_inst_sin_z[36]), .Z(round_inst_S_10__sbox_inst_com_w_inst_n484)
         );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U79 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[43])
         );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U73 ( .A1(
        round_inst_sin_z[43]), .A2(round_inst_S_10__sbox_inst_com_w_inst_n440), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U71 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_10__sbox_inst_n5), .A2(round_inst_sin_y[41]), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U69 ( .A1(
        round_inst_S_10__sbox_inst_n1), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_10__sbox_inst_n5), .A2(round_inst_S_10__sbox_inst_n1), 
        .A3(round_inst_S_10__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n439), .A2(
        round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n505), .A2(
        round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U63 ( .A(round_inst_sin_z[43]), 
        .B(round_inst_S_10__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n505) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U62 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U61 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U60 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U58 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U57 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U56 ( .A(round_inst_sin_y[41]), .B(round_inst_S_10__sbox_inst_n1), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U55 ( .A1(
        round_inst_sin_z[43]), .A2(round_inst_S_10__sbox_inst_n1), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U54 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_w_inst_U52 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n506), .A3(
        round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U51 ( .A(round_inst_sin_y[41]), 
        .B(round_inst_S_10__sbox_inst_n3), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_w_inst_U50 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n506), .A2(round_inst_sin_y[41]), 
        .A3(round_inst_S_10__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U49 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n504), .B(round_inst_sin_z[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n465) );
  INV_X1 round_inst_S_10__sbox_inst_com_w_inst_U48 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n436), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n504) );
  INV_X1 round_inst_S_10__sbox_inst_com_w_inst_U47 ( .A(round_inst_sin_y[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U45 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n520) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U44 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n421), .A2(round_inst_sin_z[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U43 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U42 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n419), .A2(
        round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U40 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_10__sbox_inst_n1), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U38 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n521) );
  INV_X1 round_inst_S_10__sbox_inst_com_w_inst_U37 ( .A(round_inst_sin_x[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n489) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U36 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U33 ( .A(round_inst_sin_x[40]), .B(round_inst_sin_z[40]), .ZN(round_inst_S_10__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U32 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n498), .A2(
        round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U31 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U30 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U29 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U28 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U27 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U26 ( .A1(
        round_inst_S_10__sbox_inst_n3), .A2(round_inst_sin_z[40]), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n522), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U24 ( .A(
        round_inst_S_10__sbox_inst_n3), .B(round_inst_S_10__sbox_inst_n1), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_10__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U22 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U21 ( .A1(
        round_inst_sin_x[40]), .A2(round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U20 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[41]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U19 ( .A(round_inst_sin_y[40]), 
        .B(round_inst_sin_z[40]), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n418) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U17 ( .A(round_inst_sin_x[40]), .B(round_inst_S_10__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U15 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n398), .A2(round_inst_sin_x[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U13 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n498), .B(
        round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_10__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_10__sbox_inst_com_w_inst_U11 ( .A(round_inst_sin_y[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_10__sbox_inst_n1), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U9 ( .A(round_inst_sin_z[43]), 
        .B(round_inst_S_10__sbox_inst_com_w_inst_n506), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n510) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U8 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U7 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_10__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_10__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U6 ( .A1(
        round_inst_S_10__sbox_inst_n3), .A2(round_inst_sin_y[40]), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U5 ( .A1(round_inst_sin_x[40]), .A2(round_inst_sin_y[41]), .ZN(round_inst_S_10__sbox_inst_com_w_inst_n477)
         );
  NAND2_X1 round_inst_S_10__sbox_inst_com_w_inst_U4 ( .A1(
        round_inst_S_10__sbox_inst_com_w_inst_n506), .A2(round_inst_sin_y[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n522) );
  INV_X1 round_inst_S_10__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_10__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_10__sbox_inst_com_w_inst_n506) );
  INV_X1 round_inst_S_10__sbox_inst_com_w_inst_U2 ( .A(round_inst_sin_x[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_w_inst_n486) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_w_inst_U1 ( .A(round_inst_n55), .B(
        round_inst_sin_z[38]), .Z(round_inst_S_10__sbox_inst_com_w_inst_n402)
         );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U144 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n519), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n518), .Z(round_inst_sout_x[40])
         );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U143 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n517), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n516), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n518) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U142 ( .A(
        round_inst_sin_y[42]), .B(round_inst_sin_y[43]), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n516) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U141 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n515), .B(round_inst_sin_z[36]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n517) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U140 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n514), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n513), .ZN(
        round_inst_srout2_x[26]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U139 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n512), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n511), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n513) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U138 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n510), .A2(round_inst_sin_z[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n511) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U137 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n509), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n510) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U136 ( .A1(
        round_inst_sin_y[42]), .A2(round_inst_S_10__sbox_inst_com_x_inst_n507), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n508) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n506), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n505), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n512) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n504), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n503), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n505) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U133 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n509), .A2(round_inst_sin_w[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U132 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n501), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n504) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n501) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_x_inst_U130 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n497), .A3(round_inst_sin_y[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n499) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U129 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n496), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n495), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n500) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_x_inst_U128 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n494), .A2(round_inst_sin_y[40]), 
        .A3(round_inst_sin_y[42]), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n495) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U127 ( .A(round_inst_sin_y[43]), .B(round_inst_sin_z[43]), .Z(round_inst_S_10__sbox_inst_com_x_inst_n494) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U126 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n493), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n496) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_x_inst_U125 ( .A1(
        round_inst_sin_y[42]), .A2(round_inst_sin_z[40]), .A3(
        round_inst_sin_z[43]), .ZN(round_inst_S_10__sbox_inst_com_x_inst_n502)
         );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U124 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n492), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n506) );
  OR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U123 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n493), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n491) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U122 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U121 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n488) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n484), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n486) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n483), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n484) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U118 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n507), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n482) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U117 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n480), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n479), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n483) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U116 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n478), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n479) );
  AND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U115 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n481), .A2(round_inst_sin_z[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n477) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U114 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .B(round_inst_sin_z[39]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n478) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_x_inst_U113 ( .A1(
        round_inst_sin_y[42]), .A2(round_inst_sin_w[40]), .A3(
        round_inst_sin_z[43]), .ZN(round_inst_S_10__sbox_inst_com_x_inst_n480)
         );
  NAND3_X1 round_inst_S_10__sbox_inst_com_x_inst_U112 ( .A1(
        round_inst_sin_y[42]), .A2(round_inst_sin_y[40]), .A3(
        round_inst_S_10__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U111 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n475), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n493), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n487) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_y[42]), .A2(round_inst_sin_z[40]), .A3(
        round_inst_sin_y[43]), .ZN(round_inst_S_10__sbox_inst_com_x_inst_n489)
         );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n519), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n474), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n514) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U108 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n473), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n519) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n471), .A2(round_inst_sin_y[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n472) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_sin_z[43]), .B(round_inst_S_10__sbox_inst_com_x_inst_n470), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n471) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U105 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n509), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n473) );
  AND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U104 ( .A1(
        round_inst_sin_z[42]), .A2(round_inst_sin_y[43]), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n509) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n468), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n467), .ZN(
        round_inst_srout2_x[24]) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n493), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n467) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U101 ( .A1(
        round_inst_sin_y[40]), .A2(round_inst_sin_z[42]), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n493) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U100 ( .A1(
        round_inst_sin_y[42]), .A2(round_inst_S_10__sbox_inst_com_x_inst_n498), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n466) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U99 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n465), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n468) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n463), .B(round_inst_sin_z[37]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n464) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n463) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U96 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n462), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n481) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U95 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n460), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n459), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n469) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U94 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n458), .A2(round_inst_sin_y[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n459) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n457), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n458) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_10__sbox_inst_n1), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n498), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n455), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n454), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n460) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U90 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n453), .A2(round_inst_sin_w[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n454) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n451), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n453) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_sin_y[42]), .A2(round_inst_S_10__sbox_inst_n1), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n452) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n450), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n449), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n455) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U86 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n448), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n447), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n449) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U85 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n446), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n445), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n447) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n443), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n445) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n497), .B(round_inst_sin_z[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n443) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U82 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n442), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n441), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n440), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n448) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U80 ( .A1(
        round_inst_sin_y[42]), .A2(round_inst_sin_z[40]), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n441) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_x_inst_U79 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n498), .A3(
        round_inst_S_10__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U78 ( .A(round_inst_sin_z[42]), 
        .B(round_inst_S_10__sbox_inst_com_x_inst_n497), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n439) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U77 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n515), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_srout2_x[27]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U76 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n437), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n436), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U75 ( .A(round_inst_sin_y[40]), .B(round_inst_S_10__sbox_inst_com_x_inst_n474), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n436) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U74 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n435), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n434), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n433), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n432), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n434) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U72 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n431), .A2(round_inst_sin_w[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n432) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U71 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n430), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n429), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n431) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U70 ( .A1(
        round_inst_S_10__sbox_inst_n1), .A2(round_inst_sin_y[43]), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n429) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U69 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_z[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n428), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n433) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U67 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n426), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n427) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n424), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n423), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n422), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n421), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n423) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U64 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n507), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n421) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U63 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n440), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n456) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .B(round_inst_sin_w[41]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n440) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U61 ( .A1(
        round_inst_sin_z[43]), .A2(round_inst_S_10__sbox_inst_com_x_inst_n442), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n422) );
  AND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U60 ( .A1(round_inst_sin_y[40]), .A2(round_inst_S_10__sbox_inst_com_x_inst_n420), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n442) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_x_inst_U59 ( .A1(
        round_inst_sin_w[41]), .A2(round_inst_S_10__sbox_inst_com_x_inst_n498), 
        .A3(round_inst_sin_y[43]), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U58 ( .A(round_inst_sin_z[40]), 
        .B(round_inst_sin_y[40]), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n498) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U57 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n419), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n426) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_10__sbox_inst_n1), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n416), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n417) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n470), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n416) );
  MUX2_X1 round_inst_S_10__sbox_inst_com_x_inst_U53 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n419), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n414), .S(
        round_inst_S_10__sbox_inst_com_x_inst_n413), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n435) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U52 ( .A1(
        round_inst_sin_y[43]), .A2(round_inst_S_10__sbox_inst_com_x_inst_n412), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n413) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_y[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n412) );
  MUX2_X1 round_inst_S_10__sbox_inst_com_x_inst_U50 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n411), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n410), .S(
        round_inst_S_10__sbox_inst_com_x_inst_n409), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n414) );
  NOR3_X1 round_inst_S_10__sbox_inst_com_x_inst_U49 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n410), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n462), .A3(
        round_inst_S_10__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n411) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n475), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n419), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n410) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U47 ( .A(round_inst_sin_z[38]), 
        .B(round_inst_S_10__sbox_inst_com_x_inst_n465), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n407), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n406), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n465) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U45 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n405), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n406) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n405) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U43 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n418), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n404) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U42 ( .A(round_inst_sin_z[43]), .B(round_inst_S_10__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n418) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U41 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n403), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n402), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n407) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_x_inst_U40 ( .A1(
        round_inst_sin_z[42]), .A2(round_inst_sin_y[43]), .A3(
        round_inst_S_10__sbox_inst_com_x_inst_n401), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n402) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U39 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n420), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n401) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U38 ( .A(
        round_inst_S_10__sbox_inst_n1), .B(round_inst_sin_w[41]), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n420) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U37 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n400), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n399), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n403) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U36 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n446), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n399) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U35 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n475), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n398), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n397), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n400) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U33 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n490), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n451), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n397) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U32 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n396), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n395), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U31 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n395) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U30 ( .A1(
        round_inst_sin_y[43]), .A2(round_inst_S_10__sbox_inst_com_x_inst_n392), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n393) );
  MUX2_X1 round_inst_S_10__sbox_inst_com_x_inst_U29 ( .A(
        round_inst_S_10__sbox_inst_n1), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .S(
        round_inst_S_10__sbox_inst_com_x_inst_n497), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n392) );
  INV_X1 round_inst_S_10__sbox_inst_com_x_inst_U28 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n497) );
  INV_X1 round_inst_S_10__sbox_inst_com_x_inst_U27 ( .A(round_inst_sin_w[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n461) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n391), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n394) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n451), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n390), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U24 ( .A1(
        round_inst_sin_y[42]), .A2(round_inst_sin_w[41]), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n390) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U23 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_z[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n451) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U22 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n409), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n389), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n396) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U21 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n446), .Z(
        round_inst_S_10__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U20 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n388), .A2(round_inst_sin_y[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n446) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_10__sbox_inst_n1), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n388) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n387), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n386), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n515) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U17 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n385), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n419), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n386) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U16 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_z[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n419) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U15 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n384), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n385) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U14 ( .A(round_inst_sin_w[41]), .B(round_inst_S_10__sbox_inst_com_x_inst_n383), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n384) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_10__sbox_inst_n1), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_10__sbox_inst_com_x_inst_U12 ( .A(round_inst_sin_z[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n409) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n382), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n387) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_x_inst_U10 ( .A1(
        round_inst_sin_z[40]), .A2(round_inst_sin_y[43]), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n415) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U9 ( .A1(
        round_inst_S_10__sbox_inst_com_x_inst_n381), .A2(
        round_inst_S_10__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n382) );
  INV_X1 round_inst_S_10__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_y[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n462) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U7 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n507), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n380), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n381) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_x_inst_U6 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_10__sbox_inst_com_x_inst_n475), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n380) );
  INV_X1 round_inst_S_10__sbox_inst_com_x_inst_U5 ( .A(round_inst_sin_y[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n475) );
  INV_X1 round_inst_S_10__sbox_inst_com_x_inst_U4 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n476) );
  INV_X1 round_inst_S_10__sbox_inst_com_x_inst_U3 ( .A(round_inst_sin_y[41]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n408) );
  INV_X1 round_inst_S_10__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_10__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_10__sbox_inst_com_x_inst_n507) );
  INV_X1 round_inst_S_10__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_w[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_x_inst_n490) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n516), .Z(round_inst_sout_y[40])
         );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n515), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U134 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n513), .B(round_inst_sin_z[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n514) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U133 ( .A(round_inst_sin_x[36]), .B(round_inst_S_10__sbox_inst_com_y_inst_n512), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n515) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n511), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_srout2_y[26]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n507), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n517) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U129 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n506), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n505), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n507) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n505) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U127 ( .A1(
        round_inst_sin_w[42]), .A2(round_inst_sin_z[43]), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n506) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U125 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_10__sbox_inst_com_y_inst_U124 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_10__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U123 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_sin_x[43]), .A2(round_inst_S_10__sbox_inst_com_y_inst_n493), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U121 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n492), .A2(round_inst_sin_z[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U120 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U119 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U118 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U117 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n486), .A2(round_inst_sin_z[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U116 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_sin_w[42]), .A2(round_inst_sin_w[40]), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U114 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n513), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U112 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U111 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_10__sbox_inst_n1), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U109 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[39]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_y_inst_U108 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n513), .A2(round_inst_sin_z[43]), 
        .A3(round_inst_sin_x[40]), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U107 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_sin_w[40]), .A2(round_inst_sin_w[43]), .A3(
        round_inst_S_10__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_10__sbox_inst_com_y_inst_U105 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_10__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U104 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[24]) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U103 ( .A1(
        round_inst_S_10__sbox_inst_n5), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n508) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U98 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U97 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_10__sbox_inst_n1), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_10__sbox_inst_com_y_inst_U95 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U94 ( .A1(
        round_inst_sin_x[40]), .A2(round_inst_sin_w[42]), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_y_inst_U93 ( .A1(
        round_inst_sin_w[40]), .A2(round_inst_S_10__sbox_inst_n3), .A3(
        round_inst_S_10__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U92 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U91 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U88 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U87 ( .A1(
        round_inst_S_10__sbox_inst_n1), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_10__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_10__sbox_inst_n5), .B(round_inst_sin_w[42]), .S(
        round_inst_S_10__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U84 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U80 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_10__sbox_inst_n1), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U78 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n478), .B(round_inst_sin_x[37]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_sin_w[42]), .A2(round_inst_S_10__sbox_inst_com_y_inst_n483), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U76 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n513), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n438), .Z(
        round_inst_srout2_y[27]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U71 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U70 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U69 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n483), .A2(
        round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_10__sbox_inst_n1), .A2(round_inst_sin_w[40]), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_y_inst_U66 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[43]), 
        .A3(round_inst_S_10__sbox_inst_n1), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U65 ( .A(round_inst_sin_w[40]), 
        .B(round_inst_sin_x[40]), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U63 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U61 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U59 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U58 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U57 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[41]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U55 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_10__sbox_inst_com_y_inst_U54 ( .A(round_inst_sin_x[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U53 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n418), .A2(round_inst_sin_z[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U51 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U50 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U49 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n414), .B(
        round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U48 ( .A(round_inst_sin_w[41]), .B(round_inst_S_10__sbox_inst_n1), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_10__sbox_inst_n1), .A2(round_inst_sin_x[40]), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U46 ( .A1(
        round_inst_S_10__sbox_inst_n1), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U45 ( .A(round_inst_sin_x[38]), 
        .B(round_inst_S_10__sbox_inst_com_y_inst_n512), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U44 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n512) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U43 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U42 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U41 ( .A(round_inst_sin_w[41]), 
        .B(round_inst_sin_x[43]), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U40 ( .A(
        round_inst_S_10__sbox_inst_n3), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_10__sbox_inst_com_y_inst_U39 ( .A(round_inst_sin_w[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U38 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[40]), 
        .Z(round_inst_S_10__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_10__sbox_inst_com_y_inst_U36 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_10__sbox_inst_com_y_inst_U35 ( .A(round_inst_sin_z[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_10__sbox_inst_n1), .B(round_inst_sin_z[43]), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U30 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U29 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_10__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U27 ( .A(
        round_inst_S_10__sbox_inst_n5), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_sin_w[41]), .A2(round_inst_sin_z[43]), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n513), .A2(round_inst_sin_w[41]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_10__sbox_inst_n1), .A2(round_inst_sin_w[43]), .A3(
        round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U22 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_10__sbox_inst_n1), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U21 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U20 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n397) );
  INV_X1 round_inst_S_10__sbox_inst_com_y_inst_U19 ( .A(round_inst_sin_w[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n396) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n503), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U17 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_z[43]), .B(round_inst_sin_w[43]), .ZN(round_inst_S_10__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U15 ( .A(round_inst_sin_z[43]), 
        .B(round_inst_S_10__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n503) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U14 ( .A(round_inst_sin_w[43]), .B(round_inst_sin_x[43]), .ZN(round_inst_S_10__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U13 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U12 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_y_inst_U11 ( .A1(
        round_inst_S_10__sbox_inst_n3), .A2(round_inst_sin_w[43]), .A3(
        round_inst_S_10__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_y_inst_U10 ( .A1(
        round_inst_sin_z[43]), .A2(round_inst_S_10__sbox_inst_com_y_inst_n389), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_10__sbox_inst_com_y_inst_U9 ( .A(round_inst_sin_w[41]), 
        .B(round_inst_S_10__sbox_inst_n3), .S(round_inst_sin_w[42]), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_10__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_10__sbox_inst_n3), .A2(
        round_inst_S_10__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_10__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U6 ( .A(round_inst_sin_z[43]), 
        .B(round_inst_sin_x[43]), .Z(
        round_inst_S_10__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_y_inst_U5 ( .A1(
        round_inst_S_10__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_10__sbox_inst_n1), .A3(round_inst_sin_x[43]), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_10__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_y_inst_U3 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n513), .B(round_inst_sin_w[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_10__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_10__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_10__sbox_inst_com_y_inst_n513) );
  INV_X1 round_inst_S_10__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U137 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n523), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n522), .ZN(round_inst_sout_z[40]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U136 ( .A(
        round_inst_sin_w[43]), .B(round_inst_S_10__sbox_inst_com_z_inst_n521), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n522) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U135 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n520), .B(round_inst_sin_w[42]), 
        .Z(round_inst_S_10__sbox_inst_com_z_inst_n523) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U134 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n519), .B(round_inst_sin_x[36]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n520) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U133 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n518), .B(round_inst_n54), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n519) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U132 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n517), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n516), .Z(
        round_inst_srout2_z[26]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n515), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n514), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n516) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n512), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n514) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U129 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n511), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n510), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n512) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U128 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n509), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n508), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n518), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n507), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n511) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n506), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n505), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_sin_w[41]), .B(round_inst_sin_x[39]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n505) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U124 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n504), .B(round_inst_sin_y[39]), 
        .Z(round_inst_S_10__sbox_inst_com_z_inst_n506) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U123 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n503), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n502), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n504) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U122 ( .A1(
        round_inst_sin_y[40]), .A2(round_inst_S_10__sbox_inst_com_z_inst_n501), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n502) );
  INV_X1 round_inst_S_10__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n500), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n501) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U120 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n499), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n498), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n503) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_z_inst_U119 ( .A1(
        round_inst_sin_x[40]), .A2(round_inst_sin_w[43]), .A3(
        round_inst_S_10__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n498) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U118 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n496), .B(
        round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n497) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U117 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n495), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n494), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n499) );
  INV_X1 round_inst_S_10__sbox_inst_com_z_inst_U116 ( .A(round_inst_sin_x[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n494) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U115 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n500), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n518) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U114 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n491), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n493) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U113 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n508), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n490), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n491) );
  INV_X1 round_inst_S_10__sbox_inst_com_z_inst_U112 ( .A(round_inst_sin_w[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n490) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U111 ( .A1(
        round_inst_sin_w[42]), .A2(round_inst_S_10__sbox_inst_com_z_inst_n489), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n513) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U110 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n488), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n508), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n488) );
  INV_X1 round_inst_S_10__sbox_inst_com_z_inst_U108 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n486) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U107 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n484), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U106 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n482), .ZN(
        round_inst_srout2_z[24]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n481), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n482) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U104 ( .A1(
        round_inst_sin_w[40]), .A2(round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n495) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n509), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n479), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n478), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n480) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U101 ( .A1(
        round_inst_sin_w[42]), .A2(round_inst_S_10__sbox_inst_com_z_inst_n485), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n478) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U100 ( .A(round_inst_sin_y[37]), .B(round_inst_sin_x[37]), .Z(round_inst_S_10__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U99 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n492), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n483) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U98 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n476), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n492) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U97 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n474), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n475) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U96 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n472), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n471), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U95 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n470), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n471) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U94 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n468), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n469) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n467), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n466), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n470) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n465), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n464), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n466) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U91 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n463), .A2(round_inst_sin_w[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n464) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U90 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n462), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U89 ( .A1(
        round_inst_S_10__sbox_inst_n3), .A2(round_inst_sin_y[40]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n462) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U88 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n461), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n460), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U87 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n459), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n458), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n460) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n458) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U85 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n455), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n459) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U84 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n453), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n509), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U83 ( .A1(
        round_inst_sin_w[40]), .A2(round_inst_sin_y[42]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n509) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_sin_w[42]), .A2(round_inst_sin_x[40]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U81 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n452), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n461) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U80 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n450), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U79 ( .A(
        round_inst_S_10__sbox_inst_n5), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n449) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U78 ( .A(round_inst_sin_y[42]), 
        .B(round_inst_sin_w[42]), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n448) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n452), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U76 ( .A(round_inst_sin_w[42]), .B(round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n452) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U75 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n446), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_srout2_z[27]) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n445) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U73 ( .A(round_inst_sin_w[40]), .B(round_inst_S_10__sbox_inst_com_z_inst_n477), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U72 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n477) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U71 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n440), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n441) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U70 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n457), .A2(round_inst_sin_w[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n439) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U69 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n474), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n457) );
  AND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U68 ( .A1(round_inst_sin_w[41]), .A2(round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n474) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n437), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n436), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U66 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n435), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n434), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n436) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U65 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n456), .A2(round_inst_sin_y[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n434) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U64 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n433), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n432), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n456) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U63 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n431), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n430), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U62 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n429), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n428), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n430) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_z_inst_U61 ( .A1(
        round_inst_S_10__sbox_inst_n3), .A2(round_inst_sin_w[43]), .A3(
        round_inst_S_10__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n428) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U60 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n427), .A2(round_inst_sin_w[41]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n429) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U59 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n426), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n425), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n427) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U58 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n424), .A2(
        round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U57 ( .A(round_inst_sin_x[43]), 
        .B(round_inst_sin_y[43]), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n424) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U56 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n422), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U55 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U54 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n419), .A2(round_inst_sin_w[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n420) );
  INV_X1 round_inst_S_10__sbox_inst_com_z_inst_U53 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n419) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U52 ( .A1(
        round_inst_sin_y[43]), .A2(round_inst_S_10__sbox_inst_com_z_inst_n438), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n421) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U51 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n418), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n500), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n423) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U50 ( .A1(
        round_inst_sin_w[43]), .A2(round_inst_S_10__sbox_inst_n5), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n500) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U49 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n417), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n432), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n437) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U48 ( .A1(
        round_inst_sin_w[41]), .A2(round_inst_sin_w[42]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n432) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U47 ( .A(round_inst_sin_x[43]), .B(round_inst_sin_w[43]), .ZN(round_inst_S_10__sbox_inst_com_z_inst_n417) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U46 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n416), .A2(round_inst_sin_x[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n442) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U45 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U44 ( .A(round_inst_sin_w[41]), .B(round_inst_S_10__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n414) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U43 ( .A1(
        round_inst_S_10__sbox_inst_n3), .A2(round_inst_sin_w[42]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n433) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n413), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n415) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U41 ( .A1(
        round_inst_sin_y[41]), .A2(round_inst_sin_w[42]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n413) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U40 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n412), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n438) );
  INV_X1 round_inst_S_10__sbox_inst_com_z_inst_U39 ( .A(round_inst_sin_y[42]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n496) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U38 ( .A(round_inst_n55), .B(
        round_inst_sin_x[38]), .Z(round_inst_S_10__sbox_inst_com_z_inst_n444)
         );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n521), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n517), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n411), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n410), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n517) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U35 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n409), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n408), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n410) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U34 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n407), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n406), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n408) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n405), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n406) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U32 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n403), .A2(round_inst_sin_y[43]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n404) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n402), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n401), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n405) );
  MUX2_X1 round_inst_S_10__sbox_inst_com_z_inst_U30 ( .A(round_inst_sin_x[43]), 
        .B(round_inst_sin_w[43]), .S(
        round_inst_S_10__sbox_inst_com_z_inst_n400), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n401) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_sin_w[41]), .A2(round_inst_S_10__sbox_inst_com_z_inst_n485), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n400) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U28 ( .A(round_inst_sin_w[40]), 
        .B(round_inst_sin_x[40]), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n485) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_z_inst_U27 ( .A1(
        round_inst_sin_w[43]), .A2(round_inst_S_10__sbox_inst_n3), .A3(
        round_inst_S_10__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n402) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U26 ( .A(round_inst_sin_w[40]), 
        .B(round_inst_sin_y[40]), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n473) );
  NAND3_X1 round_inst_S_10__sbox_inst_com_z_inst_U25 ( .A1(
        round_inst_sin_w[40]), .A2(round_inst_sin_x[43]), .A3(
        round_inst_S_10__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n407) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U24 ( .A(
        round_inst_S_10__sbox_inst_n3), .B(round_inst_sin_y[41]), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n454) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U23 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n484), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n409) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_sin_w[40]), .A2(round_inst_sin_y[41]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n447) );
  INV_X1 round_inst_S_10__sbox_inst_com_z_inst_U21 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n425), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n484) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U20 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n399), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n398), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n411) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U19 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n418), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n398) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U18 ( .A(round_inst_sin_y[41]), .B(round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n418) );
  NOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U17 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_10__sbox_inst_com_z_inst_n412), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n399) );
  INV_X1 round_inst_S_10__sbox_inst_com_z_inst_U16 ( .A(round_inst_sin_w[41]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n412) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U15 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n395), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U14 ( .A1(
        round_inst_sin_x[43]), .A2(round_inst_sin_y[40]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n487) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U13 ( .A1(
        round_inst_sin_y[43]), .A2(round_inst_sin_x[40]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n395) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U12 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n394), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n393), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n521) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U11 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n392), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U10 ( .A1(
        round_inst_sin_x[40]), .A2(round_inst_sin_w[41]), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n450) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U9 ( .A1(
        round_inst_S_10__sbox_inst_com_z_inst_n391), .A2(round_inst_sin_w[40]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n392) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U8 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n508), .B(round_inst_sin_y[41]), 
        .ZN(round_inst_S_10__sbox_inst_com_z_inst_n391) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U7 ( .A(round_inst_sin_x[43]), 
        .B(round_inst_S_10__sbox_inst_com_z_inst_n425), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n508) );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U6 ( .A(round_inst_sin_w[43]), 
        .B(round_inst_sin_y[43]), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n425) );
  XNOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U5 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n394) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U4 ( .A1(round_inst_sin_w[43]), .A2(round_inst_sin_x[40]), .ZN(round_inst_S_10__sbox_inst_com_z_inst_n397)
         );
  XOR2_X1 round_inst_S_10__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_10__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_10__sbox_inst_com_z_inst_n451), .Z(
        round_inst_S_10__sbox_inst_com_z_inst_n403) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U2 ( .A1(round_inst_sin_w[40]), .A2(round_inst_S_10__sbox_inst_n3), .ZN(
        round_inst_S_10__sbox_inst_com_z_inst_n451) );
  NAND2_X1 round_inst_S_10__sbox_inst_com_z_inst_U1 ( .A1(round_inst_sin_w[40]), .A2(round_inst_sin_w[41]), .ZN(round_inst_S_10__sbox_inst_com_z_inst_n468)
         );
  INV_X1 round_inst_S_11__sbox_inst_U6 ( .A(round_inst_sin_x[45]), .ZN(
        round_inst_S_11__sbox_inst_n4) );
  INV_X1 round_inst_S_11__sbox_inst_U5 ( .A(round_inst_sin_x[46]), .ZN(
        round_inst_S_11__sbox_inst_n6) );
  INV_X1 round_inst_S_11__sbox_inst_U4 ( .A(round_inst_sin_z[45]), .ZN(
        round_inst_S_11__sbox_inst_n2) );
  INV_X2 round_inst_S_11__sbox_inst_U3 ( .A(round_inst_S_11__sbox_inst_n6), 
        .ZN(round_inst_S_11__sbox_inst_n5) );
  INV_X2 round_inst_S_11__sbox_inst_U2 ( .A(round_inst_S_11__sbox_inst_n2), 
        .ZN(round_inst_S_11__sbox_inst_n1) );
  INV_X2 round_inst_S_11__sbox_inst_U1 ( .A(round_inst_S_11__sbox_inst_n4), 
        .ZN(round_inst_S_11__sbox_inst_n3) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n531), .ZN(round_inst_sout_w[47]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U139 ( .A1(
        round_inst_sin_z[44]), .A2(round_inst_S_11__sbox_inst_com_w_inst_n528), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n526), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n524), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n526) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[46]), .A2(round_inst_S_11__sbox_inst_com_w_inst_n523), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n525) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n518), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n516), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n518) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n514), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n513), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n512), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n513) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_w_inst_U128 ( .A1(
        round_inst_S_11__sbox_inst_n5), .A2(round_inst_sin_x[44]), .A3(
        round_inst_S_11__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n511) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U127 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n509), .A2(round_inst_sin_y[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n508), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n507), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U125 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n508) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_sin_z[47]), .A2(round_inst_S_11__sbox_inst_com_w_inst_n504), 
        .A3(round_inst_sin_x[44]), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U122 ( .A(
        round_inst_sin_y[43]), .B(round_inst_S_11__sbox_inst_com_w_inst_n501), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U121 ( .A(
        round_inst_S_11__sbox_inst_n3), .B(round_inst_sin_z[43]), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n501) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U120 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[45]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[41]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[41]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U113 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[44]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_11__sbox_inst_n5), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U110 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n528), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U105 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_11__sbox_inst_n5), .B(round_inst_sin_z[46]), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_11__sbox_inst_n1), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U99 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n504), .A2(round_inst_sin_x[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_11__sbox_inst_n5), .A2(round_inst_sin_y[44]), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n507) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U94 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n461), .A2(
        round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U88 ( .A1(round_inst_sin_z[44]), .A2(round_inst_S_11__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_w_inst_U85 ( .A1(
        round_inst_sin_y[45]), .A2(round_inst_sin_y[44]), .A3(
        round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_w_inst_U84 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_11__sbox_inst_n3), .A3(round_inst_sin_y[44]), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n528) );
  OR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_11__sbox_inst_n5), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U80 ( .A(round_inst_sin_y[40]), 
        .B(round_inst_sin_z[40]), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n484) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U79 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[47])
         );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U73 ( .A1(
        round_inst_sin_z[47]), .A2(round_inst_S_11__sbox_inst_com_w_inst_n440), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U71 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n504), .A2(
        round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_11__sbox_inst_n5), .A2(round_inst_sin_y[45]), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U69 ( .A1(
        round_inst_S_11__sbox_inst_n1), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_11__sbox_inst_n5), .A2(round_inst_S_11__sbox_inst_n1), 
        .A3(round_inst_S_11__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n439), .A2(
        round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n505), .A2(
        round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U63 ( .A(round_inst_sin_z[47]), 
        .B(round_inst_S_11__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n505) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U62 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U61 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U60 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U58 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U57 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U56 ( .A(round_inst_sin_y[45]), .B(round_inst_S_11__sbox_inst_n1), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U55 ( .A1(
        round_inst_sin_z[47]), .A2(round_inst_S_11__sbox_inst_n1), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U54 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_w_inst_U52 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n506), .A3(
        round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U51 ( .A(round_inst_sin_y[45]), 
        .B(round_inst_S_11__sbox_inst_n3), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_w_inst_U50 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n506), .A2(round_inst_sin_y[45]), 
        .A3(round_inst_S_11__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U49 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n504), .B(round_inst_sin_z[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n465) );
  INV_X1 round_inst_S_11__sbox_inst_com_w_inst_U48 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n436), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n504) );
  INV_X1 round_inst_S_11__sbox_inst_com_w_inst_U47 ( .A(round_inst_sin_y[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U45 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n520) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U44 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n421), .A2(round_inst_sin_z[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U43 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U42 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n419), .A2(
        round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U40 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_11__sbox_inst_n1), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U38 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n521) );
  INV_X1 round_inst_S_11__sbox_inst_com_w_inst_U37 ( .A(round_inst_sin_x[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n489) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U36 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U33 ( .A(round_inst_sin_x[44]), .B(round_inst_sin_z[44]), .ZN(round_inst_S_11__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U32 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n498), .A2(
        round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U31 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U30 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U29 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U28 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U27 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U26 ( .A1(
        round_inst_S_11__sbox_inst_n3), .A2(round_inst_sin_z[44]), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n522), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U24 ( .A(
        round_inst_S_11__sbox_inst_n3), .B(round_inst_S_11__sbox_inst_n1), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_11__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U22 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U21 ( .A1(
        round_inst_sin_x[44]), .A2(round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U20 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[45]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U19 ( .A(round_inst_sin_y[44]), 
        .B(round_inst_sin_z[44]), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n418) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U17 ( .A(round_inst_sin_x[44]), .B(round_inst_S_11__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U15 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n398), .A2(round_inst_sin_x[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U13 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n498), .B(
        round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_11__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_11__sbox_inst_com_w_inst_U11 ( .A(round_inst_sin_y[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_11__sbox_inst_n1), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U9 ( .A(round_inst_sin_z[47]), 
        .B(round_inst_S_11__sbox_inst_com_w_inst_n506), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n510) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U8 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U7 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_11__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U6 ( .A1(
        round_inst_S_11__sbox_inst_n3), .A2(round_inst_sin_y[44]), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U5 ( .A1(round_inst_sin_x[44]), .A2(round_inst_sin_y[45]), .ZN(round_inst_S_11__sbox_inst_com_w_inst_n477)
         );
  NAND2_X1 round_inst_S_11__sbox_inst_com_w_inst_U4 ( .A1(
        round_inst_S_11__sbox_inst_com_w_inst_n506), .A2(round_inst_sin_y[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n522) );
  INV_X1 round_inst_S_11__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_11__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_11__sbox_inst_com_w_inst_n506) );
  INV_X1 round_inst_S_11__sbox_inst_com_w_inst_U2 ( .A(round_inst_sin_x[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_w_inst_n486) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_w_inst_U1 ( .A(round_inst_sin_y[42]), 
        .B(round_inst_sin_z[42]), .Z(
        round_inst_S_11__sbox_inst_com_w_inst_n402) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U144 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n519), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n518), .Z(round_inst_sout_x[44])
         );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U143 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n517), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n516), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n518) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U142 ( .A(
        round_inst_sin_y[46]), .B(round_inst_sin_y[47]), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n516) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U141 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n515), .B(round_inst_sin_z[40]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n517) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U140 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n514), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n513), .ZN(
        round_inst_srout2_x[46]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U139 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n512), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n511), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n513) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U138 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n510), .A2(round_inst_sin_z[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n511) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U137 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n509), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n510) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U136 ( .A1(
        round_inst_sin_y[46]), .A2(round_inst_S_11__sbox_inst_com_x_inst_n507), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n508) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n506), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n505), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n512) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n504), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n503), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n505) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U133 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n509), .A2(round_inst_sin_w[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U132 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n501), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n504) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n501) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_x_inst_U130 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n497), .A3(round_inst_sin_y[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n499) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U129 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n496), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n495), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n500) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_x_inst_U128 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n494), .A2(round_inst_sin_y[44]), 
        .A3(round_inst_sin_y[46]), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n495) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U127 ( .A(round_inst_sin_y[47]), .B(round_inst_sin_z[47]), .Z(round_inst_S_11__sbox_inst_com_x_inst_n494) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U126 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n493), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n496) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_x_inst_U125 ( .A1(
        round_inst_sin_y[46]), .A2(round_inst_sin_z[44]), .A3(
        round_inst_sin_z[47]), .ZN(round_inst_S_11__sbox_inst_com_x_inst_n502)
         );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U124 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n492), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n506) );
  OR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U123 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n493), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n491) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U122 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U121 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n488) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n484), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n486) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n483), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n484) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U118 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n507), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n482) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U117 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n480), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n479), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n483) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U116 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n478), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n479) );
  AND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U115 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n481), .A2(round_inst_sin_z[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n477) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U114 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .B(round_inst_sin_z[43]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n478) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_x_inst_U113 ( .A1(
        round_inst_sin_y[46]), .A2(round_inst_sin_w[44]), .A3(
        round_inst_sin_z[47]), .ZN(round_inst_S_11__sbox_inst_com_x_inst_n480)
         );
  NAND3_X1 round_inst_S_11__sbox_inst_com_x_inst_U112 ( .A1(
        round_inst_sin_y[46]), .A2(round_inst_sin_y[44]), .A3(
        round_inst_S_11__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U111 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n475), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n493), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n487) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_y[46]), .A2(round_inst_sin_z[44]), .A3(
        round_inst_sin_y[47]), .ZN(round_inst_S_11__sbox_inst_com_x_inst_n489)
         );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n519), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n474), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n514) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U108 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n473), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n519) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n471), .A2(round_inst_sin_y[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n472) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_sin_z[47]), .B(round_inst_S_11__sbox_inst_com_x_inst_n470), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n471) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U105 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n509), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n473) );
  AND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U104 ( .A1(
        round_inst_sin_z[46]), .A2(round_inst_sin_y[47]), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n509) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n468), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n467), .ZN(
        round_inst_srout2_x[44]) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n493), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n467) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U101 ( .A1(
        round_inst_sin_y[44]), .A2(round_inst_sin_z[46]), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n493) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U100 ( .A1(
        round_inst_sin_y[46]), .A2(round_inst_S_11__sbox_inst_com_x_inst_n498), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n466) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U99 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n465), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n468) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n463), .B(round_inst_sin_z[41]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n464) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n463) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U96 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n462), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n481) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U95 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n460), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n459), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n469) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U94 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n458), .A2(round_inst_sin_y[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n459) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n457), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n458) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_11__sbox_inst_n1), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n498), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n455), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n454), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n460) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U90 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n453), .A2(round_inst_sin_w[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n454) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n451), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n453) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_sin_y[46]), .A2(round_inst_S_11__sbox_inst_n1), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n452) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n450), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n449), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n455) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U86 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n448), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n447), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n449) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U85 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n446), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n445), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n447) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n443), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n445) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n497), .B(round_inst_sin_z[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n443) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U82 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n442), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n441), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n440), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n448) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U80 ( .A1(
        round_inst_sin_y[46]), .A2(round_inst_sin_z[44]), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n441) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_x_inst_U79 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n498), .A3(
        round_inst_S_11__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U78 ( .A(round_inst_sin_z[46]), 
        .B(round_inst_S_11__sbox_inst_com_x_inst_n497), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n439) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U77 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n515), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_srout2_x[47]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U76 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n437), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n436), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U75 ( .A(round_inst_sin_y[44]), .B(round_inst_S_11__sbox_inst_com_x_inst_n474), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n436) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U74 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n435), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n434), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n433), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n432), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n434) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U72 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n431), .A2(round_inst_sin_w[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n432) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U71 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n430), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n429), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n431) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U70 ( .A1(
        round_inst_S_11__sbox_inst_n1), .A2(round_inst_sin_y[47]), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n429) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U69 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_z[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n428), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n433) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U67 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n426), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n427) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n424), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n423), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n422), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n421), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n423) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U64 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n507), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n421) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U63 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n440), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n456) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .B(round_inst_sin_w[45]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n440) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U61 ( .A1(
        round_inst_sin_z[47]), .A2(round_inst_S_11__sbox_inst_com_x_inst_n442), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n422) );
  AND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U60 ( .A1(round_inst_sin_y[44]), .A2(round_inst_S_11__sbox_inst_com_x_inst_n420), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n442) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_x_inst_U59 ( .A1(
        round_inst_sin_w[45]), .A2(round_inst_S_11__sbox_inst_com_x_inst_n498), 
        .A3(round_inst_sin_y[47]), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U58 ( .A(round_inst_sin_z[44]), 
        .B(round_inst_sin_y[44]), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n498) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U57 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n419), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n426) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_11__sbox_inst_n1), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n416), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n417) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n470), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n416) );
  MUX2_X1 round_inst_S_11__sbox_inst_com_x_inst_U53 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n419), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n414), .S(
        round_inst_S_11__sbox_inst_com_x_inst_n413), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n435) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U52 ( .A1(
        round_inst_sin_y[47]), .A2(round_inst_S_11__sbox_inst_com_x_inst_n412), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n413) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_y[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n412) );
  MUX2_X1 round_inst_S_11__sbox_inst_com_x_inst_U50 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n411), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n410), .S(
        round_inst_S_11__sbox_inst_com_x_inst_n409), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n414) );
  NOR3_X1 round_inst_S_11__sbox_inst_com_x_inst_U49 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n410), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n462), .A3(
        round_inst_S_11__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n411) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n475), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n419), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n410) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U47 ( .A(round_inst_sin_z[42]), 
        .B(round_inst_S_11__sbox_inst_com_x_inst_n465), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n407), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n406), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n465) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U45 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n405), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n406) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n405) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U43 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n418), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n404) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U42 ( .A(round_inst_sin_z[47]), .B(round_inst_S_11__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n418) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U41 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n403), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n402), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n407) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_x_inst_U40 ( .A1(
        round_inst_sin_z[46]), .A2(round_inst_sin_y[47]), .A3(
        round_inst_S_11__sbox_inst_com_x_inst_n401), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n402) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U39 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n420), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n401) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U38 ( .A(
        round_inst_S_11__sbox_inst_n1), .B(round_inst_sin_w[45]), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n420) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U37 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n400), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n399), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n403) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U36 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n446), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n399) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U35 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n475), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n398), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n397), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n400) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U33 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n490), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n451), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n397) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U32 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n396), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n395), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U31 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n395) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U30 ( .A1(
        round_inst_sin_y[47]), .A2(round_inst_S_11__sbox_inst_com_x_inst_n392), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n393) );
  MUX2_X1 round_inst_S_11__sbox_inst_com_x_inst_U29 ( .A(
        round_inst_S_11__sbox_inst_n1), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .S(
        round_inst_S_11__sbox_inst_com_x_inst_n497), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n392) );
  INV_X1 round_inst_S_11__sbox_inst_com_x_inst_U28 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n497) );
  INV_X1 round_inst_S_11__sbox_inst_com_x_inst_U27 ( .A(round_inst_sin_w[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n461) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n391), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n394) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n451), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n390), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U24 ( .A1(
        round_inst_sin_y[46]), .A2(round_inst_sin_w[45]), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n390) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U23 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_z[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n451) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U22 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n409), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n389), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n396) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U21 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n446), .Z(
        round_inst_S_11__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U20 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n388), .A2(round_inst_sin_y[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n446) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_11__sbox_inst_n1), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n388) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n387), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n386), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n515) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U17 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n385), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n419), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n386) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U16 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_z[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n419) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U15 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n384), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n385) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U14 ( .A(round_inst_sin_w[45]), .B(round_inst_S_11__sbox_inst_com_x_inst_n383), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n384) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_11__sbox_inst_n1), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_11__sbox_inst_com_x_inst_U12 ( .A(round_inst_sin_z[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n409) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n382), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n387) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_x_inst_U10 ( .A1(
        round_inst_sin_z[44]), .A2(round_inst_sin_y[47]), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n415) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U9 ( .A1(
        round_inst_S_11__sbox_inst_com_x_inst_n381), .A2(
        round_inst_S_11__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n382) );
  INV_X1 round_inst_S_11__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_y[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n462) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U7 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n507), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n380), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n381) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_x_inst_U6 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_11__sbox_inst_com_x_inst_n475), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n380) );
  INV_X1 round_inst_S_11__sbox_inst_com_x_inst_U5 ( .A(round_inst_sin_y[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n475) );
  INV_X1 round_inst_S_11__sbox_inst_com_x_inst_U4 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n476) );
  INV_X1 round_inst_S_11__sbox_inst_com_x_inst_U3 ( .A(round_inst_sin_y[45]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n408) );
  INV_X1 round_inst_S_11__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_11__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_11__sbox_inst_com_x_inst_n507) );
  INV_X1 round_inst_S_11__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_w[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_x_inst_n490) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n516), .Z(round_inst_sout_y[44])
         );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n515), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U134 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n513), .B(round_inst_sin_z[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n514) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U133 ( .A(round_inst_sin_x[40]), .B(round_inst_S_11__sbox_inst_com_y_inst_n512), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n515) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n511), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_srout2_y[46]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n507), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n517) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U129 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n506), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n505), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n507) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n505) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U127 ( .A1(
        round_inst_sin_w[46]), .A2(round_inst_sin_z[47]), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n506) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U125 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_11__sbox_inst_com_y_inst_U124 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_11__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U123 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_sin_x[47]), .A2(round_inst_S_11__sbox_inst_com_y_inst_n493), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U121 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n492), .A2(round_inst_sin_z[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U120 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U119 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U118 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U117 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n486), .A2(round_inst_sin_z[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U116 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_sin_w[46]), .A2(round_inst_sin_w[44]), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U114 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n513), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U112 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U111 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_11__sbox_inst_n1), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U109 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[43]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_y_inst_U108 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n513), .A2(round_inst_sin_z[47]), 
        .A3(round_inst_sin_x[44]), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U107 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_sin_w[44]), .A2(round_inst_sin_w[47]), .A3(
        round_inst_S_11__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_11__sbox_inst_com_y_inst_U105 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_11__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U104 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[44]) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U103 ( .A1(
        round_inst_S_11__sbox_inst_n5), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n508) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U98 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U97 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_11__sbox_inst_n1), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_11__sbox_inst_com_y_inst_U95 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U94 ( .A1(
        round_inst_sin_x[44]), .A2(round_inst_sin_w[46]), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_y_inst_U93 ( .A1(
        round_inst_sin_w[44]), .A2(round_inst_S_11__sbox_inst_n3), .A3(
        round_inst_S_11__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U92 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U91 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U88 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U87 ( .A1(
        round_inst_S_11__sbox_inst_n1), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_11__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_11__sbox_inst_n5), .B(round_inst_sin_w[46]), .S(
        round_inst_S_11__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U84 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U80 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_11__sbox_inst_n1), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U78 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n478), .B(round_inst_sin_x[41]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_sin_w[46]), .A2(round_inst_S_11__sbox_inst_com_y_inst_n483), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U76 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n513), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n438), .Z(
        round_inst_srout2_y[47]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U71 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U70 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U69 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n483), .A2(
        round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_11__sbox_inst_n1), .A2(round_inst_sin_w[44]), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_y_inst_U66 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[47]), 
        .A3(round_inst_S_11__sbox_inst_n1), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U65 ( .A(round_inst_sin_w[44]), 
        .B(round_inst_sin_x[44]), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U63 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U61 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U59 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U58 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U57 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[45]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U55 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_11__sbox_inst_com_y_inst_U54 ( .A(round_inst_sin_x[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U53 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n418), .A2(round_inst_sin_z[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U51 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U50 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U49 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n414), .B(
        round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U48 ( .A(round_inst_sin_w[45]), .B(round_inst_S_11__sbox_inst_n1), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_11__sbox_inst_n1), .A2(round_inst_sin_x[44]), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U46 ( .A1(
        round_inst_S_11__sbox_inst_n1), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U45 ( .A(round_inst_sin_x[42]), 
        .B(round_inst_S_11__sbox_inst_com_y_inst_n512), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U44 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n512) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U43 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U42 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U41 ( .A(round_inst_sin_w[45]), 
        .B(round_inst_sin_x[47]), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U40 ( .A(
        round_inst_S_11__sbox_inst_n3), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_11__sbox_inst_com_y_inst_U39 ( .A(round_inst_sin_w[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U38 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[44]), 
        .Z(round_inst_S_11__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_11__sbox_inst_com_y_inst_U36 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_11__sbox_inst_com_y_inst_U35 ( .A(round_inst_sin_z[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_11__sbox_inst_n1), .B(round_inst_sin_z[47]), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U30 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U29 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_11__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U27 ( .A(
        round_inst_S_11__sbox_inst_n5), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_sin_w[45]), .A2(round_inst_sin_z[47]), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n513), .A2(round_inst_sin_w[45]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_11__sbox_inst_n1), .A2(round_inst_sin_w[47]), .A3(
        round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U22 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_11__sbox_inst_n1), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U21 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U20 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n397) );
  INV_X1 round_inst_S_11__sbox_inst_com_y_inst_U19 ( .A(round_inst_sin_w[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n396) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n503), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U17 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_z[47]), .B(round_inst_sin_w[47]), .ZN(round_inst_S_11__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U15 ( .A(round_inst_sin_z[47]), 
        .B(round_inst_S_11__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n503) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U14 ( .A(round_inst_sin_w[47]), .B(round_inst_sin_x[47]), .ZN(round_inst_S_11__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U13 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U12 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_y_inst_U11 ( .A1(
        round_inst_S_11__sbox_inst_n3), .A2(round_inst_sin_w[47]), .A3(
        round_inst_S_11__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_y_inst_U10 ( .A1(
        round_inst_sin_z[47]), .A2(round_inst_S_11__sbox_inst_com_y_inst_n389), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_11__sbox_inst_com_y_inst_U9 ( .A(round_inst_sin_w[45]), 
        .B(round_inst_S_11__sbox_inst_n3), .S(round_inst_sin_w[46]), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_11__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_11__sbox_inst_n3), .A2(
        round_inst_S_11__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_11__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U6 ( .A(round_inst_sin_z[47]), 
        .B(round_inst_sin_x[47]), .Z(
        round_inst_S_11__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_y_inst_U5 ( .A1(
        round_inst_S_11__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_11__sbox_inst_n1), .A3(round_inst_sin_x[47]), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_11__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_y_inst_U3 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n513), .B(round_inst_sin_w[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_11__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_11__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_11__sbox_inst_com_y_inst_n513) );
  INV_X1 round_inst_S_11__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U137 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n523), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n522), .ZN(round_inst_sout_z[44]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U136 ( .A(
        round_inst_sin_w[47]), .B(round_inst_S_11__sbox_inst_com_z_inst_n521), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n522) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U135 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n520), .B(round_inst_sin_w[46]), 
        .Z(round_inst_S_11__sbox_inst_com_z_inst_n523) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U134 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n519), .B(round_inst_sin_x[40]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n520) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U133 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n518), .B(round_inst_sin_y[40]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n519) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U132 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n517), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n516), .Z(
        round_inst_srout2_z[46]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n515), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n514), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n516) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n512), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n514) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U129 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n511), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n510), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n512) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U128 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n509), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n508), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n518), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n507), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n511) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n506), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n505), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_sin_w[45]), .B(round_inst_sin_x[43]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n505) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U124 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n504), .B(round_inst_sin_y[43]), 
        .Z(round_inst_S_11__sbox_inst_com_z_inst_n506) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U123 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n503), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n502), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n504) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U122 ( .A1(
        round_inst_sin_y[44]), .A2(round_inst_S_11__sbox_inst_com_z_inst_n501), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n502) );
  INV_X1 round_inst_S_11__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n500), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n501) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U120 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n499), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n498), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n503) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_z_inst_U119 ( .A1(
        round_inst_sin_x[44]), .A2(round_inst_sin_w[47]), .A3(
        round_inst_S_11__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n498) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U118 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n496), .B(
        round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n497) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U117 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n495), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n494), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n499) );
  INV_X1 round_inst_S_11__sbox_inst_com_z_inst_U116 ( .A(round_inst_sin_x[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n494) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U115 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n500), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n518) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U114 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n491), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n493) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U113 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n508), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n490), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n491) );
  INV_X1 round_inst_S_11__sbox_inst_com_z_inst_U112 ( .A(round_inst_sin_w[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n490) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U111 ( .A1(
        round_inst_sin_w[46]), .A2(round_inst_S_11__sbox_inst_com_z_inst_n489), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n513) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U110 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n488), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n508), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n488) );
  INV_X1 round_inst_S_11__sbox_inst_com_z_inst_U108 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n486) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U107 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n484), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U106 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n482), .ZN(
        round_inst_srout2_z[44]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n481), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n482) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U104 ( .A1(
        round_inst_sin_w[44]), .A2(round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n495) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n509), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n479), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n478), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n480) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U101 ( .A1(
        round_inst_sin_w[46]), .A2(round_inst_S_11__sbox_inst_com_z_inst_n485), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n478) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U100 ( .A(round_inst_sin_y[41]), .B(round_inst_sin_x[41]), .Z(round_inst_S_11__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U99 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n492), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n483) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U98 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n476), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n492) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U97 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n474), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n475) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U96 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n472), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n471), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U95 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n470), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n471) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U94 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n496), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n468), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n469) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n467), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n466), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n470) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n465), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n464), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n466) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U91 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n463), .A2(round_inst_sin_w[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n464) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U90 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n462), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U89 ( .A1(
        round_inst_S_11__sbox_inst_n3), .A2(round_inst_sin_y[44]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n462) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U88 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n461), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n460), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U87 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n459), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n458), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n460) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n458) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U85 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n455), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n459) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U84 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n453), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n509), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U83 ( .A1(
        round_inst_sin_w[44]), .A2(round_inst_sin_y[46]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n509) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_sin_w[46]), .A2(round_inst_sin_x[44]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U81 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n452), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n461) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U80 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n450), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U79 ( .A(
        round_inst_S_11__sbox_inst_n5), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n449) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U78 ( .A(round_inst_sin_y[46]), 
        .B(round_inst_sin_w[46]), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n448) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n452), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U76 ( .A(round_inst_sin_w[46]), .B(round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n452) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U75 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n446), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_srout2_z[47]) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n445) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U73 ( .A(round_inst_sin_w[44]), .B(round_inst_S_11__sbox_inst_com_z_inst_n477), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U72 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n477) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U71 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n440), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n441) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U70 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n457), .A2(round_inst_sin_w[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n439) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U69 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n474), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n457) );
  AND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U68 ( .A1(round_inst_sin_w[45]), .A2(round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n474) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n437), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n436), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U66 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n435), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n434), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n436) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U65 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n456), .A2(round_inst_sin_y[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n434) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U64 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n433), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n432), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n456) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U63 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n431), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n430), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U62 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n429), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n428), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n430) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_z_inst_U61 ( .A1(
        round_inst_S_11__sbox_inst_n3), .A2(round_inst_sin_w[47]), .A3(
        round_inst_S_11__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n428) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U60 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n427), .A2(round_inst_sin_w[45]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n429) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U59 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n426), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n425), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n427) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U58 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n424), .A2(
        round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U57 ( .A(round_inst_sin_x[47]), 
        .B(round_inst_sin_y[47]), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n424) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U56 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n422), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U55 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U54 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n419), .A2(round_inst_sin_w[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n420) );
  INV_X1 round_inst_S_11__sbox_inst_com_z_inst_U53 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n419) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U52 ( .A1(
        round_inst_sin_y[47]), .A2(round_inst_S_11__sbox_inst_com_z_inst_n438), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n421) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U51 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n418), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n500), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n423) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U50 ( .A1(
        round_inst_sin_w[47]), .A2(round_inst_S_11__sbox_inst_n5), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n500) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U49 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n417), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n432), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n437) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U48 ( .A1(
        round_inst_sin_w[45]), .A2(round_inst_sin_w[46]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n432) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U47 ( .A(round_inst_sin_x[47]), .B(round_inst_sin_w[47]), .ZN(round_inst_S_11__sbox_inst_com_z_inst_n417) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U46 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n416), .A2(round_inst_sin_x[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n442) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U45 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U44 ( .A(round_inst_sin_w[45]), .B(round_inst_S_11__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n414) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U43 ( .A1(
        round_inst_S_11__sbox_inst_n3), .A2(round_inst_sin_w[46]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n433) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n413), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n415) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U41 ( .A1(
        round_inst_sin_y[45]), .A2(round_inst_sin_w[46]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n413) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U40 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n412), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n438) );
  INV_X1 round_inst_S_11__sbox_inst_com_z_inst_U39 ( .A(round_inst_sin_y[46]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n496) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U38 ( .A(round_inst_sin_y[42]), 
        .B(round_inst_sin_x[42]), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n521), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n517), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n411), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n410), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n517) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U35 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n409), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n408), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n410) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U34 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n407), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n406), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n408) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n405), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n406) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U32 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n403), .A2(round_inst_sin_y[47]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n404) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n402), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n401), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n405) );
  MUX2_X1 round_inst_S_11__sbox_inst_com_z_inst_U30 ( .A(round_inst_sin_x[47]), 
        .B(round_inst_sin_w[47]), .S(
        round_inst_S_11__sbox_inst_com_z_inst_n400), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n401) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_sin_w[45]), .A2(round_inst_S_11__sbox_inst_com_z_inst_n485), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n400) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U28 ( .A(round_inst_sin_w[44]), 
        .B(round_inst_sin_x[44]), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n485) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_z_inst_U27 ( .A1(
        round_inst_sin_w[47]), .A2(round_inst_S_11__sbox_inst_n3), .A3(
        round_inst_S_11__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n402) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U26 ( .A(round_inst_sin_w[44]), 
        .B(round_inst_sin_y[44]), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n473) );
  NAND3_X1 round_inst_S_11__sbox_inst_com_z_inst_U25 ( .A1(
        round_inst_sin_w[44]), .A2(round_inst_sin_x[47]), .A3(
        round_inst_S_11__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n407) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U24 ( .A(
        round_inst_S_11__sbox_inst_n3), .B(round_inst_sin_y[45]), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n454) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U23 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n484), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n409) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_sin_w[44]), .A2(round_inst_sin_y[45]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n447) );
  INV_X1 round_inst_S_11__sbox_inst_com_z_inst_U21 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n425), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n484) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U20 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n399), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n398), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n411) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U19 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n418), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n398) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U18 ( .A(round_inst_sin_y[45]), .B(round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n418) );
  NOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U17 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_11__sbox_inst_com_z_inst_n412), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n399) );
  INV_X1 round_inst_S_11__sbox_inst_com_z_inst_U16 ( .A(round_inst_sin_w[45]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n412) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U15 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n395), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U14 ( .A1(
        round_inst_sin_x[47]), .A2(round_inst_sin_y[44]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n487) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U13 ( .A1(
        round_inst_sin_y[47]), .A2(round_inst_sin_x[44]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n395) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U12 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n394), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n393), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n521) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U11 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n392), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U10 ( .A1(
        round_inst_sin_x[44]), .A2(round_inst_sin_w[45]), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n450) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U9 ( .A1(
        round_inst_S_11__sbox_inst_com_z_inst_n391), .A2(round_inst_sin_w[44]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n392) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U8 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n508), .B(round_inst_sin_y[45]), 
        .ZN(round_inst_S_11__sbox_inst_com_z_inst_n391) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U7 ( .A(round_inst_sin_x[47]), 
        .B(round_inst_S_11__sbox_inst_com_z_inst_n425), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n508) );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U6 ( .A(round_inst_sin_w[47]), 
        .B(round_inst_sin_y[47]), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n425) );
  XNOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U5 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n394) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U4 ( .A1(round_inst_sin_w[47]), .A2(round_inst_sin_x[44]), .ZN(round_inst_S_11__sbox_inst_com_z_inst_n397)
         );
  XOR2_X1 round_inst_S_11__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_11__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_11__sbox_inst_com_z_inst_n451), .Z(
        round_inst_S_11__sbox_inst_com_z_inst_n403) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U2 ( .A1(round_inst_sin_w[44]), .A2(round_inst_S_11__sbox_inst_n3), .ZN(
        round_inst_S_11__sbox_inst_com_z_inst_n451) );
  NAND2_X1 round_inst_S_11__sbox_inst_com_z_inst_U1 ( .A1(round_inst_sin_w[44]), .A2(round_inst_sin_w[45]), .ZN(round_inst_S_11__sbox_inst_com_z_inst_n468)
         );
  INV_X1 round_inst_S_12__sbox_inst_U6 ( .A(round_inst_sin_x[50]), .ZN(
        round_inst_S_12__sbox_inst_n6) );
  INV_X1 round_inst_S_12__sbox_inst_U5 ( .A(round_inst_sin_z[49]), .ZN(
        round_inst_S_12__sbox_inst_n2) );
  INV_X1 round_inst_S_12__sbox_inst_U4 ( .A(round_inst_sin_z[51]), .ZN(
        round_inst_S_12__sbox_inst_n4) );
  INV_X2 round_inst_S_12__sbox_inst_U3 ( .A(round_inst_S_12__sbox_inst_n2), 
        .ZN(round_inst_S_12__sbox_inst_n1) );
  INV_X2 round_inst_S_12__sbox_inst_U2 ( .A(round_inst_S_12__sbox_inst_n4), 
        .ZN(round_inst_S_12__sbox_inst_n3) );
  INV_X2 round_inst_S_12__sbox_inst_U1 ( .A(round_inst_S_12__sbox_inst_n6), 
        .ZN(round_inst_S_12__sbox_inst_n5) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n529), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n528), .ZN(round_inst_sout_w[51]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n526), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n528) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[48]), .A2(round_inst_S_12__sbox_inst_com_w_inst_n525), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n526) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n524), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n523), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n523) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U133 ( .A1(
        round_inst_sin_z[50]), .A2(round_inst_S_12__sbox_inst_com_w_inst_n520), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n521) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U132 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n519), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n518), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n520) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n517), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n516), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n522) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n515), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n514), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n516) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U129 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n518), .A2(
        round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U128 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n513), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n512), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U127 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n511), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n512) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U126 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n508), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n510) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_w_inst_U125 ( .A1(
        round_inst_S_12__sbox_inst_n5), .A2(round_inst_sin_x[48]), .A3(
        round_inst_S_12__sbox_inst_com_w_inst_n507), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n508) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n506), .A2(round_inst_n56), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n509) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U123 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n505), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n511) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U122 ( .A(
        round_inst_sin_x[51]), .B(round_inst_S_12__sbox_inst_com_w_inst_n503), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n505) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_w_inst_U121 ( .A1(
        round_inst_S_12__sbox_inst_n3), .A2(round_inst_n57), .A3(
        round_inst_sin_x[48]), .ZN(round_inst_S_12__sbox_inst_com_w_inst_n513)
         );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U120 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n502), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_sin_y[47]), .B(round_inst_S_12__sbox_inst_com_w_inst_n500), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n501) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U118 ( .A(round_inst_n67), .B(
        round_inst_sin_z[47]), .Z(round_inst_S_12__sbox_inst_com_w_inst_n500)
         );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U117 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n499), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n502) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_sin_x[51]), .B(round_inst_sin_y[51]), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n499) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[49]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U113 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[45]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[45]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U110 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[48]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_12__sbox_inst_n5), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n529), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U105 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n529) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U104 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U102 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_12__sbox_inst_n5), .B(round_inst_sin_z[50]), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U99 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_12__sbox_inst_n1), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n504), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U96 ( .A1(round_inst_n57), 
        .A2(round_inst_sin_x[48]), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n498) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U95 ( .A1(
        round_inst_S_12__sbox_inst_n5), .A2(round_inst_n56), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n504) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U94 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U93 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[50]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U90 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U89 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U88 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n461), .A2(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[50]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U86 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U85 ( .A1(round_inst_sin_z[48]), .A2(round_inst_S_12__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U84 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_sin_y[49]), .A2(round_inst_n56), .A3(
        round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_w_inst_U81 ( .A1(round_inst_n57), 
        .A2(round_inst_n67), .A3(round_inst_n56), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U80 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n525) );
  OR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U79 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_12__sbox_inst_n5), .B(round_inst_n57), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U77 ( .A(round_inst_sin_y[44]), 
        .B(round_inst_sin_z[44]), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n484) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[51])
         );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U73 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U71 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_12__sbox_inst_n3), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U69 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U68 ( .A1(round_inst_n57), 
        .A2(round_inst_n67), .ZN(round_inst_S_12__sbox_inst_com_w_inst_n456)
         );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_12__sbox_inst_n5), .A2(round_inst_sin_y[49]), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U66 ( .A1(
        round_inst_S_12__sbox_inst_n1), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_w_inst_U65 ( .A1(
        round_inst_S_12__sbox_inst_n5), .A2(round_inst_S_12__sbox_inst_n1), 
        .A3(round_inst_sin_x[51]), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n439), .A2(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U62 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U61 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n503), .A2(
        round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U60 ( .A(
        round_inst_S_12__sbox_inst_n3), .B(round_inst_sin_y[51]), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n503) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n506) );
  INV_X1 round_inst_S_12__sbox_inst_com_w_inst_U58 ( .A(round_inst_sin_x[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n486) );
  INV_X1 round_inst_S_12__sbox_inst_com_w_inst_U57 ( .A(round_inst_n57), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U56 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U55 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U54 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U52 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U51 ( .A(round_inst_sin_y[49]), .B(round_inst_S_12__sbox_inst_n1), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U50 ( .A1(
        round_inst_S_12__sbox_inst_n3), .A2(round_inst_S_12__sbox_inst_n1), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U49 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U48 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_w_inst_U47 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n425), .A2(round_inst_sin_x[51]), 
        .A3(round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U46 ( .A(round_inst_sin_y[49]), 
        .B(round_inst_n67), .Z(round_inst_S_12__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_w_inst_U45 ( .A1(
        round_inst_sin_x[51]), .A2(round_inst_sin_y[49]), .A3(
        round_inst_S_12__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U44 ( .A(round_inst_n57), .B(
        round_inst_sin_z[50]), .ZN(round_inst_S_12__sbox_inst_com_w_inst_n465)
         );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U43 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U42 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n517) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U41 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n421), .A2(
        round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U40 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n419), .A2(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U38 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U37 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U36 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n518), .A2(
        round_inst_S_12__sbox_inst_n1), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U35 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n518) );
  INV_X1 round_inst_S_12__sbox_inst_com_w_inst_U34 ( .A(round_inst_sin_x[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n489) );
  INV_X1 round_inst_S_12__sbox_inst_com_w_inst_U33 ( .A(round_inst_sin_y[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n434) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U32 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U31 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U30 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U29 ( .A(round_inst_sin_x[48]), .B(round_inst_sin_z[48]), .ZN(round_inst_S_12__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U28 ( .A1(
        round_inst_sin_y[51]), .A2(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U27 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U26 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n407), .A2(round_inst_sin_y[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U24 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_x[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U23 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U22 ( .A1(round_inst_n67), 
        .A2(round_inst_sin_z[48]), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U21 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_12__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U20 ( .A(round_inst_n67), .B(
        round_inst_S_12__sbox_inst_n1), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U19 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n404), .A2(round_inst_sin_x[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U17 ( .A1(
        round_inst_sin_x[48]), .A2(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U16 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[49]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U15 ( .A(round_inst_n56), .B(
        round_inst_sin_z[48]), .Z(round_inst_S_12__sbox_inst_com_w_inst_n418)
         );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U13 ( .A(round_inst_sin_x[48]), .B(round_inst_S_12__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U11 ( .A1(
        round_inst_S_12__sbox_inst_com_w_inst_n398), .A2(round_inst_sin_x[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U9 ( .A(round_inst_sin_y[51]), 
        .B(round_inst_n67), .ZN(round_inst_S_12__sbox_inst_com_w_inst_n396) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U8 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_12__sbox_inst_n1), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U7 ( .A(
        round_inst_S_12__sbox_inst_n3), .B(round_inst_sin_x[51]), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n507) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U6 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n519), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_12__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U5 ( .A(
        round_inst_S_12__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_12__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U4 ( .A1(round_inst_n67), 
        .A2(round_inst_n56), .ZN(round_inst_S_12__sbox_inst_com_w_inst_n475)
         );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U3 ( .A1(round_inst_sin_x[48]), .A2(round_inst_sin_y[49]), .ZN(round_inst_S_12__sbox_inst_com_w_inst_n477)
         );
  NAND2_X1 round_inst_S_12__sbox_inst_com_w_inst_U2 ( .A1(round_inst_sin_x[51]), .A2(round_inst_n56), .ZN(round_inst_S_12__sbox_inst_com_w_inst_n519) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_w_inst_U1 ( .A(round_inst_sin_y[46]), 
        .B(round_inst_sin_z[46]), .Z(
        round_inst_S_12__sbox_inst_com_w_inst_n402) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U136 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n512), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n511), .ZN(round_inst_sout_x[48]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n510), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n509), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n511) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U134 ( .A(round_inst_n57), 
        .B(round_inst_S_12__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U133 ( .A(round_inst_sin_z[44]), .B(round_inst_S_12__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n510) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U132 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n512), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n506), .Z(round_inst_srout2_x[2]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U130 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n503), .A2(round_inst_sin_z[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U129 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U127 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U126 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U125 ( .A1(round_inst_n57), 
        .A2(round_inst_sin_w[48]), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U124 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U122 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U121 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U118 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n508), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n487) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U115 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n481) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_x_inst_U114 ( .A1(
        round_inst_sin_z[50]), .A2(round_inst_sin_w[48]), .A3(
        round_inst_S_12__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n489) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n478), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n475), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n477) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n474), .B(round_inst_sin_z[47]), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n475) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_w[50]), .A2(round_inst_S_12__sbox_inst_com_x_inst_n508), 
        .A3(round_inst_sin_z[48]), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n473), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n478) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n470), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n473) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n468), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n512) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n467), .A2(round_inst_n57), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n468) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n467) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n469) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n465), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n463), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_srout2_x[0]) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U100 ( .A1(round_inst_n56), 
        .A2(round_inst_sin_z[50]), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[45]), .B(round_inst_S_12__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n461), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n462) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n466), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n460) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n458), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n457), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_12__sbox_inst_n1), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n459), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n456), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n455), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n454), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n453), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n455) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n452), .A2(round_inst_sin_w[50]), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n451), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n450), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n454) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n449), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n448), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n447), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n446), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n448) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n445), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n446) );
  MUX2_X1 round_inst_S_12__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n444), .B(round_inst_n57), .S(
        round_inst_n56), .Z(round_inst_S_12__sbox_inst_com_x_inst_n445) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n443), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_12__sbox_inst_com_x_inst_U85 ( .A(round_inst_n57), .B(
        round_inst_sin_z[50]), .S(round_inst_sin_z[48]), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n443) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n442), .A2(round_inst_sin_w[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n449) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n441), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n440), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n451) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_w[48]), 
        .A3(round_inst_sin_z[50]), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n440) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n439), .A2(round_inst_sin_w[49]), 
        .A3(round_inst_n57), .ZN(round_inst_S_12__sbox_inst_com_x_inst_n441)
         );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U80 ( .A(round_inst_n56), .B(
        round_inst_sin_z[48]), .Z(round_inst_S_12__sbox_inst_com_x_inst_n439)
         );
  NAND3_X1 round_inst_S_12__sbox_inst_com_x_inst_U79 ( .A1(round_inst_n56), 
        .A2(round_inst_S_12__sbox_inst_com_x_inst_n444), .A3(
        round_inst_S_12__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n456) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n459) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U77 ( .A1(round_inst_n56), 
        .A2(round_inst_n57), .ZN(round_inst_S_12__sbox_inst_com_x_inst_n482)
         );
  AND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U76 ( .A1(round_inst_n57), 
        .A2(round_inst_sin_z[48]), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n490) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n461) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U74 ( .A1(round_inst_n56), 
        .A2(round_inst_sin_w[50]), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n497) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n436), .ZN(
        round_inst_srout2_x[3]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n435), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n434), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n436) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U71 ( .A(round_inst_n56), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n434) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n433), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n432), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U69 ( .A1(
        round_inst_sin_z[48]), .A2(round_inst_S_12__sbox_inst_com_x_inst_n508), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n432) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n431), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n430), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n433) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n429), .A2(round_inst_n56), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n428), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n427) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_12__sbox_inst_n1), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n431) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n452) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[46]), 
        .B(round_inst_S_12__sbox_inst_com_x_inst_n437), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n435) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n424), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n423), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n422), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n421), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n423) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n420), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n419), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n421) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n418), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n419) );
  NOR3_X1 round_inst_S_12__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n470), .A3(
        round_inst_S_12__sbox_inst_com_x_inst_n416), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n417) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n415), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n414), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n418) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n413), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n414) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U53 ( .A1(round_inst_n57), 
        .A2(round_inst_S_12__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n412) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U52 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n442), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_12__sbox_inst_n1), .A2(round_inst_n57), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n442) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_x_inst_U50 ( .A1(round_inst_n57), 
        .A2(round_inst_S_12__sbox_inst_com_x_inst_n476), .A3(
        round_inst_S_12__sbox_inst_com_x_inst_n411), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n420) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U49 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n410), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n422) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U48 ( .A1(round_inst_n57), 
        .A2(round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n464) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U47 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n410) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n409), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n407), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n406), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n405), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n404), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n406) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U43 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n465), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n404) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U42 ( .A(round_inst_sin_w[49]), 
        .B(round_inst_S_12__sbox_inst_n1), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n438) );
  AND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U41 ( .A1(round_inst_sin_z[50]), .A2(round_inst_S_12__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n465) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U40 ( .A1(
        round_inst_S_12__sbox_inst_n3), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n405) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n476), .A3(
        round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n407) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U38 ( .A(round_inst_sin_z[50]), 
        .B(round_inst_sin_w[50]), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U37 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n403), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n402), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U36 ( .A(round_inst_sin_w[50]), 
        .B(round_inst_n57), .Z(round_inst_S_12__sbox_inst_com_x_inst_n402) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U35 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n401), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n400), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n399), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n400) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U33 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n398) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U32 ( .A1(
        round_inst_sin_z[48]), .A2(round_inst_S_12__sbox_inst_com_x_inst_n476), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n425) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U31 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n479), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n471) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_12__sbox_inst_n3), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n426), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n399) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U28 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n401) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_12__sbox_inst_n1), .A3(round_inst_n56), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n396) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n411), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U23 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n392), .A2(round_inst_sin_w[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U21 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_x_inst_U19 ( .A1(
        round_inst_sin_z[48]), .A2(round_inst_S_12__sbox_inst_com_x_inst_n508), 
        .A3(round_inst_sin_w[49]), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n388) );
  MUX2_X1 round_inst_S_12__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n411), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n508), .S(
        round_inst_S_12__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U17 ( .A1(round_inst_n56), 
        .A2(round_inst_S_12__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n491), .B(
        round_inst_S_12__sbox_inst_n3), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n411) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U15 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U14 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n384), .A2(round_inst_sin_z[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n403), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U10 ( .A(round_inst_sin_w[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U9 ( .A1(
        round_inst_S_12__sbox_inst_n1), .A2(
        round_inst_S_12__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n403) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U8 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n508) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U7 ( .A(round_inst_sin_y[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n413) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_12__sbox_inst_com_x_inst_n426), .Z(
        round_inst_S_12__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U4 ( .A1(round_inst_n56), 
        .A2(round_inst_sin_w[49]), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n426) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_12__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_w[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_12__sbox_inst_com_x_inst_n416), .ZN(
        round_inst_S_12__sbox_inst_com_x_inst_n476) );
  INV_X1 round_inst_S_12__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_y[49]), 
        .ZN(round_inst_S_12__sbox_inst_com_x_inst_n416) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U138 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n519), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n518), .Z(round_inst_sout_y[48])
         );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n516), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n518) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n515), .B(
        round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n516) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U135 ( .A(round_inst_sin_x[44]), .B(round_inst_S_12__sbox_inst_com_y_inst_n514), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U134 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n513), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n512), .ZN(
        round_inst_srout2_y[2]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n519), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n510), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n519) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n507), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n509) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U130 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n506), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n507) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n508) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U128 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n503), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n502), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n513) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n501), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n500), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n502) );
  NOR3_X1 round_inst_S_12__sbox_inst_com_y_inst_U126 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n499), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n498), .A3(
        round_inst_S_12__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n500) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U125 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n496), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n495), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n501) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U124 ( .A1(
        round_inst_sin_x[51]), .A2(round_inst_S_12__sbox_inst_com_y_inst_n494), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n495) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U123 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n493), .A2(
        round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U122 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n492), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n491), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U121 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n490), .A2(round_inst_sin_w[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n492) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U120 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n489), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n488), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n503) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U119 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n487), .A2(
        round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n488) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U118 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n486), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n485), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n487) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U117 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n504), .A2(round_inst_sin_w[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n485) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n515), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n486) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U115 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n482), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n489) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n481), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n480), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n482) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U113 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n479), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U112 ( .A(
        round_inst_S_12__sbox_inst_n1), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n478), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n481) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n477), .B(round_inst_sin_x[47]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n478) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_y_inst_U110 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n515), .A2(
        round_inst_S_12__sbox_inst_n3), .A3(
        round_inst_S_12__sbox_inst_com_y_inst_n476), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n477) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U109 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n483) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_y_inst_U108 ( .A1(
        round_inst_sin_w[48]), .A2(round_inst_sin_w[51]), .A3(
        round_inst_S_12__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_12__sbox_inst_com_y_inst_U107 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n506), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_12__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U106 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[0]) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U105 ( .A1(
        round_inst_S_12__sbox_inst_n5), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U104 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n510), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U99 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_12__sbox_inst_n1), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U98 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U96 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n476), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n491) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_y_inst_U95 ( .A1(
        round_inst_sin_w[48]), .A2(round_inst_n67), .A3(
        round_inst_S_12__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U94 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U93 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U92 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U89 ( .A1(
        round_inst_S_12__sbox_inst_n1), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_12__sbox_inst_com_y_inst_U88 ( .A(
        round_inst_S_12__sbox_inst_n5), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n504), .S(
        round_inst_S_12__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U87 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U85 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U81 ( .A(
        round_inst_S_12__sbox_inst_n1), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n479), .B(round_inst_sin_x[45]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U79 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n479) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n515), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U77 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n438), .Z(round_inst_srout2_y[3]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n484), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U72 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U71 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U70 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n484), .A2(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_12__sbox_inst_n1), .A2(round_inst_sin_w[48]), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[51]), 
        .A3(round_inst_S_12__sbox_inst_n1), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U67 ( .A(round_inst_sin_w[48]), 
        .B(round_inst_S_12__sbox_inst_com_y_inst_n476), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U66 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U64 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U62 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U60 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U59 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U58 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n484), .A2(round_inst_sin_w[49]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n422) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n418), .A2(
        round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U55 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U54 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U53 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n414), .B(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U51 ( .A(round_inst_sin_w[49]), .B(round_inst_S_12__sbox_inst_n1), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U50 ( .A1(
        round_inst_S_12__sbox_inst_n1), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n476), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n444) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U49 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n473), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n476) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U48 ( .A(round_inst_sin_x[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_12__sbox_inst_n1), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U46 ( .A(round_inst_sin_x[46]), 
        .B(round_inst_S_12__sbox_inst_com_y_inst_n514), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n514) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[49]), 
        .B(round_inst_sin_x[51]), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U41 ( .A(round_inst_n67), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n499) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n484), .B(round_inst_sin_w[48]), 
        .Z(round_inst_S_12__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n484) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U36 ( .A(round_inst_sin_z[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n497) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_12__sbox_inst_n1), .B(round_inst_S_12__sbox_inst_n3), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n490), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n498) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_12__sbox_inst_n5), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n506), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n490) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U27 ( .A1(
        round_inst_sin_w[49]), .A2(round_inst_S_12__sbox_inst_n3), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n515), .A2(round_inst_sin_w[49]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_12__sbox_inst_n1), .A2(round_inst_sin_w[51]), .A3(
        round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_12__sbox_inst_n1), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n505), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n506), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_12__sbox_inst_n3), .B(round_inst_sin_w[51]), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U17 ( .A(
        round_inst_S_12__sbox_inst_n3), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[51]), .B(round_inst_sin_x[51]), .ZN(round_inst_S_12__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_y_inst_U13 ( .A1(round_inst_n67), 
        .A2(round_inst_sin_w[51]), .A3(
        round_inst_S_12__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_y_inst_U12 ( .A1(
        round_inst_S_12__sbox_inst_n3), .A2(
        round_inst_S_12__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_12__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[49]), 
        .B(round_inst_n67), .S(round_inst_S_12__sbox_inst_com_y_inst_n504), 
        .Z(round_inst_S_12__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_y_inst_U9 ( .A1(round_inst_n67), 
        .A2(round_inst_S_12__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_12__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_12__sbox_inst_n3), .B(round_inst_sin_x[51]), .Z(
        round_inst_S_12__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_12__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_12__sbox_inst_n1), .A3(round_inst_sin_x[51]), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n515), .B(
        round_inst_S_12__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n504) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[50]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_12__sbox_inst_com_y_inst_n506), .ZN(
        round_inst_S_12__sbox_inst_com_y_inst_n515) );
  INV_X1 round_inst_S_12__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[50]), 
        .ZN(round_inst_S_12__sbox_inst_com_y_inst_n506) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U132 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n517), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n516), .ZN(round_inst_sout_z[48]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n515), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n514), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_sin_w[50]), .B(round_inst_sin_w[51]), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n514) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_x[44]), .B(round_inst_sin_y[44]), .Z(round_inst_S_12__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U128 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n512), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n517) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_srout2_z[2]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n510), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n509), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n511) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n508), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n507), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n509) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U124 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n506), .A2(round_inst_n56), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U123 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n505), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n504), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n508) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n503), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n502), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_sin_w[49]), .B(round_inst_sin_x[47]), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U120 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n501), .B(round_inst_sin_y[47]), 
        .Z(round_inst_S_12__sbox_inst_com_z_inst_n503) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U119 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n500), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n499), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n501) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U118 ( .A1(round_inst_n57), 
        .A2(round_inst_S_12__sbox_inst_com_z_inst_n498), .A3(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n499) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U117 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_x[48]), 
        .A3(round_inst_sin_w[51]), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n500) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U116 ( .A(
        round_inst_S_12__sbox_inst_n5), .B(round_inst_n57), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n496) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U115 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_12__sbox_inst_n5), .A3(
        round_inst_S_12__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n505) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U114 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n491), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n493) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n490), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n489), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n491) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U111 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n488), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n486), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n490) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_sin_w[50]), .A2(round_inst_S_12__sbox_inst_com_z_inst_n495), 
        .A3(round_inst_n56), .ZN(round_inst_S_12__sbox_inst_com_z_inst_n492)
         );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U108 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n484), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n513) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U107 ( .A1(
        round_inst_sin_w[50]), .A2(round_inst_S_12__sbox_inst_com_z_inst_n498), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U106 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n506), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n484) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n482), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n481), .Z(round_inst_srout2_z[0]) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n479), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n478), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n483), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n483) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U101 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n475), .A2(round_inst_sin_x[48]), 
        .A3(round_inst_sin_w[50]), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U100 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n474), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n477) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U99 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n472), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .A3(round_inst_n57), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n473) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U98 ( .A(round_inst_sin_w[49]), 
        .B(round_inst_sin_y[49]), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U97 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n471), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n474) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U96 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n469), .A2(
        round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n470) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U95 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n467), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n471) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n466), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n465), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n464), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n463), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n462), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n461), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U91 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n460), .A2(round_inst_n57), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n461) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U90 ( .A1(round_inst_n67), 
        .A2(round_inst_S_12__sbox_inst_n5), .A3(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n462) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U89 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n459), .A2(round_inst_n56), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_w[50]), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n466) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U87 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U85 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n453), .A2(round_inst_n57), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n454) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U84 ( .A(round_inst_sin_w[49]), .B(round_inst_S_12__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U83 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n451), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_sin_w[50]), .A2(round_inst_sin_x[48]), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n478) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U81 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n487), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n448) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U79 ( .A(round_inst_sin_y[45]), 
        .B(round_inst_sin_x[45]), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n447) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U78 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n487) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n446), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U76 ( .A(round_inst_sin_w[50]), .B(round_inst_n57), .ZN(round_inst_S_12__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U75 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_srout2_z[3]) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n512), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U72 ( .A1(
        round_inst_sin_x[48]), .A2(round_inst_sin_w[51]), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n441) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U71 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n458), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n440), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n442) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U70 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n498), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U69 ( .A(round_inst_sin_w[51]), .B(round_inst_S_12__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n498) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U68 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n494) );
  MUX2_X1 round_inst_S_12__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n495), .B(round_inst_sin_w[51]), 
        .S(round_inst_S_12__sbox_inst_com_z_inst_n436), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n437) );
  OR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U66 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n436) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U65 ( .A(round_inst_sin_x[48]), .B(round_inst_S_12__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n486) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U64 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n438) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U63 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n495), .A3(
        round_inst_S_12__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U62 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n430), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n429) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U59 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n426), .A2(round_inst_sin_w[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U58 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n422), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n424) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U56 ( .A1(
        round_inst_sin_x[48]), .A2(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U55 ( .A1(
        round_inst_sin_y[49]), .A2(round_inst_sin_x[48]), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n425) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U54 ( .A1(round_inst_n56), 
        .A2(round_inst_S_12__sbox_inst_com_z_inst_n495), .A3(
        round_inst_sin_w[49]), .ZN(round_inst_S_12__sbox_inst_com_z_inst_n428)
         );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U53 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_y[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U52 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n460), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n423), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n469) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U50 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .A2(round_inst_sin_y[49]), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n423) );
  AND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U49 ( .A1(round_inst_sin_w[49]), .A2(round_inst_sin_x[48]), .ZN(round_inst_S_12__sbox_inst_com_z_inst_n460)
         );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U48 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n421) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U47 ( .A1(
        round_inst_sin_w[49]), .A2(round_inst_S_12__sbox_inst_com_z_inst_n497), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U46 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .A2(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n419), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n418), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n432) );
  INV_X1 round_inst_S_12__sbox_inst_com_z_inst_U44 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U43 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .B(round_inst_n56), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n451) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n417), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U41 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n497), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n449) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U39 ( .A1(
        round_inst_sin_w[51]), .A2(round_inst_S_12__sbox_inst_com_z_inst_n413), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n414) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U38 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n415) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U35 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n506), .A2(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n409) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U34 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n407) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U32 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n405) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n404) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U30 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n506), .A2(round_inst_sin_y[49]), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n402) );
  AND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_S_12__sbox_inst_n5), .A2(round_inst_sin_w[51]), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n506) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n401), .A2(round_inst_n57), .A3(
        round_inst_sin_w[49]), .ZN(round_inst_S_12__sbox_inst_com_z_inst_n403)
         );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U27 ( .A(round_inst_sin_w[51]), 
        .B(round_inst_S_12__sbox_inst_com_z_inst_n495), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n401) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U26 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n399), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n406) );
  MUX2_X1 round_inst_S_12__sbox_inst_com_z_inst_U25 ( .A(round_inst_sin_y[51]), 
        .B(round_inst_S_12__sbox_inst_com_z_inst_n398), .S(
        round_inst_S_12__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U24 ( .A1(
        round_inst_sin_w[49]), .A2(round_inst_S_12__sbox_inst_n5), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U23 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n398) );
  NOR3_X1 round_inst_S_12__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n488), .A3(
        round_inst_S_12__sbox_inst_com_z_inst_n395), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U21 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n394), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n395) );
  INV_X1 round_inst_S_12__sbox_inst_com_z_inst_U20 ( .A(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n394) );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U19 ( .A(round_inst_sin_w[51]), .B(round_inst_sin_y[51]), .ZN(round_inst_S_12__sbox_inst_com_z_inst_n488) );
  AND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U18 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n459), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U17 ( .A1(
        round_inst_sin_w[50]), .A2(round_inst_n67), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n459) );
  INV_X1 round_inst_S_12__sbox_inst_com_z_inst_U16 ( .A(round_inst_sin_w[49]), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U15 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n393), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U14 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n391), .A2(round_inst_n57), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U13 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_12__sbox_inst_com_z_inst_n390), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U12 ( .A1(
        round_inst_sin_w[49]), .A2(round_inst_sin_y[51]), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n390) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U11 ( .A1(round_inst_n67), 
        .A2(round_inst_sin_w[51]), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n418) );
  NOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U10 ( .A1(
        round_inst_S_12__sbox_inst_com_z_inst_n439), .A2(
        round_inst_S_12__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_12__sbox_inst_com_z_inst_U9 ( .A1(round_inst_sin_w[50]), .A2(round_inst_sin_w[49]), .ZN(round_inst_S_12__sbox_inst_com_z_inst_n456)
         );
  XNOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U8 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n495), .B(round_inst_sin_y[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n439) );
  NAND3_X1 round_inst_S_12__sbox_inst_com_z_inst_U7 ( .A1(round_inst_sin_w[50]), .A2(round_inst_S_12__sbox_inst_com_z_inst_n495), .A3(
        round_inst_S_12__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U6 ( .A(round_inst_n67), .B(
        round_inst_sin_y[49]), .Z(round_inst_S_12__sbox_inst_com_z_inst_n475)
         );
  INV_X1 round_inst_S_12__sbox_inst_com_z_inst_U5 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n495) );
  INV_X1 round_inst_S_12__sbox_inst_com_z_inst_U4 ( .A(round_inst_sin_x[51]), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n397) );
  INV_X1 round_inst_S_12__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_12__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_12__sbox_inst_com_z_inst_n497) );
  INV_X1 round_inst_S_12__sbox_inst_com_z_inst_U2 ( .A(round_inst_sin_w[48]), 
        .ZN(round_inst_S_12__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_12__sbox_inst_com_z_inst_U1 ( .A(round_inst_sin_y[46]), 
        .B(round_inst_sin_x[46]), .Z(
        round_inst_S_12__sbox_inst_com_z_inst_n417) );
  INV_X1 round_inst_S_13__sbox_inst_U4 ( .A(round_inst_sin_x[53]), .ZN(
        round_inst_S_13__sbox_inst_n4) );
  INV_X1 round_inst_S_13__sbox_inst_U3 ( .A(round_inst_sin_z[53]), .ZN(
        round_inst_S_13__sbox_inst_n2) );
  INV_X2 round_inst_S_13__sbox_inst_U2 ( .A(round_inst_S_13__sbox_inst_n2), 
        .ZN(round_inst_S_13__sbox_inst_n1) );
  INV_X2 round_inst_S_13__sbox_inst_U1 ( .A(round_inst_S_13__sbox_inst_n4), 
        .ZN(round_inst_S_13__sbox_inst_n3) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n531), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n530), .ZN(round_inst_sout_w[55]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U139 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n529), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n528), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n530) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U138 ( .A1(
        round_inst_sin_z[52]), .A2(round_inst_S_13__sbox_inst_com_w_inst_n527), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n528) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n526), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n525), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n529) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U136 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n524), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n523), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n525) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U135 ( .A1(
        round_inst_sin_z[54]), .A2(round_inst_S_13__sbox_inst_com_w_inst_n522), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n521), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n522) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n519), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n518), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U132 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n517), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n516), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n518) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U131 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n520), .A2(round_inst_n68), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n515), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n514), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n513), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n512), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U128 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n511), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n512) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_w_inst_U127 ( .A1(round_inst_n68), 
        .A2(round_inst_sin_x[52]), .A3(
        round_inst_S_13__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n510) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n508), .A2(round_inst_sin_y[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n511) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U125 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n507), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n513) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U124 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n507) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_w_inst_U123 ( .A1(
        round_inst_sin_z[55]), .A2(round_inst_n58), .A3(round_inst_sin_x[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U122 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n526) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U121 ( .A(
        round_inst_sin_y[51]), .B(round_inst_S_13__sbox_inst_com_w_inst_n501), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U120 ( .A(
        round_inst_S_13__sbox_inst_n3), .B(round_inst_sin_z[51]), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n501) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U119 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n505), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[53]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[49]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U113 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[49]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U112 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[52]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U110 ( .A(round_inst_n68), 
        .B(round_inst_S_13__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n531), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n531) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U105 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U103 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U102 ( .A(round_inst_n68), 
        .B(round_inst_sin_z[54]), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U101 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U100 ( .A1(
        round_inst_S_13__sbox_inst_n1), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U99 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U98 ( .A1(round_inst_n58), 
        .A2(round_inst_sin_x[52]), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U97 ( .A1(round_inst_n68), 
        .A2(round_inst_sin_y[52]), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n506) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U94 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U92 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U91 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U90 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n461), .A2(
        round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U89 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U88 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n459), .A2(round_inst_n68), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U87 ( .A1(round_inst_sin_z[52]), .A2(round_inst_S_13__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U85 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_w_inst_U84 ( .A1(
        round_inst_sin_y[53]), .A2(round_inst_sin_y[52]), .A3(round_inst_n68), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_w_inst_U83 ( .A1(round_inst_n58), 
        .A2(round_inst_S_13__sbox_inst_n3), .A3(round_inst_sin_y[52]), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U82 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n527) );
  OR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U81 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U80 ( .A(round_inst_n68), .B(
        round_inst_n58), .ZN(round_inst_S_13__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U79 ( .A(round_inst_n56), .B(
        round_inst_sin_z[48]), .Z(round_inst_S_13__sbox_inst_com_w_inst_n484)
         );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[55])
         );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U73 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U72 ( .A1(
        round_inst_sin_z[55]), .A2(round_inst_S_13__sbox_inst_com_w_inst_n440), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U71 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U70 ( .A1(round_inst_n58), 
        .A2(round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U69 ( .A1(round_inst_n68), 
        .A2(round_inst_sin_y[53]), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_13__sbox_inst_n1), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n508), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_w_inst_U67 ( .A1(round_inst_n68), 
        .A2(round_inst_S_13__sbox_inst_n1), .A3(
        round_inst_S_13__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U66 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n439), .A2(
        round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U64 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n508), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U63 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n504), .A2(round_inst_n68), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U62 ( .A(round_inst_sin_z[55]), 
        .B(round_inst_S_13__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n504) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U61 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n508) );
  INV_X1 round_inst_S_13__sbox_inst_com_w_inst_U60 ( .A(round_inst_n58), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U59 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U58 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U57 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n433), .A2(round_inst_n68), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U56 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U55 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U54 ( .A(round_inst_sin_y[53]), .B(round_inst_S_13__sbox_inst_n1), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U53 ( .A1(
        round_inst_sin_z[55]), .A2(round_inst_S_13__sbox_inst_n1), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U52 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U51 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_w_inst_U50 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n505), .A3(round_inst_n68), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U49 ( .A(round_inst_sin_y[53]), 
        .B(round_inst_S_13__sbox_inst_n3), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_w_inst_U48 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n505), .A2(round_inst_sin_y[53]), 
        .A3(round_inst_S_13__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U47 ( .A(round_inst_n58), .B(
        round_inst_sin_z[54]), .ZN(round_inst_S_13__sbox_inst_com_w_inst_n465)
         );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U45 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U44 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n421), .A2(round_inst_sin_z[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U43 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U42 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n419), .A2(
        round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U40 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n520), .A2(
        round_inst_S_13__sbox_inst_n1), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U38 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n520) );
  INV_X1 round_inst_S_13__sbox_inst_com_w_inst_U37 ( .A(round_inst_sin_x[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n489) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U36 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U33 ( .A(round_inst_sin_x[52]), .B(round_inst_sin_z[52]), .ZN(round_inst_S_13__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U32 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n498), .A2(
        round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U31 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U30 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U29 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U28 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U27 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U26 ( .A1(
        round_inst_S_13__sbox_inst_n3), .A2(round_inst_sin_z[52]), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U24 ( .A(
        round_inst_S_13__sbox_inst_n3), .B(round_inst_S_13__sbox_inst_n1), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_13__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U22 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U21 ( .A1(
        round_inst_sin_x[52]), .A2(round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U20 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[53]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U19 ( .A(round_inst_sin_y[52]), 
        .B(round_inst_sin_z[52]), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n418) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U17 ( .A(round_inst_sin_x[52]), .B(round_inst_S_13__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U15 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n398), .A2(round_inst_sin_x[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U13 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n498), .B(
        round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_13__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_13__sbox_inst_com_w_inst_U11 ( .A(round_inst_sin_y[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_13__sbox_inst_n1), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U9 ( .A(round_inst_sin_z[55]), 
        .B(round_inst_S_13__sbox_inst_com_w_inst_n505), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U8 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n521), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U7 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_13__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_13__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U6 ( .A1(
        round_inst_S_13__sbox_inst_n3), .A2(round_inst_sin_y[52]), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U5 ( .A1(round_inst_sin_x[52]), .A2(round_inst_sin_y[53]), .ZN(round_inst_S_13__sbox_inst_com_w_inst_n477)
         );
  NAND2_X1 round_inst_S_13__sbox_inst_com_w_inst_U4 ( .A1(
        round_inst_S_13__sbox_inst_com_w_inst_n505), .A2(round_inst_sin_y[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n521) );
  INV_X1 round_inst_S_13__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_13__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_13__sbox_inst_com_w_inst_n505) );
  INV_X1 round_inst_S_13__sbox_inst_com_w_inst_U2 ( .A(round_inst_sin_x[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_w_inst_n486) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_w_inst_U1 ( .A(round_inst_n57), .B(
        round_inst_sin_z[50]), .Z(round_inst_S_13__sbox_inst_com_w_inst_n402)
         );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U143 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n518), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n517), .Z(round_inst_sout_x[52])
         );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U142 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n516), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n515), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n517) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U141 ( .A(round_inst_n58), 
        .B(round_inst_sin_y[55]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n515) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U140 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n514), .B(round_inst_sin_z[48]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n516) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U139 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n513), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n512), .ZN(
        round_inst_srout2_x[22]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U138 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n510), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n512) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U137 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n509), .A2(round_inst_sin_z[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n510) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U136 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n509) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U135 ( .A1(round_inst_n58), 
        .A2(round_inst_S_13__sbox_inst_com_x_inst_n506), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n507) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n504), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n511) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U133 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n503), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n502), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n504) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U132 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n508), .A2(round_inst_sin_w[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n502) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n501), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n500), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U130 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n499), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n498), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n500) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_x_inst_U129 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n497), .A2(round_inst_sin_w[54]), 
        .A3(round_inst_sin_y[55]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n498) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n496), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n495), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n499) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_x_inst_U127 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n494), .A2(round_inst_sin_y[52]), 
        .A3(round_inst_n58), .ZN(round_inst_S_13__sbox_inst_com_x_inst_n495)
         );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U126 ( .A(round_inst_sin_y[55]), .B(round_inst_sin_z[55]), .Z(round_inst_S_13__sbox_inst_com_x_inst_n494) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U125 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n493), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n496) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_x_inst_U124 ( .A1(round_inst_n58), 
        .A2(round_inst_sin_z[52]), .A3(round_inst_sin_z[55]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n501) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n492), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n505) );
  OR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U122 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n493), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n491) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U121 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n488) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n484), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n486) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U118 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n483), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n484) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n506), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n482) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U116 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n480), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n479), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n483) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U115 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n478), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n479) );
  AND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U114 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n481), .A2(round_inst_sin_z[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n477) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .B(round_inst_sin_z[51]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n478) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_x_inst_U112 ( .A1(round_inst_n58), 
        .A2(round_inst_sin_w[52]), .A3(round_inst_sin_z[55]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n480) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_x_inst_U111 ( .A1(round_inst_n58), 
        .A2(round_inst_sin_y[52]), .A3(
        round_inst_S_13__sbox_inst_com_x_inst_n506), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n475), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n493), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n487) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_x_inst_U109 ( .A1(round_inst_n58), 
        .A2(round_inst_sin_z[52]), .A3(round_inst_sin_y[55]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n489) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U108 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n518), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n474), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n513) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U107 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n473), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n518) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U106 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n471), .A2(round_inst_n58), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n472) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U105 ( .A(
        round_inst_sin_z[55]), .B(round_inst_S_13__sbox_inst_com_x_inst_n470), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n471) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n508), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n473) );
  AND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U103 ( .A1(
        round_inst_sin_z[54]), .A2(round_inst_sin_y[55]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n508) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n468), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n467), .ZN(
        round_inst_srout2_x[20]) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n493), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n467) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U100 ( .A1(
        round_inst_sin_y[52]), .A2(round_inst_sin_z[54]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n493) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U99 ( .A1(round_inst_n58), 
        .A2(round_inst_S_13__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n466) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n465), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n468) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n463), .B(round_inst_sin_z[49]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n464) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n463) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n462), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n481) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n460), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n459), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n469) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U93 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n458), .A2(round_inst_n58), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n459) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U92 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n457), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n458) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U91 ( .A1(
        round_inst_S_13__sbox_inst_n1), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n455), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n454), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n460) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U89 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n453), .A2(round_inst_sin_w[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n454) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U88 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n451), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n453) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U87 ( .A1(round_inst_n58), 
        .A2(round_inst_S_13__sbox_inst_n1), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n452) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U86 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n450), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n449), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n455) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U85 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n448), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n447), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n449) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U84 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n446), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n445), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n447) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U83 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n443), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n445) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U82 ( .A(round_inst_sin_w[54]), .B(round_inst_sin_z[54]), .ZN(round_inst_S_13__sbox_inst_com_x_inst_n443) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U81 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n442), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U80 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n441), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n440), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n448) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U79 ( .A1(round_inst_n58), 
        .A2(round_inst_sin_z[52]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n441) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_x_inst_U78 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n497), .A3(
        round_inst_S_13__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U77 ( .A(round_inst_sin_z[54]), 
        .B(round_inst_sin_w[54]), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n439) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U76 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n514), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_srout2_x[23]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n437), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n436), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U74 ( .A(round_inst_sin_y[52]), .B(round_inst_S_13__sbox_inst_com_x_inst_n474), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n436) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n435), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n434), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n433), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n432), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n434) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U71 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n431), .A2(round_inst_sin_w[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n432) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n430), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n429), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n431) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U69 ( .A1(
        round_inst_S_13__sbox_inst_n1), .A2(round_inst_sin_y[55]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n429) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U68 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_z[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U67 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n428), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n433) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n426), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n427) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n424), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n423), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n422), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n421), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n423) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U63 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n506), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n421) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U62 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n440), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n456) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U61 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .B(round_inst_sin_w[53]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n440) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U60 ( .A1(
        round_inst_sin_z[55]), .A2(round_inst_S_13__sbox_inst_com_x_inst_n442), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n422) );
  AND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U59 ( .A1(round_inst_sin_y[52]), .A2(round_inst_S_13__sbox_inst_com_x_inst_n420), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n442) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_x_inst_U58 ( .A1(
        round_inst_sin_w[53]), .A2(round_inst_S_13__sbox_inst_com_x_inst_n497), 
        .A3(round_inst_sin_y[55]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U57 ( .A(round_inst_sin_z[52]), 
        .B(round_inst_sin_y[52]), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n497) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n419), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n426) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U55 ( .A1(
        round_inst_S_13__sbox_inst_n1), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U54 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n416), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n417) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U53 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n470), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n416) );
  MUX2_X1 round_inst_S_13__sbox_inst_com_x_inst_U52 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n419), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n414), .S(
        round_inst_S_13__sbox_inst_com_x_inst_n413), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n435) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_sin_y[55]), .A2(round_inst_S_13__sbox_inst_com_x_inst_n412), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n413) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U50 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_y[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n412) );
  MUX2_X1 round_inst_S_13__sbox_inst_com_x_inst_U49 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n411), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n410), .S(
        round_inst_S_13__sbox_inst_com_x_inst_n409), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n414) );
  NOR3_X1 round_inst_S_13__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n410), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n462), .A3(
        round_inst_S_13__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n411) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U47 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n475), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n419), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n410) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U46 ( .A(round_inst_sin_z[50]), 
        .B(round_inst_S_13__sbox_inst_com_x_inst_n465), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n407), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n406), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n465) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U44 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n405), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n406) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U43 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n405) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U42 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n418), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n404) );
  INV_X1 round_inst_S_13__sbox_inst_com_x_inst_U41 ( .A(round_inst_sin_w[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n461) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U40 ( .A(round_inst_sin_z[55]), .B(round_inst_S_13__sbox_inst_com_x_inst_n506), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n418) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U39 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n403), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n402), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n407) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_x_inst_U38 ( .A1(
        round_inst_sin_z[54]), .A2(round_inst_sin_y[55]), .A3(
        round_inst_S_13__sbox_inst_com_x_inst_n401), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n402) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U37 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n420), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n401) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U36 ( .A(
        round_inst_S_13__sbox_inst_n1), .B(round_inst_sin_w[53]), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n420) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U35 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n400), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n399), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n403) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U34 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n446), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n399) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U33 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n475), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n506), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U32 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n398), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n397), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n400) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U31 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n490), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n451), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n397) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n396), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n395), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U29 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n395) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U28 ( .A1(
        round_inst_sin_y[55]), .A2(round_inst_S_13__sbox_inst_com_x_inst_n392), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n393) );
  MUX2_X1 round_inst_S_13__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_13__sbox_inst_n1), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .S(round_inst_sin_w[54]), 
        .Z(round_inst_S_13__sbox_inst_com_x_inst_n392) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n391), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n394) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n451), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n390), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U24 ( .A1(round_inst_n58), 
        .A2(round_inst_sin_w[53]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n390) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U23 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_z[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n451) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U22 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n409), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n389), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n396) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U21 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n446), .Z(
        round_inst_S_13__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U20 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n388), .A2(round_inst_n58), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n446) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_13__sbox_inst_n1), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n388) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n387), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n386), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n514) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U17 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n385), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n419), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n386) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U16 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_z[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n419) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U15 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n384), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n385) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U14 ( .A(round_inst_sin_w[53]), .B(round_inst_S_13__sbox_inst_com_x_inst_n383), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n384) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_13__sbox_inst_n1), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_13__sbox_inst_com_x_inst_U12 ( .A(round_inst_sin_z[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n409) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n382), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n387) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_x_inst_U10 ( .A1(
        round_inst_sin_z[52]), .A2(round_inst_sin_y[55]), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n415) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U9 ( .A1(
        round_inst_S_13__sbox_inst_com_x_inst_n381), .A2(
        round_inst_S_13__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n382) );
  INV_X1 round_inst_S_13__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_y[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n462) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U7 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n506), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n380), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n381) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_x_inst_U6 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_13__sbox_inst_com_x_inst_n475), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n380) );
  INV_X1 round_inst_S_13__sbox_inst_com_x_inst_U5 ( .A(round_inst_sin_y[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n475) );
  INV_X1 round_inst_S_13__sbox_inst_com_x_inst_U4 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n476) );
  INV_X1 round_inst_S_13__sbox_inst_com_x_inst_U3 ( .A(round_inst_sin_y[53]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n408) );
  INV_X1 round_inst_S_13__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_13__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_13__sbox_inst_com_x_inst_n506) );
  INV_X1 round_inst_S_13__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_w[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_x_inst_n490) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n516), .Z(round_inst_sout_y[52])
         );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n515), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U134 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n513), .B(round_inst_sin_z[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n514) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U133 ( .A(round_inst_sin_x[48]), .B(round_inst_S_13__sbox_inst_com_y_inst_n512), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n515) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n511), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_srout2_y[22]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n507), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n517) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U129 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n506), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n505), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n507) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n505) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U127 ( .A1(
        round_inst_sin_w[54]), .A2(round_inst_sin_z[55]), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n506) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U125 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_13__sbox_inst_com_y_inst_U124 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_13__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U123 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_sin_x[55]), .A2(round_inst_S_13__sbox_inst_com_y_inst_n493), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U121 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n492), .A2(round_inst_sin_z[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U120 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U119 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U118 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U117 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n486), .A2(round_inst_sin_z[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U116 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_sin_w[54]), .A2(round_inst_sin_w[52]), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U114 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n513), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U112 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U111 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_13__sbox_inst_n1), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U109 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[51]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_y_inst_U108 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n513), .A2(round_inst_sin_z[55]), 
        .A3(round_inst_sin_x[52]), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U107 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_sin_w[52]), .A2(round_inst_sin_w[55]), .A3(
        round_inst_S_13__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_13__sbox_inst_com_y_inst_U105 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_13__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U104 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[20]) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U103 ( .A1(round_inst_n68), 
        .A2(round_inst_S_13__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n508) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U98 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U97 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_13__sbox_inst_n1), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_13__sbox_inst_com_y_inst_U95 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U94 ( .A1(
        round_inst_sin_x[52]), .A2(round_inst_sin_w[54]), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_y_inst_U93 ( .A1(
        round_inst_sin_w[52]), .A2(round_inst_S_13__sbox_inst_n3), .A3(
        round_inst_S_13__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U92 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U91 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n457), .A2(round_inst_n68), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U88 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U87 ( .A1(
        round_inst_S_13__sbox_inst_n1), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_13__sbox_inst_com_y_inst_U86 ( .A(round_inst_n68), .B(
        round_inst_sin_w[54]), .S(round_inst_S_13__sbox_inst_com_y_inst_n483), 
        .Z(round_inst_S_13__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U84 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U80 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_13__sbox_inst_n1), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U78 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n478), .B(round_inst_n67), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_sin_w[54]), .A2(round_inst_S_13__sbox_inst_com_y_inst_n483), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U76 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n513), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n438), .Z(
        round_inst_srout2_y[23]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U71 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U70 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U69 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n483), .A2(
        round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_13__sbox_inst_n1), .A2(round_inst_sin_w[52]), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_y_inst_U66 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[55]), 
        .A3(round_inst_S_13__sbox_inst_n1), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U65 ( .A(round_inst_sin_w[52]), 
        .B(round_inst_sin_x[52]), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U63 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U61 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U59 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U58 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U57 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[53]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U55 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_13__sbox_inst_com_y_inst_U54 ( .A(round_inst_sin_x[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U53 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n418), .A2(round_inst_sin_z[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U51 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U50 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U49 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n414), .B(
        round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U48 ( .A(round_inst_sin_w[53]), .B(round_inst_S_13__sbox_inst_n1), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_13__sbox_inst_n1), .A2(round_inst_sin_x[52]), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U46 ( .A1(
        round_inst_S_13__sbox_inst_n1), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U45 ( .A(round_inst_sin_x[50]), 
        .B(round_inst_S_13__sbox_inst_com_y_inst_n512), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U44 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n512) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U43 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U42 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U41 ( .A(round_inst_sin_w[53]), 
        .B(round_inst_sin_x[55]), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U40 ( .A(
        round_inst_S_13__sbox_inst_n3), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_13__sbox_inst_com_y_inst_U39 ( .A(round_inst_sin_w[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U38 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[52]), 
        .Z(round_inst_S_13__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_13__sbox_inst_com_y_inst_U36 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_13__sbox_inst_com_y_inst_U35 ( .A(round_inst_sin_z[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_13__sbox_inst_n1), .B(round_inst_sin_z[55]), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U30 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U29 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_13__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U27 ( .A(round_inst_n68), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_sin_w[53]), .A2(round_inst_sin_z[55]), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n513), .A2(round_inst_sin_w[53]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_13__sbox_inst_n1), .A2(round_inst_sin_w[55]), .A3(
        round_inst_n68), .ZN(round_inst_S_13__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U22 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_13__sbox_inst_n1), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U21 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U20 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n397) );
  INV_X1 round_inst_S_13__sbox_inst_com_y_inst_U19 ( .A(round_inst_sin_w[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n396) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n503), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U17 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_z[55]), .B(round_inst_sin_w[55]), .ZN(round_inst_S_13__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U15 ( .A(round_inst_sin_z[55]), 
        .B(round_inst_S_13__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n503) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U14 ( .A(round_inst_sin_w[55]), .B(round_inst_sin_x[55]), .ZN(round_inst_S_13__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U13 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U12 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_y_inst_U11 ( .A1(
        round_inst_S_13__sbox_inst_n3), .A2(round_inst_sin_w[55]), .A3(
        round_inst_S_13__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_y_inst_U10 ( .A1(
        round_inst_sin_z[55]), .A2(round_inst_S_13__sbox_inst_com_y_inst_n389), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_13__sbox_inst_com_y_inst_U9 ( .A(round_inst_sin_w[53]), 
        .B(round_inst_S_13__sbox_inst_n3), .S(round_inst_sin_w[54]), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_13__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_13__sbox_inst_n3), .A2(
        round_inst_S_13__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_13__sbox_inst_com_y_inst_n513), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U6 ( .A(round_inst_sin_z[55]), 
        .B(round_inst_sin_x[55]), .Z(
        round_inst_S_13__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_y_inst_U5 ( .A1(
        round_inst_S_13__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_13__sbox_inst_n1), .A3(round_inst_sin_x[55]), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_13__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_y_inst_U3 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n513), .B(round_inst_sin_w[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_13__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_13__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_13__sbox_inst_com_y_inst_n513) );
  INV_X1 round_inst_S_13__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U128 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n512), .ZN(round_inst_sout_z[52]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n511), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n510), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n513) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n509), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n508), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n511) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_sin_w[54]), .B(round_inst_sin_w[55]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n508) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U124 ( .A(round_inst_sin_x[48]), .B(round_inst_n56), .Z(round_inst_S_13__sbox_inst_com_z_inst_n509) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U123 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n510), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n507), .ZN(
        round_inst_srout2_z[22]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n506), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n505), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n504), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n503), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n505) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U120 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n502), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n501), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n503) );
  NOR3_X1 round_inst_S_13__sbox_inst_com_z_inst_U119 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n500), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n499), .A3(
        round_inst_S_13__sbox_inst_com_z_inst_n498), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n501) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U118 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n496), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n502) );
  INV_X1 round_inst_S_13__sbox_inst_com_z_inst_U117 ( .A(round_inst_sin_w[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n496) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U116 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n495), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n494), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n497) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U115 ( .A1(
        round_inst_sin_y[52]), .A2(round_inst_sin_x[55]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n494) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U114 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n493), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n492), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n495) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n491), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n490), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n506) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n489), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n488), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n490) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_z_inst_U111 ( .A1(round_inst_n68), 
        .A2(round_inst_sin_x[55]), .A3(round_inst_sin_w[52]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n488) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_sin_y[52]), .A2(round_inst_S_13__sbox_inst_com_z_inst_n487), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n489) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U109 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n486), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n491) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U108 ( .A(
        round_inst_sin_w[53]), .B(round_inst_sin_x[51]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U107 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n484), .B(round_inst_sin_y[51]), 
        .Z(round_inst_S_13__sbox_inst_com_z_inst_n486) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U106 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n482), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n484) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_z_inst_U105 ( .A1(round_inst_n58), 
        .A2(round_inst_S_13__sbox_inst_com_z_inst_n493), .A3(
        round_inst_sin_w[52]), .ZN(round_inst_S_13__sbox_inst_com_z_inst_n482)
         );
  NAND3_X1 round_inst_S_13__sbox_inst_com_z_inst_U104 ( .A1(
        round_inst_sin_x[52]), .A2(round_inst_sin_w[55]), .A3(
        round_inst_S_13__sbox_inst_com_z_inst_n481), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n483) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n479), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n510) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n487), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n478), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n479) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U101 ( .A1(
        round_inst_sin_w[54]), .A2(round_inst_S_13__sbox_inst_com_z_inst_n493), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U100 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n478), .ZN(
        round_inst_srout2_z[20]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U99 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n476), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n478) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U98 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n474), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n475) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U97 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n472), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n471), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n473) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U96 ( .A1(round_inst_n68), 
        .A2(round_inst_S_13__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n471) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U95 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n469), .A2(round_inst_n58), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n472) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U94 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n468), .A2(round_inst_sin_w[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n474) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n467), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n466), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n465), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n464), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U91 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n463), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n462), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U90 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n461), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n460), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n462) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U89 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n470), .A2(round_inst_n58), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n460) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U88 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n459), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n458), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n461) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U87 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U85 ( .A1(
        round_inst_sin_w[54]), .A2(round_inst_sin_w[53]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n454) );
  AND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U84 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n466), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n481), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n455) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U83 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n453), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n451), .A2(round_inst_n68), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n452) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U81 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n451) );
  INV_X1 round_inst_S_13__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n469) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U79 ( .A1(
        round_inst_sin_y[52]), .A2(round_inst_sin_w[53]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U78 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n448), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n453) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U77 ( .A(round_inst_sin_x[52]), .B(round_inst_sin_y[52]), .ZN(round_inst_S_13__sbox_inst_com_z_inst_n448) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U76 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n446), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n477) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U75 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n481), .A2(round_inst_sin_w[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n443), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n443) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U72 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n492), .A2(round_inst_sin_w[54]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n441) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U71 ( .A(round_inst_sin_y[49]), 
        .B(round_inst_n67), .Z(round_inst_S_13__sbox_inst_com_z_inst_n442) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U70 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n440), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_srout2_z[23]) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U69 ( .A(round_inst_sin_w[52]), .B(round_inst_sin_x[50]), .ZN(round_inst_S_13__sbox_inst_com_z_inst_n439) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U68 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n438), .B(round_inst_n57), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n512), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n438) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U66 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n504), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n437) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U65 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n436), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n435), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U64 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n435) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U63 ( .A1(
        round_inst_sin_y[55]), .A2(round_inst_S_13__sbox_inst_com_z_inst_n466), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U62 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n434) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U61 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n430), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n430) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U59 ( .A1(
        round_inst_S_13__sbox_inst_n3), .A2(round_inst_sin_y[52]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U58 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n466), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n426), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n428) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U57 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n499), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n425), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n466) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U56 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n424), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n492), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n432) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U55 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n422), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n424) );
  AND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U54 ( .A1(round_inst_sin_w[53]), .A2(round_inst_sin_x[55]), .ZN(round_inst_S_13__sbox_inst_com_z_inst_n423)
         );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U53 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n436) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U52 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n419), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n418), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U51 ( .A1(
        round_inst_sin_y[55]), .A2(round_inst_S_13__sbox_inst_com_z_inst_n417), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n418) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U50 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n417) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U49 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n426), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n416), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n470) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U48 ( .A1(
        round_inst_sin_y[53]), .A2(round_inst_sin_w[52]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n416) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_z_inst_U47 ( .A1(
        round_inst_sin_w[53]), .A2(round_inst_sin_y[52]), .A3(
        round_inst_sin_x[55]), .ZN(round_inst_S_13__sbox_inst_com_z_inst_n419)
         );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U46 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n414), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n421) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n465), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n414) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U44 ( .A1(
        round_inst_sin_y[53]), .A2(round_inst_S_13__sbox_inst_com_z_inst_n492), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n465) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U43 ( .A(round_inst_sin_w[52]), 
        .B(round_inst_sin_x[52]), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n492) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U42 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n413), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n499), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n415) );
  INV_X1 round_inst_S_13__sbox_inst_com_z_inst_U41 ( .A(round_inst_sin_w[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n499) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U39 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U38 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n487), .A2(round_inst_sin_y[53]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n409) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n407), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n407) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U35 ( .A1(
        round_inst_sin_y[55]), .A2(round_inst_S_13__sbox_inst_com_z_inst_n459), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n405) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U34 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n404), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n403), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n406) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n402), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n401), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n403) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U32 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n487), .A2(
        round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n401) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U31 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n498), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n487) );
  INV_X1 round_inst_S_13__sbox_inst_com_z_inst_U30 ( .A(round_inst_sin_w[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n429) );
  MUX2_X1 round_inst_S_13__sbox_inst_com_z_inst_U29 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n413), .S(round_inst_sin_w[54]), 
        .Z(round_inst_S_13__sbox_inst_com_z_inst_n402) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_sin_x[55]), .A2(round_inst_S_13__sbox_inst_com_z_inst_n399), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n413) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U27 ( .A(round_inst_sin_y[53]), 
        .B(round_inst_S_13__sbox_inst_n3), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U26 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n493), .A2(round_inst_sin_w[53]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n400) );
  NAND3_X1 round_inst_S_13__sbox_inst_com_z_inst_U25 ( .A1(
        round_inst_sin_w[53]), .A2(round_inst_S_13__sbox_inst_com_z_inst_n481), 
        .A3(round_inst_sin_x[55]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n404) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U24 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n498), .B(round_inst_n58), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U23 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n398), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_sin_y[55]), .A2(round_inst_S_13__sbox_inst_com_z_inst_n456), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n397) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U21 ( .A1(round_inst_n58), 
        .A2(round_inst_S_13__sbox_inst_com_z_inst_n422), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n398) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U20 ( .A1(
        round_inst_S_13__sbox_inst_n3), .A2(round_inst_sin_w[55]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U19 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n396), .A2(round_inst_sin_w[55]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U18 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n456), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n459), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n396) );
  XOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U17 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n447), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n395), .Z(
        round_inst_S_13__sbox_inst_com_z_inst_n459) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U16 ( .A1(
        round_inst_sin_w[53]), .A2(round_inst_n58), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n395) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U15 ( .A1(
        round_inst_sin_w[54]), .A2(round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n447) );
  NOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U14 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n425), .A2(
        round_inst_S_13__sbox_inst_com_z_inst_n498), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n456) );
  INV_X1 round_inst_S_13__sbox_inst_com_z_inst_U13 ( .A(round_inst_n68), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n498) );
  INV_X1 round_inst_S_13__sbox_inst_com_z_inst_U12 ( .A(round_inst_sin_w[53]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n425) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U11 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n394), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n393), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U10 ( .A1(
        round_inst_S_13__sbox_inst_com_z_inst_n392), .A2(round_inst_sin_w[52]), 
        .ZN(round_inst_S_13__sbox_inst_com_z_inst_n393) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U9 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n391), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n392) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U8 ( .A(round_inst_sin_x[55]), 
        .B(round_inst_S_13__sbox_inst_com_z_inst_n500), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n493) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U7 ( .A(round_inst_sin_w[55]), 
        .B(round_inst_sin_y[55]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n500) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U6 ( .A(round_inst_sin_w[53]), 
        .B(round_inst_sin_y[53]), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n391) );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U5 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n464), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n390), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n394) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U4 ( .A1(round_inst_sin_x[52]), .A2(round_inst_sin_w[55]), .ZN(round_inst_S_13__sbox_inst_com_z_inst_n390)
         );
  XNOR2_X1 round_inst_S_13__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_13__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_13__sbox_inst_com_z_inst_n426), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U2 ( .A1(round_inst_sin_x[52]), .A2(round_inst_sin_w[53]), .ZN(round_inst_S_13__sbox_inst_com_z_inst_n426)
         );
  NAND2_X1 round_inst_S_13__sbox_inst_com_z_inst_U1 ( .A1(round_inst_sin_w[52]), .A2(round_inst_S_13__sbox_inst_n3), .ZN(
        round_inst_S_13__sbox_inst_com_z_inst_n449) );
  INV_X1 round_inst_S_14__sbox_inst_U6 ( .A(round_inst_sin_x[58]), .ZN(
        round_inst_S_14__sbox_inst_n6) );
  INV_X1 round_inst_S_14__sbox_inst_U5 ( .A(round_inst_sin_z[57]), .ZN(
        round_inst_S_14__sbox_inst_n2) );
  INV_X1 round_inst_S_14__sbox_inst_U4 ( .A(round_inst_sin_z[59]), .ZN(
        round_inst_S_14__sbox_inst_n4) );
  INV_X2 round_inst_S_14__sbox_inst_U3 ( .A(round_inst_S_14__sbox_inst_n4), 
        .ZN(round_inst_S_14__sbox_inst_n3) );
  INV_X2 round_inst_S_14__sbox_inst_U2 ( .A(round_inst_S_14__sbox_inst_n2), 
        .ZN(round_inst_S_14__sbox_inst_n1) );
  INV_X2 round_inst_S_14__sbox_inst_U1 ( .A(round_inst_S_14__sbox_inst_n6), 
        .ZN(round_inst_S_14__sbox_inst_n5) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n529), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n528), .ZN(round_inst_sout_w[59]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n526), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n528) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U136 ( .A1(
        round_inst_sin_z[56]), .A2(round_inst_S_14__sbox_inst_com_w_inst_n525), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n526) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n524), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n523), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n523) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U133 ( .A1(
        round_inst_sin_z[58]), .A2(round_inst_S_14__sbox_inst_com_w_inst_n520), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n521) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U132 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n519), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n518), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n520) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n517), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n516), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n522) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n515), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n514), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n516) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U129 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n518), .A2(
        round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U128 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n513), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n512), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U127 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n511), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n512) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U126 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n508), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n510) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_w_inst_U125 ( .A1(
        round_inst_S_14__sbox_inst_n5), .A2(round_inst_sin_x[56]), .A3(
        round_inst_S_14__sbox_inst_com_w_inst_n507), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n508) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n506), .A2(round_inst_n59), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n509) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U123 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n505), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n511) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U122 ( .A(
        round_inst_sin_x[59]), .B(round_inst_S_14__sbox_inst_com_w_inst_n503), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n505) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_w_inst_U121 ( .A1(
        round_inst_S_14__sbox_inst_n3), .A2(round_inst_n60), .A3(
        round_inst_sin_x[56]), .ZN(round_inst_S_14__sbox_inst_com_w_inst_n513)
         );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U120 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n502), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n501), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_sin_y[55]), .B(round_inst_S_14__sbox_inst_com_w_inst_n500), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n501) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U118 ( .A(round_inst_n69), .B(
        round_inst_sin_z[55]), .Z(round_inst_S_14__sbox_inst_com_w_inst_n500)
         );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U117 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n499), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n502) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_sin_x[59]), .B(round_inst_sin_y[59]), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n499) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[57]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U113 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[53]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[53]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U110 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[56]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_14__sbox_inst_n5), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n529), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U105 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n529) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U104 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U102 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_14__sbox_inst_n5), .B(round_inst_sin_z[58]), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U99 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_14__sbox_inst_n1), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n504), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U96 ( .A1(round_inst_n60), 
        .A2(round_inst_sin_x[56]), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n498) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U95 ( .A1(
        round_inst_S_14__sbox_inst_n5), .A2(round_inst_n59), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n504) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U94 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U93 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_z[58]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U90 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U89 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U88 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n461), .A2(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n460), .B(round_inst_sin_z[58]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U86 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U85 ( .A1(round_inst_sin_z[56]), .A2(round_inst_S_14__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U84 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_sin_y[57]), .A2(round_inst_n59), .A3(
        round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_w_inst_U81 ( .A1(round_inst_n60), 
        .A2(round_inst_n69), .A3(round_inst_n59), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U80 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n525) );
  OR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U79 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_14__sbox_inst_n5), .B(round_inst_n60), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U77 ( .A(round_inst_sin_y[52]), 
        .B(round_inst_sin_z[52]), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n484) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[59])
         );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U73 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U71 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_14__sbox_inst_n3), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U69 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U68 ( .A1(round_inst_n60), 
        .A2(round_inst_n69), .ZN(round_inst_S_14__sbox_inst_com_w_inst_n456)
         );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_14__sbox_inst_n5), .A2(round_inst_sin_y[57]), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U66 ( .A1(
        round_inst_S_14__sbox_inst_n1), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_w_inst_U65 ( .A1(
        round_inst_S_14__sbox_inst_n5), .A2(round_inst_S_14__sbox_inst_n1), 
        .A3(round_inst_sin_x[59]), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n439), .A2(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U62 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U61 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n503), .A2(
        round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U60 ( .A(
        round_inst_S_14__sbox_inst_n3), .B(round_inst_sin_y[59]), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n503) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n506) );
  INV_X1 round_inst_S_14__sbox_inst_com_w_inst_U58 ( .A(round_inst_sin_x[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n486) );
  INV_X1 round_inst_S_14__sbox_inst_com_w_inst_U57 ( .A(round_inst_n60), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U56 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U55 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U54 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U52 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U51 ( .A(round_inst_sin_y[57]), .B(round_inst_S_14__sbox_inst_n1), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U50 ( .A1(
        round_inst_S_14__sbox_inst_n3), .A2(round_inst_S_14__sbox_inst_n1), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U49 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U48 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_w_inst_U47 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n425), .A2(round_inst_sin_x[59]), 
        .A3(round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U46 ( .A(round_inst_sin_y[57]), 
        .B(round_inst_n69), .Z(round_inst_S_14__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_w_inst_U45 ( .A1(
        round_inst_sin_x[59]), .A2(round_inst_sin_y[57]), .A3(
        round_inst_S_14__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U44 ( .A(round_inst_n60), .B(
        round_inst_sin_z[58]), .ZN(round_inst_S_14__sbox_inst_com_w_inst_n465)
         );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U43 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U42 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n517) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U41 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n421), .A2(
        round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U40 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n419), .A2(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U38 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U37 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U36 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n518), .A2(
        round_inst_S_14__sbox_inst_n1), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U35 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n518) );
  INV_X1 round_inst_S_14__sbox_inst_com_w_inst_U34 ( .A(round_inst_sin_x[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n489) );
  INV_X1 round_inst_S_14__sbox_inst_com_w_inst_U33 ( .A(round_inst_sin_y[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n434) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U32 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U31 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U30 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U29 ( .A(round_inst_sin_x[56]), .B(round_inst_sin_z[56]), .ZN(round_inst_S_14__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U28 ( .A1(
        round_inst_sin_y[59]), .A2(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U27 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U26 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n407), .A2(round_inst_sin_y[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U24 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n466), .A2(round_inst_sin_x[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U23 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U22 ( .A1(round_inst_n69), 
        .A2(round_inst_sin_z[56]), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U21 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_14__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U20 ( .A(round_inst_n69), .B(
        round_inst_S_14__sbox_inst_n1), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U19 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n404), .A2(round_inst_sin_x[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U17 ( .A1(
        round_inst_sin_x[56]), .A2(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U16 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n418), .A2(round_inst_sin_y[57]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U15 ( .A(round_inst_n59), .B(
        round_inst_sin_z[56]), .Z(round_inst_S_14__sbox_inst_com_w_inst_n418)
         );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U13 ( .A(round_inst_sin_x[56]), .B(round_inst_S_14__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U11 ( .A1(
        round_inst_S_14__sbox_inst_com_w_inst_n398), .A2(round_inst_sin_x[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U9 ( .A(round_inst_sin_y[59]), 
        .B(round_inst_n69), .ZN(round_inst_S_14__sbox_inst_com_w_inst_n396) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U8 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_14__sbox_inst_n1), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U7 ( .A(
        round_inst_S_14__sbox_inst_n3), .B(round_inst_sin_x[59]), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n507) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U6 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n519), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_14__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U5 ( .A(
        round_inst_S_14__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_14__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_14__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U4 ( .A1(round_inst_n69), 
        .A2(round_inst_n59), .ZN(round_inst_S_14__sbox_inst_com_w_inst_n475)
         );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U3 ( .A1(round_inst_sin_x[56]), .A2(round_inst_sin_y[57]), .ZN(round_inst_S_14__sbox_inst_com_w_inst_n477)
         );
  NAND2_X1 round_inst_S_14__sbox_inst_com_w_inst_U2 ( .A1(round_inst_sin_x[59]), .A2(round_inst_n59), .ZN(round_inst_S_14__sbox_inst_com_w_inst_n519) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_w_inst_U1 ( .A(round_inst_n58), .B(
        round_inst_sin_z[54]), .Z(round_inst_S_14__sbox_inst_com_w_inst_n402)
         );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U136 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n512), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n511), .ZN(round_inst_sout_x[56]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n510), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n509), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n511) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U134 ( .A(round_inst_n60), 
        .B(round_inst_S_14__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U133 ( .A(round_inst_sin_z[52]), .B(round_inst_S_14__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n510) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U132 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n512), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n506), .Z(
        round_inst_srout2_x[42]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U130 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n503), .A2(round_inst_sin_z[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U129 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U127 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U126 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U125 ( .A1(round_inst_n60), 
        .A2(round_inst_sin_w[56]), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n496) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U124 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U122 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U121 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U118 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n508), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U117 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n487) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U115 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n481) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_x_inst_U114 ( .A1(
        round_inst_sin_z[58]), .A2(round_inst_sin_w[56]), .A3(
        round_inst_S_14__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n489) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n478), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n475), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n477) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n474), .B(round_inst_sin_z[55]), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n475) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_w[58]), .A2(round_inst_S_14__sbox_inst_com_x_inst_n508), 
        .A3(round_inst_sin_z[56]), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n473), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n478) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n470), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n473) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n469), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n468), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n512) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n467), .A2(round_inst_n60), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n468) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n467) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n469) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n465), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n463), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_srout2_x[40]) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U100 ( .A1(round_inst_n59), 
        .A2(round_inst_sin_z[58]), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[53]), .B(round_inst_S_14__sbox_inst_com_x_inst_n462), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n461), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n462) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n466), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n460) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n458), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n457), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_14__sbox_inst_n1), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n459), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n456), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n455), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n454), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n453), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n455) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n452), .A2(round_inst_sin_w[58]), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n451), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n450), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n454) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n449), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n448), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n447), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n446), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n448) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n445), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n446) );
  MUX2_X1 round_inst_S_14__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n444), .B(round_inst_n60), .S(
        round_inst_n59), .Z(round_inst_S_14__sbox_inst_com_x_inst_n445) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n443), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_14__sbox_inst_com_x_inst_U85 ( .A(round_inst_n60), .B(
        round_inst_sin_z[58]), .S(round_inst_sin_z[56]), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n443) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n442), .A2(round_inst_sin_w[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n449) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n441), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n440), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n451) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_w[56]), 
        .A3(round_inst_sin_z[58]), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n440) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n439), .A2(round_inst_sin_w[57]), 
        .A3(round_inst_n60), .ZN(round_inst_S_14__sbox_inst_com_x_inst_n441)
         );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U80 ( .A(round_inst_n59), .B(
        round_inst_sin_z[56]), .Z(round_inst_S_14__sbox_inst_com_x_inst_n439)
         );
  NAND3_X1 round_inst_S_14__sbox_inst_com_x_inst_U79 ( .A1(round_inst_n59), 
        .A2(round_inst_S_14__sbox_inst_com_x_inst_n444), .A3(
        round_inst_S_14__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n456) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n459) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U77 ( .A1(round_inst_n59), 
        .A2(round_inst_n60), .ZN(round_inst_S_14__sbox_inst_com_x_inst_n482)
         );
  AND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U76 ( .A1(round_inst_n60), 
        .A2(round_inst_sin_z[56]), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n490) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n461) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U74 ( .A1(round_inst_n59), 
        .A2(round_inst_sin_w[58]), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n497) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n436), .ZN(
        round_inst_srout2_x[43]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n435), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n434), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n436) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U71 ( .A(round_inst_n59), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n434) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n433), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n432), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U69 ( .A1(
        round_inst_sin_z[56]), .A2(round_inst_S_14__sbox_inst_com_x_inst_n508), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n432) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n431), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n430), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n433) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n429), .A2(round_inst_n59), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n428), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n476), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n427) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_14__sbox_inst_n1), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n431) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n452) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[54]), 
        .B(round_inst_S_14__sbox_inst_com_x_inst_n437), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n435) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n424), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n423), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n422), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n421), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n423) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n420), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n419), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n421) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n418), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n419) );
  NOR3_X1 round_inst_S_14__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n470), .A3(
        round_inst_S_14__sbox_inst_com_x_inst_n416), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n417) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n415), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n414), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n418) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n413), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n414) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U53 ( .A1(round_inst_n60), 
        .A2(round_inst_S_14__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n412) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U52 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n442), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_14__sbox_inst_n1), .A2(round_inst_n60), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n442) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_x_inst_U50 ( .A1(round_inst_n60), 
        .A2(round_inst_S_14__sbox_inst_com_x_inst_n476), .A3(
        round_inst_S_14__sbox_inst_com_x_inst_n411), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n420) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U49 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n410), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n464), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n422) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U48 ( .A1(round_inst_n60), 
        .A2(round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n464) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U47 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n410) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n409), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n408), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n407), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n406), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n405), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n404), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n406) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U43 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n465), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n404) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U42 ( .A(round_inst_sin_w[57]), 
        .B(round_inst_S_14__sbox_inst_n1), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n438) );
  AND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U41 ( .A1(round_inst_sin_z[58]), .A2(round_inst_S_14__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n465) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U40 ( .A1(
        round_inst_S_14__sbox_inst_n3), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n405) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n444), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n476), .A3(
        round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n407) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U38 ( .A(round_inst_sin_z[58]), 
        .B(round_inst_sin_w[58]), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U37 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n403), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n402), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U36 ( .A(round_inst_sin_w[58]), 
        .B(round_inst_n60), .Z(round_inst_S_14__sbox_inst_com_x_inst_n402) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U35 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n401), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n400), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n399), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n400) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U33 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n425), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n398) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U32 ( .A1(
        round_inst_sin_z[56]), .A2(round_inst_S_14__sbox_inst_com_x_inst_n476), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n425) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U31 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n479), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n471) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_14__sbox_inst_n3), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n426), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n470), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n399) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U28 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n401) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_14__sbox_inst_n1), .A3(round_inst_n59), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n396) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n508), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n411), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U23 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n392), .A2(round_inst_sin_w[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U21 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_x_inst_U19 ( .A1(
        round_inst_sin_z[56]), .A2(round_inst_S_14__sbox_inst_com_x_inst_n508), 
        .A3(round_inst_sin_w[57]), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n388) );
  MUX2_X1 round_inst_S_14__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n411), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n508), .S(
        round_inst_S_14__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U17 ( .A1(round_inst_n59), 
        .A2(round_inst_S_14__sbox_inst_com_x_inst_n476), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n491), .B(
        round_inst_S_14__sbox_inst_n3), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n411) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U15 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U14 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n384), .A2(round_inst_sin_z[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n403), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n476), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U10 ( .A(round_inst_sin_w[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U9 ( .A1(
        round_inst_S_14__sbox_inst_n1), .A2(
        round_inst_S_14__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n403) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U8 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n508) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U7 ( .A(round_inst_sin_y[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n413) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_14__sbox_inst_com_x_inst_n426), .Z(
        round_inst_S_14__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U4 ( .A1(round_inst_n59), 
        .A2(round_inst_sin_w[57]), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n426) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_14__sbox_inst_com_x_inst_n476), .A2(round_inst_sin_w[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_14__sbox_inst_com_x_inst_n416), .ZN(
        round_inst_S_14__sbox_inst_com_x_inst_n476) );
  INV_X1 round_inst_S_14__sbox_inst_com_x_inst_U1 ( .A(round_inst_sin_y[57]), 
        .ZN(round_inst_S_14__sbox_inst_com_x_inst_n416) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U138 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n519), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n518), .Z(round_inst_sout_y[56])
         );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n517), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n516), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n518) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n515), .B(
        round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n516) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U135 ( .A(round_inst_sin_x[52]), .B(round_inst_S_14__sbox_inst_com_y_inst_n514), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U134 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n513), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n512), .ZN(
        round_inst_srout2_y[42]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n519), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n510), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n509), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n519) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n508), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n507), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n509) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U130 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n506), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n507) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n508) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U128 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n503), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n502), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n513) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n501), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n500), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n502) );
  NOR3_X1 round_inst_S_14__sbox_inst_com_y_inst_U126 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n499), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n498), .A3(
        round_inst_S_14__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n500) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U125 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n496), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n495), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n501) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U124 ( .A1(
        round_inst_sin_x[59]), .A2(round_inst_S_14__sbox_inst_com_y_inst_n494), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n495) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U123 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n493), .A2(
        round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U122 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n492), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n491), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U121 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n490), .A2(round_inst_sin_w[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n492) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U120 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n489), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n488), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n503) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U119 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n487), .A2(
        round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n488) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U118 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n486), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n485), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n487) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U117 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n504), .A2(round_inst_sin_w[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n485) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n515), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n486) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U115 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n482), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n489) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n481), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n480), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n482) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U113 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n479), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U112 ( .A(
        round_inst_S_14__sbox_inst_n1), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n478), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n481) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n477), .B(round_inst_sin_x[55]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n478) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_y_inst_U110 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n515), .A2(
        round_inst_S_14__sbox_inst_n3), .A3(
        round_inst_S_14__sbox_inst_com_y_inst_n476), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n477) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U109 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n483) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_y_inst_U108 ( .A1(
        round_inst_sin_w[56]), .A2(round_inst_sin_w[59]), .A3(
        round_inst_S_14__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_14__sbox_inst_com_y_inst_U107 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n506), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_14__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U106 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[40]) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U105 ( .A1(
        round_inst_S_14__sbox_inst_n5), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U104 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n510), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U99 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_14__sbox_inst_n1), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U98 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U96 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n476), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n491) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_y_inst_U95 ( .A1(
        round_inst_sin_w[56]), .A2(round_inst_n69), .A3(
        round_inst_S_14__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U94 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U93 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U92 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U89 ( .A1(
        round_inst_S_14__sbox_inst_n1), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_14__sbox_inst_com_y_inst_U88 ( .A(
        round_inst_S_14__sbox_inst_n5), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n504), .S(
        round_inst_S_14__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U87 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U85 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U81 ( .A(
        round_inst_S_14__sbox_inst_n1), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n479), .B(round_inst_sin_x[53]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U79 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n504), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n479) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n515), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U77 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n438), .Z(
        round_inst_srout2_y[43]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n484), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U72 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U71 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U70 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n484), .A2(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_14__sbox_inst_n1), .A2(round_inst_sin_w[56]), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n443), .A2(round_inst_sin_x[59]), 
        .A3(round_inst_S_14__sbox_inst_n1), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U67 ( .A(round_inst_sin_w[56]), 
        .B(round_inst_S_14__sbox_inst_com_y_inst_n476), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U66 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U64 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U62 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U60 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U59 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U58 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n484), .A2(round_inst_sin_w[57]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n422) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n418), .A2(
        round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U55 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U54 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U53 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n414), .B(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U51 ( .A(round_inst_sin_w[57]), .B(round_inst_S_14__sbox_inst_n1), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U50 ( .A1(
        round_inst_S_14__sbox_inst_n1), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n476), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n444) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U49 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n473), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n476) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U48 ( .A(round_inst_sin_x[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_14__sbox_inst_n1), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n484), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U46 ( .A(round_inst_n68), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n514), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n514) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[57]), 
        .B(round_inst_sin_x[59]), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U41 ( .A(round_inst_n69), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n499) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n484), .B(round_inst_sin_w[56]), 
        .Z(round_inst_S_14__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n484) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U36 ( .A(round_inst_sin_z[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n497) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_14__sbox_inst_n1), .B(round_inst_S_14__sbox_inst_n3), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n490), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n498) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_14__sbox_inst_n5), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n506), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n490) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U27 ( .A1(
        round_inst_sin_w[57]), .A2(round_inst_S_14__sbox_inst_n3), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n515), .A2(round_inst_sin_w[57]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_14__sbox_inst_n1), .A2(round_inst_sin_w[59]), .A3(
        round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_14__sbox_inst_n1), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n505), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n506), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_14__sbox_inst_n3), .B(round_inst_sin_w[59]), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U17 ( .A(
        round_inst_S_14__sbox_inst_n3), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[59]), .B(round_inst_sin_x[59]), .ZN(round_inst_S_14__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_y_inst_U13 ( .A1(round_inst_n69), 
        .A2(round_inst_sin_w[59]), .A3(
        round_inst_S_14__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_y_inst_U12 ( .A1(
        round_inst_S_14__sbox_inst_n3), .A2(
        round_inst_S_14__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_14__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[57]), 
        .B(round_inst_n69), .S(round_inst_S_14__sbox_inst_com_y_inst_n504), 
        .Z(round_inst_S_14__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_y_inst_U9 ( .A1(round_inst_n69), 
        .A2(round_inst_S_14__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_14__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_14__sbox_inst_n3), .B(round_inst_sin_x[59]), .Z(
        round_inst_S_14__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_14__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_14__sbox_inst_n1), .A3(round_inst_sin_x[59]), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n515), .B(
        round_inst_S_14__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n504) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[58]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_14__sbox_inst_com_y_inst_n506), .ZN(
        round_inst_S_14__sbox_inst_com_y_inst_n515) );
  INV_X1 round_inst_S_14__sbox_inst_com_y_inst_U1 ( .A(round_inst_sin_z[58]), 
        .ZN(round_inst_S_14__sbox_inst_com_y_inst_n506) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U132 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n517), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n516), .ZN(round_inst_sout_z[56]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n515), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n514), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_sin_w[58]), .B(round_inst_sin_w[59]), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n514) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_x[52]), .B(round_inst_sin_y[52]), .Z(round_inst_S_14__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U128 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n512), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n517) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_srout2_z[42]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n510), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n509), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n511) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n508), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n507), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n509) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U124 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n506), .A2(round_inst_n59), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U123 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n505), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n504), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n508) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n503), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n502), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_sin_w[57]), .B(round_inst_sin_x[55]), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U120 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n501), .B(round_inst_sin_y[55]), 
        .Z(round_inst_S_14__sbox_inst_com_z_inst_n503) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U119 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n500), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n499), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n501) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U118 ( .A1(round_inst_n60), 
        .A2(round_inst_S_14__sbox_inst_com_z_inst_n498), .A3(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n499) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U117 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n496), .A2(round_inst_sin_x[56]), 
        .A3(round_inst_sin_w[59]), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n500) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U116 ( .A(
        round_inst_S_14__sbox_inst_n5), .B(round_inst_n60), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n496) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U115 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_14__sbox_inst_n5), .A3(
        round_inst_S_14__sbox_inst_com_z_inst_n495), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n505) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U114 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n493), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n492), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n491), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n493) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n490), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n489), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n491) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U111 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n488), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n489) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n486), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n490) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_sin_w[58]), .A2(round_inst_S_14__sbox_inst_com_z_inst_n495), 
        .A3(round_inst_n59), .ZN(round_inst_S_14__sbox_inst_com_z_inst_n492)
         );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U108 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n484), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n485), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n513) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U107 ( .A1(
        round_inst_sin_w[58]), .A2(round_inst_S_14__sbox_inst_com_z_inst_n498), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U106 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n506), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n484) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n482), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n481), .Z(
        round_inst_srout2_z[40]) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n480), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n479), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n478), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n483), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n477), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n483) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U101 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n475), .A2(round_inst_sin_x[56]), 
        .A3(round_inst_sin_w[58]), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n476) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U100 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n474), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n473), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n477) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U99 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n472), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .A3(round_inst_n60), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n473) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U98 ( .A(round_inst_sin_w[57]), 
        .B(round_inst_sin_y[57]), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U97 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n471), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n474) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U96 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n469), .A2(
        round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n470) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U95 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n468), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n467), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n471) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n466), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n465), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n464), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n463), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n465) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n462), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n461), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n463) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U91 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n460), .A2(round_inst_n60), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n461) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U90 ( .A1(round_inst_n69), 
        .A2(round_inst_S_14__sbox_inst_n5), .A3(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n462) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U89 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n459), .A2(round_inst_n59), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_w[58]), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n466) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U87 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U85 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n453), .A2(round_inst_n60), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n454) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U84 ( .A(round_inst_sin_w[57]), .B(round_inst_S_14__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U83 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n451), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_sin_w[58]), .A2(round_inst_sin_x[56]), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n478) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U81 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n487), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n448) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U79 ( .A(round_inst_sin_y[53]), 
        .B(round_inst_sin_x[53]), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n447) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U78 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n487) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n446), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U76 ( .A(round_inst_sin_w[58]), .B(round_inst_n60), .ZN(round_inst_S_14__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U75 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_srout2_z[43]) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n494), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n512), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U72 ( .A1(
        round_inst_sin_x[56]), .A2(round_inst_sin_w[59]), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n441) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U71 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n458), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n440), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n442) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U70 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n498), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U69 ( .A(round_inst_sin_w[59]), .B(round_inst_S_14__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n498) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U68 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n494) );
  MUX2_X1 round_inst_S_14__sbox_inst_com_z_inst_U67 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n495), .B(round_inst_sin_w[59]), 
        .S(round_inst_S_14__sbox_inst_com_z_inst_n436), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n437) );
  OR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U66 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n436) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U65 ( .A(round_inst_sin_x[56]), .B(round_inst_S_14__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n486) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U64 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n438) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U63 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n495), .A3(
        round_inst_S_14__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U62 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n430), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n429) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U59 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n426), .A2(round_inst_sin_w[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U58 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n422), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n424) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U56 ( .A1(
        round_inst_sin_x[56]), .A2(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U55 ( .A1(
        round_inst_sin_y[57]), .A2(round_inst_sin_x[56]), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n425) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U54 ( .A1(round_inst_n59), 
        .A2(round_inst_S_14__sbox_inst_com_z_inst_n495), .A3(
        round_inst_sin_w[57]), .ZN(round_inst_S_14__sbox_inst_com_z_inst_n428)
         );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U53 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_y[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U52 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n469), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n460), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n423), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n469) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U50 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .A2(round_inst_sin_y[57]), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n423) );
  AND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U49 ( .A1(round_inst_sin_w[57]), .A2(round_inst_sin_x[56]), .ZN(round_inst_S_14__sbox_inst_com_z_inst_n460)
         );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U48 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n421) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U47 ( .A1(
        round_inst_sin_w[57]), .A2(round_inst_S_14__sbox_inst_com_z_inst_n497), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U46 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .A2(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n419), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n418), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n432) );
  INV_X1 round_inst_S_14__sbox_inst_com_z_inst_U44 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U43 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .B(round_inst_n59), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n451) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n417), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U41 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n497), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n449) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U39 ( .A1(
        round_inst_sin_w[59]), .A2(round_inst_S_14__sbox_inst_com_z_inst_n413), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n414) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U38 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n415) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U35 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n506), .A2(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n409) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U34 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n407) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U32 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n405) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n404) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U30 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n506), .A2(round_inst_sin_y[57]), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n402) );
  AND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_S_14__sbox_inst_n5), .A2(round_inst_sin_w[59]), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n506) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n401), .A2(round_inst_n60), .A3(
        round_inst_sin_w[57]), .ZN(round_inst_S_14__sbox_inst_com_z_inst_n403)
         );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U27 ( .A(round_inst_sin_w[59]), 
        .B(round_inst_S_14__sbox_inst_com_z_inst_n495), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n401) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U26 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n399), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n406) );
  MUX2_X1 round_inst_S_14__sbox_inst_com_z_inst_U25 ( .A(round_inst_sin_y[59]), 
        .B(round_inst_S_14__sbox_inst_com_z_inst_n398), .S(
        round_inst_S_14__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U24 ( .A1(
        round_inst_sin_w[57]), .A2(round_inst_S_14__sbox_inst_n5), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U23 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n398) );
  NOR3_X1 round_inst_S_14__sbox_inst_com_z_inst_U22 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n488), .A3(
        round_inst_S_14__sbox_inst_com_z_inst_n395), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U21 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n394), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n395) );
  INV_X1 round_inst_S_14__sbox_inst_com_z_inst_U20 ( .A(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n394) );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U19 ( .A(round_inst_sin_w[59]), .B(round_inst_sin_y[59]), .ZN(round_inst_S_14__sbox_inst_com_z_inst_n488) );
  AND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U18 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n459), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U17 ( .A1(
        round_inst_sin_w[58]), .A2(round_inst_n69), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n459) );
  INV_X1 round_inst_S_14__sbox_inst_com_z_inst_U16 ( .A(round_inst_sin_w[57]), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U15 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n393), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U14 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n391), .A2(round_inst_n60), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U13 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_14__sbox_inst_com_z_inst_n390), .Z(
        round_inst_S_14__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U12 ( .A1(
        round_inst_sin_w[57]), .A2(round_inst_sin_y[59]), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n390) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U11 ( .A1(round_inst_n69), 
        .A2(round_inst_sin_w[59]), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n418) );
  NOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U10 ( .A1(
        round_inst_S_14__sbox_inst_com_z_inst_n439), .A2(
        round_inst_S_14__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_14__sbox_inst_com_z_inst_U9 ( .A1(round_inst_sin_w[58]), .A2(round_inst_sin_w[57]), .ZN(round_inst_S_14__sbox_inst_com_z_inst_n456)
         );
  XNOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U8 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n495), .B(round_inst_sin_y[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n439) );
  NAND3_X1 round_inst_S_14__sbox_inst_com_z_inst_U7 ( .A1(round_inst_sin_w[58]), .A2(round_inst_S_14__sbox_inst_com_z_inst_n495), .A3(
        round_inst_S_14__sbox_inst_com_z_inst_n475), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U6 ( .A(round_inst_n69), .B(
        round_inst_sin_y[57]), .Z(round_inst_S_14__sbox_inst_com_z_inst_n475)
         );
  INV_X1 round_inst_S_14__sbox_inst_com_z_inst_U5 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n495) );
  INV_X1 round_inst_S_14__sbox_inst_com_z_inst_U4 ( .A(round_inst_sin_x[59]), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n397) );
  INV_X1 round_inst_S_14__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_14__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_14__sbox_inst_com_z_inst_n497) );
  INV_X1 round_inst_S_14__sbox_inst_com_z_inst_U2 ( .A(round_inst_sin_w[56]), 
        .ZN(round_inst_S_14__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_14__sbox_inst_com_z_inst_U1 ( .A(round_inst_n58), .B(
        round_inst_n68), .Z(round_inst_S_14__sbox_inst_com_z_inst_n417) );
  INV_X1 round_inst_S_15__sbox_inst_U6 ( .A(bout[2]), .ZN(
        round_inst_S_15__sbox_inst_n6) );
  INV_X1 round_inst_S_15__sbox_inst_U5 ( .A(dout[1]), .ZN(
        round_inst_S_15__sbox_inst_n2) );
  INV_X1 round_inst_S_15__sbox_inst_U4 ( .A(dout[3]), .ZN(
        round_inst_S_15__sbox_inst_n4) );
  INV_X2 round_inst_S_15__sbox_inst_U3 ( .A(round_inst_S_15__sbox_inst_n2), 
        .ZN(round_inst_S_15__sbox_inst_n1) );
  INV_X2 round_inst_S_15__sbox_inst_U2 ( .A(round_inst_S_15__sbox_inst_n4), 
        .ZN(round_inst_S_15__sbox_inst_n3) );
  INV_X2 round_inst_S_15__sbox_inst_U1 ( .A(round_inst_S_15__sbox_inst_n6), 
        .ZN(round_inst_S_15__sbox_inst_n5) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U141 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n531), .ZN(round_inst_sout_w[63]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U140 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n530), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n529), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n531) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U139 ( .A1(dout[0]), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n528), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n529) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U138 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n527), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n526), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n530) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U137 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n525), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n524), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n526) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U136 ( .A1(dout[2]), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n523), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n524) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U135 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n521), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n523) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U134 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n520), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n519), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n525) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U133 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n518), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n517), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n519) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U132 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n517) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U131 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n516), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n515), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n518) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U130 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n514), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n513), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n515) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U129 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n512), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n511), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n513) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_w_inst_U128 ( .A1(
        round_inst_S_15__sbox_inst_n5), .A2(bout[0]), .A3(
        round_inst_S_15__sbox_inst_com_w_inst_n510), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n511) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U127 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n509), .A2(cout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n512) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U126 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n508), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n507), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n514) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U125 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n505), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n508) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_w_inst_U124 ( .A1(
        round_inst_S_15__sbox_inst_n3), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n504), .A3(bout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n516) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U123 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n503), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n502), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n527) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U122 ( .A(
        round_inst_sin_y[59]), .B(round_inst_S_15__sbox_inst_com_w_inst_n501), 
        .ZN(round_inst_S_15__sbox_inst_com_w_inst_n502) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U121 ( .A(bout[1]), .B(
        round_inst_sin_z[59]), .Z(round_inst_S_15__sbox_inst_com_w_inst_n501)
         );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U120 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n500), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n499), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n503) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U119 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n506), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n500) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U118 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n497), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n496), .ZN(round_inst_sout_w[61]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U117 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n495), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n494), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n496) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U116 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n493), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n492), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n494) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U115 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n491), .B(round_inst_sin_z[57]), 
        .ZN(round_inst_S_15__sbox_inst_com_w_inst_n492) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U114 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n490), .B(round_inst_sin_y[57]), 
        .ZN(round_inst_S_15__sbox_inst_com_w_inst_n491) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U113 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n489), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n488), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n495) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U112 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n487), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n486), .ZN(round_inst_sout_w[60]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U111 ( .A(
        round_inst_S_15__sbox_inst_n5), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n485), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n487) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U110 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n484), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n483), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n485) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U109 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n532), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n483) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U108 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n528), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n497), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n532) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U107 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n481), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n480), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n497) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U106 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n479), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n478), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n480) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U105 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n477), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n478) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U104 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n488), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n475), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n479) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U103 ( .A(
        round_inst_S_15__sbox_inst_n5), .B(dout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n488) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U102 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n474), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n473), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n481) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U101 ( .A1(
        round_inst_S_15__sbox_inst_n1), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n490), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n473) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U100 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n507), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n499), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n490) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U99 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n504), .A2(bout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n499) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U98 ( .A1(
        round_inst_S_15__sbox_inst_n5), .A2(cout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n507) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U97 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n472), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n471), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n474) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U96 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n470), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n469), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n471) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U95 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n468), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n467), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n469) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U94 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n466), .A2(dout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n467) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U93 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n465), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n468) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U92 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n463), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n462), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n470) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U91 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n461), .A2(bout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n462) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U90 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n460), .B(dout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n461) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U89 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n459), .A2(
        round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n460) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U88 ( .A1(dout[0]), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n458), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n463) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U87 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n456), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n458) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U86 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n455), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n454), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n472) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_w_inst_U85 ( .A1(cout[1]), .A2(
        cout[0]), .A3(round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n454) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_w_inst_U84 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n504), .A2(bout[1]), .A3(cout[0]), .ZN(round_inst_S_15__sbox_inst_com_w_inst_n455) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U83 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n453), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n452), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n528) );
  OR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U82 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n486), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n476), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n453) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U81 ( .A(
        round_inst_S_15__sbox_inst_n5), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n504), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n476) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U80 ( .A(round_inst_n59), .B(
        round_inst_sin_z[56]), .Z(round_inst_S_15__sbox_inst_com_w_inst_n484)
         );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U79 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n451), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n493), .ZN(round_inst_xin_w[63])
         );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U78 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n450), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n449), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n493) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U77 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n448), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n447), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n449) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U76 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n446), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n445), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n447) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U75 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n444), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n443), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n445) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U74 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n442), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n441), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n443) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U73 ( .A1(
        round_inst_S_15__sbox_inst_n3), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n440), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n441) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U72 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n457), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n456), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n440) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U71 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n504), .A2(bout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n456) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U70 ( .A1(
        round_inst_S_15__sbox_inst_n5), .A2(cout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n457) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U69 ( .A1(
        round_inst_S_15__sbox_inst_n1), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n509), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n442) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_w_inst_U68 ( .A1(
        round_inst_S_15__sbox_inst_n5), .A2(round_inst_S_15__sbox_inst_n1), 
        .A3(round_inst_S_15__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n444) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U67 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n439), .A2(bout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n446) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U66 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n438), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n437), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n439) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U65 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n509), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n452), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n437) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U64 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n505), .A2(
        round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n452) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U63 ( .A(
        round_inst_S_15__sbox_inst_n3), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n498), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n505) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U62 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n436), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n509) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U61 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n435), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n438) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U60 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n435) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U59 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n433), .A2(
        round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n448) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U58 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n432), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n431), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n433) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U57 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n430), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n431) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U56 ( .A(cout[1]), .B(
        round_inst_S_15__sbox_inst_n1), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n430) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U55 ( .A1(
        round_inst_S_15__sbox_inst_n3), .A2(round_inst_S_15__sbox_inst_n1), 
        .ZN(round_inst_S_15__sbox_inst_com_w_inst_n432) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U54 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n429), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n428), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n450) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U53 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n427), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n426), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n428) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_w_inst_U52 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n425), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n506), .A3(
        round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n426) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U51 ( .A(cout[1]), .B(bout[1]), 
        .Z(round_inst_S_15__sbox_inst_com_w_inst_n425) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_w_inst_U50 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n506), .A2(cout[1]), .A3(
        round_inst_S_15__sbox_inst_com_w_inst_n465), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n429) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U49 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n504), .B(dout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n465) );
  INV_X1 round_inst_S_15__sbox_inst_com_w_inst_U48 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n436), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n504) );
  INV_X1 round_inst_S_15__sbox_inst_com_w_inst_U47 ( .A(cout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n436) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U46 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n424), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n520), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n451) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U45 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n423), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n422), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n520) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U44 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n421), .A2(
        round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n422) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U43 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n420), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n421) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U42 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n419), .A2(bout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n420) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U41 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n489), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n418), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n419) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U40 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n417), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n416), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n423) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U39 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n521), .A2(
        round_inst_S_15__sbox_inst_n1), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n416) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U38 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n434), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n489), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n521) );
  INV_X1 round_inst_S_15__sbox_inst_com_w_inst_U37 ( .A(bout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n489) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U36 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n415), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n414), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n417) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U35 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n413), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n412), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n414) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U34 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n427), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n459), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n412) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U33 ( .A(bout[0]), .B(dout[0]), .ZN(round_inst_S_15__sbox_inst_com_w_inst_n459) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U32 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n498), .A2(bout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n427) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U31 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n411), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n410), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n413) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U30 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n409), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n408), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n410) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U29 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n407), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n498), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n408) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U28 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n466), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n409) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U27 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n406), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n466) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U26 ( .A1(bout[1]), .A2(
        dout[0]), .ZN(round_inst_S_15__sbox_inst_com_w_inst_n406) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U25 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n405), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n522), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n411) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U24 ( .A(bout[1]), .B(
        round_inst_S_15__sbox_inst_n1), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n405) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U23 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n404), .A2(
        round_inst_S_15__sbox_inst_com_w_inst_n506), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n415) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U22 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n403), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n464), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n404) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U21 ( .A1(bout[0]), .A2(
        bout[1]), .ZN(round_inst_S_15__sbox_inst_com_w_inst_n464) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U20 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n418), .A2(cout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n403) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U19 ( .A(cout[0]), .B(dout[0]), 
        .Z(round_inst_S_15__sbox_inst_com_w_inst_n418) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U18 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n402), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n401), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n424) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U17 ( .A(bout[0]), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n482), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n401) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U16 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n400), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n399), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n482) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U15 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n398), .A2(bout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n399) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U14 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n397), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n396), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n398) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U13 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n498), .B(bout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n396) );
  INV_X1 round_inst_S_15__sbox_inst_com_w_inst_U12 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n434), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n498) );
  INV_X1 round_inst_S_15__sbox_inst_com_w_inst_U11 ( .A(cout[3]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n434) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U10 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n510), .B(
        round_inst_S_15__sbox_inst_n1), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n397) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U9 ( .A(
        round_inst_S_15__sbox_inst_n3), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n506), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n510) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U8 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n522), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n407), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n400) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U7 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n477), .B(
        round_inst_S_15__sbox_inst_com_w_inst_n475), .Z(
        round_inst_S_15__sbox_inst_com_w_inst_n407) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U6 ( .A1(bout[1]), .A2(
        cout[0]), .ZN(round_inst_S_15__sbox_inst_com_w_inst_n475) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U5 ( .A1(bout[0]), .A2(
        cout[1]), .ZN(round_inst_S_15__sbox_inst_com_w_inst_n477) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_w_inst_U4 ( .A1(
        round_inst_S_15__sbox_inst_com_w_inst_n506), .A2(cout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n522) );
  INV_X1 round_inst_S_15__sbox_inst_com_w_inst_U3 ( .A(
        round_inst_S_15__sbox_inst_com_w_inst_n486), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n506) );
  INV_X1 round_inst_S_15__sbox_inst_com_w_inst_U2 ( .A(bout[3]), .ZN(
        round_inst_S_15__sbox_inst_com_w_inst_n486) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_w_inst_U1 ( .A(round_inst_n60), .B(
        round_inst_sin_z[58]), .Z(round_inst_S_15__sbox_inst_com_w_inst_n402)
         );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U135 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n510), .ZN(round_inst_sout_x[60]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U134 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n509), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n508), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n510) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U133 ( .A(cout[2]), .B(
        cout[3]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n508) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U132 ( .A(round_inst_sin_z[56]), .B(round_inst_S_15__sbox_inst_com_x_inst_n507), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n509) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U131 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n511), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n506), .Z(
        round_inst_srout2_x[62]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U130 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n505), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n504), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n506) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U129 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n503), .A2(dout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n504) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U128 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n502), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n501), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n505) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U127 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n500), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n499), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n501) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U126 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n498), .A2(
        round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n499) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U125 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n496), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n498) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U124 ( .A1(cout[2]), .A2(
        round_inst_sin_w[60]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n496)
         );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U123 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n494), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n500) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U122 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n493), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n492), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n494) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U121 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n491), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n492) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U120 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n489), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n488), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n493) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U119 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n487), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n486), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n488) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U118 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n485), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n484), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n486) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U117 ( .A1(cout[3]), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n490), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n484) );
  OR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U116 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n483), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n485) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U115 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n481), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n487) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_x_inst_U114 ( .A1(dout[2]), .A2(
        round_inst_sin_w[60]), .A3(cout[3]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n489) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U113 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n479), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n478), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n502) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U112 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n476), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n478) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U111 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n475), .B(round_inst_sin_z[59]), 
        .ZN(round_inst_S_15__sbox_inst_com_x_inst_n476) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_x_inst_U110 ( .A1(
        round_inst_sin_w[62]), .A2(cout[3]), .A3(dout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n475) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U109 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n474), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n473), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n479) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U108 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n473) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U107 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n471), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n497), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n474) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U106 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n470), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n469), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n511) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U105 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n468), .A2(cout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n469) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U104 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n468) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U103 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n467), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n503), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n470) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U102 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n466), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n503) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U101 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n464), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n480), .ZN(
        round_inst_srout2_x[60]) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U100 ( .A1(cout[0]), .A2(
        dout[2]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n480) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U99 ( .A(round_inst_sin_z[57]), .B(round_inst_S_15__sbox_inst_com_x_inst_n463), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n464) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U98 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n462), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n461), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n463) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U97 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n460), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n467), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n461) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U96 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n459), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n458), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n467) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U95 ( .A1(
        round_inst_S_15__sbox_inst_n1), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n460), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n458) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U94 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n457), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n456), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n459) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U93 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n455), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n454), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n456) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U92 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n453), .A2(round_inst_sin_w[62]), 
        .ZN(round_inst_S_15__sbox_inst_com_x_inst_n454) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U91 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n452), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n451), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n455) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U90 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n450), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n449), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n451) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U89 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n448), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n447), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n449) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U88 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n446), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n447) );
  MUX2_X1 round_inst_S_15__sbox_inst_com_x_inst_U87 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n445), .B(cout[2]), .S(cout[0]), 
        .Z(round_inst_S_15__sbox_inst_com_x_inst_n446) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U86 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n444), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n448) );
  MUX2_X1 round_inst_S_15__sbox_inst_com_x_inst_U85 ( .A(cout[2]), .B(dout[2]), 
        .S(dout[0]), .Z(round_inst_S_15__sbox_inst_com_x_inst_n444) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U84 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n443), .A2(round_inst_sin_w[60]), 
        .ZN(round_inst_S_15__sbox_inst_com_x_inst_n450) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U83 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n442), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n441), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n452) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_x_inst_U82 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[60]), 
        .A3(dout[2]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n441) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_x_inst_U81 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n440), .A2(round_inst_sin_w[61]), 
        .A3(cout[2]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n442) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U80 ( .A(cout[0]), .B(dout[0]), 
        .Z(round_inst_S_15__sbox_inst_com_x_inst_n440) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_x_inst_U79 ( .A1(cout[0]), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n445), .A3(
        round_inst_S_15__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n457) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U78 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n490), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n482), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n460) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U77 ( .A1(cout[0]), .A2(
        cout[2]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n482) );
  AND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U76 ( .A1(cout[2]), .A2(
        dout[0]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n490) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U75 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n497), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n438), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n462) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U74 ( .A1(cout[0]), .A2(
        round_inst_sin_w[62]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n497)
         );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U73 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n495), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n437), .ZN(
        round_inst_srout2_x[63]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U72 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n436), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n435), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n437) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U71 ( .A(cout[0]), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n507), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n435) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U70 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n434), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n433), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n507) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U69 ( .A1(dout[0]), .A2(
        cout[3]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n433) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U68 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n432), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n431), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n434) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U67 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n430), .A2(cout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n431) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U66 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n429), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n428), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n430) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U65 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n428) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U64 ( .A(
        round_inst_S_15__sbox_inst_n1), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n472), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n429) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U63 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n453), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n427), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n432) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U62 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n453) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U61 ( .A(round_inst_sin_z[58]), 
        .B(round_inst_S_15__sbox_inst_com_x_inst_n438), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n436) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U60 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n425), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n424), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n438) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U59 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n423), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n422), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n424) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U58 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n421), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n420), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n422) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U57 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n419), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n418), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n420) );
  NOR3_X1 round_inst_S_15__sbox_inst_com_x_inst_U56 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n471), .A3(
        round_inst_S_15__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n418) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U55 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n416), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n415), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n419) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U54 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n414), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n413), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n415) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U53 ( .A1(cout[2]), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n413) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U52 ( .A(cout[3]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n414) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U51 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n443), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n416) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U50 ( .A1(
        round_inst_S_15__sbox_inst_n1), .A2(cout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n443) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_x_inst_U49 ( .A1(cout[2]), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_15__sbox_inst_com_x_inst_n412), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n421) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U48 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n411), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n465), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n423) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U47 ( .A1(cout[2]), .A2(
        round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n465) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U46 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n411) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U45 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n410), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n409), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n425) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U44 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n408), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n407), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n409) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U43 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n406), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n405), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n407) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U42 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n466), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n439), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n405) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U41 ( .A(round_inst_sin_w[61]), 
        .B(round_inst_S_15__sbox_inst_n1), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n439) );
  AND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U40 ( .A1(dout[2]), .A2(
        cout[3]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n466) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U39 ( .A1(
        round_inst_S_15__sbox_inst_n3), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n406) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_x_inst_U38 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n445), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .A3(
        round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n408) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U37 ( .A(dout[2]), .B(
        round_inst_sin_w[62]), .Z(round_inst_S_15__sbox_inst_com_x_inst_n445)
         );
  NOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U36 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n404), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n403), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n410) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U35 ( .A(round_inst_sin_w[62]), 
        .B(cout[2]), .Z(round_inst_S_15__sbox_inst_com_x_inst_n403) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U34 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n402), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n401), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n495) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U33 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n400), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n399), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n401) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U32 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n472), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n426), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n399) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U31 ( .A1(dout[0]), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n426) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U30 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n398), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n472) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U29 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n427), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n471), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n400) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U28 ( .A(cout[3]), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n471) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U27 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n397), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n396), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n402) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_x_inst_U26 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n395), .A2(
        round_inst_S_15__sbox_inst_n1), .A3(cout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n396) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U25 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n481), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n395) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U24 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n398), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n481) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U23 ( .A(cout[3]), .B(
        round_inst_S_15__sbox_inst_n3), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n398) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U22 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n394), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n393), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n397) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U21 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n392), .A2(round_inst_sin_w[60]), 
        .ZN(round_inst_S_15__sbox_inst_com_x_inst_n393) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U20 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n404), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n392) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U19 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n391), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n390), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n394) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U18 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n389), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n388), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n390) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_x_inst_U17 ( .A1(dout[0]), .A2(
        cout[3]), .A3(round_inst_sin_w[61]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n388) );
  MUX2_X1 round_inst_S_15__sbox_inst_com_x_inst_U16 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n412), .B(cout[3]), .S(
        round_inst_S_15__sbox_inst_com_x_inst_n387), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n389) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U15 ( .A1(cout[0]), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n387) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U14 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n491), .B(
        round_inst_S_15__sbox_inst_n3), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n412) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U13 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n386), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n385), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n391) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U12 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n384), .A2(dout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n385) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U11 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n404), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n383), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n384) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U10 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .A2(
        round_inst_S_15__sbox_inst_com_x_inst_n491), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n383) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U9 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n483), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n491) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U8 ( .A(round_inst_sin_w[63]), 
        .ZN(round_inst_S_15__sbox_inst_com_x_inst_n483) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U7 ( .A1(
        round_inst_S_15__sbox_inst_n1), .A2(cout[3]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n404) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U6 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n382), .A2(
        round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n386) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_x_inst_U5 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n381), .B(
        round_inst_S_15__sbox_inst_com_x_inst_n427), .Z(
        round_inst_S_15__sbox_inst_com_x_inst_n382) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U4 ( .A1(cout[0]), .A2(
        round_inst_sin_w[61]), .ZN(round_inst_S_15__sbox_inst_com_x_inst_n427)
         );
  NAND2_X1 round_inst_S_15__sbox_inst_com_x_inst_U3 ( .A1(
        round_inst_S_15__sbox_inst_com_x_inst_n477), .A2(round_inst_sin_w[60]), 
        .ZN(round_inst_S_15__sbox_inst_com_x_inst_n381) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U2 ( .A(
        round_inst_S_15__sbox_inst_com_x_inst_n417), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n477) );
  INV_X1 round_inst_S_15__sbox_inst_com_x_inst_U1 ( .A(cout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_x_inst_n417) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U137 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n517), .Z(round_inst_sout_y[60])
         );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U136 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n516), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n515), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n517) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U135 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n515) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U134 ( .A(round_inst_sin_x[56]), .B(round_inst_S_15__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n516) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U133 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n512), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n511), .ZN(
        round_inst_srout2_y[62]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U132 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n518), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n511) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U131 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n508), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n518) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U130 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n507), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n506), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n508) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U129 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n506) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U128 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n507) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U127 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n502), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n501), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n512) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U126 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n500), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n499), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n501) );
  NOR3_X1 round_inst_S_15__sbox_inst_com_y_inst_U125 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n498), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n497), .A3(
        round_inst_S_15__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n499) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U124 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n495), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n494), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n500) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U123 ( .A1(bout[3]), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n494) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U122 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n492), .A2(
        round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n495) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U121 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n491), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n490), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n492) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U120 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n489), .A2(round_inst_sin_w[60]), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n491) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U119 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n488), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n487), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n502) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U118 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n486), .A2(
        round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n487) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U117 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n485), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n484), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n486) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U116 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n503), .A2(round_inst_sin_w[60]), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n484) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U115 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n485) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U114 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n482), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n481), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n488) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U113 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n480), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n479), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n481) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U112 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n478), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n504), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n479) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U111 ( .A(
        round_inst_S_15__sbox_inst_n1), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n477), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n480) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U110 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n476), .B(round_inst_sin_x[59]), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n477) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_y_inst_U109 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_15__sbox_inst_n3), .A3(bout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n476) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U108 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n475), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n474), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n482) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_y_inst_U107 ( .A1(
        round_inst_sin_w[60]), .A2(round_inst_sin_w[63]), .A3(
        round_inst_S_15__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n474) );
  OR3_X1 round_inst_S_15__sbox_inst_com_y_inst_U106 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n473), .A3(
        round_inst_S_15__sbox_inst_com_y_inst_n472), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n475) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U105 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n471), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n470), .ZN(
        round_inst_srout2_y[60]) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U104 ( .A1(
        round_inst_S_15__sbox_inst_n5), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n470) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U103 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n469), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n468), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n471) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U102 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n467), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n466), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n468) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U101 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n509), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n465), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n466) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U100 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n464), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n463), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n509) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U99 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n462), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n461), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n463) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U98 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n460), .A2(
        round_inst_S_15__sbox_inst_n1), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n461) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U97 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n490), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n493), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n460) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U96 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n469), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n493) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U95 ( .A1(bout[0]), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n490) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_y_inst_U94 ( .A1(
        round_inst_sin_w[60]), .A2(bout[1]), .A3(
        round_inst_S_15__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n462) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U93 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n459), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n458), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n464) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U92 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n457), .A2(
        round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n458) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U91 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n455), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n457) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U90 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n454), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n453), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n459) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U89 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n452), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n451), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n453) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U88 ( .A1(
        round_inst_S_15__sbox_inst_n1), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n450), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n451) );
  MUX2_X1 round_inst_S_15__sbox_inst_com_y_inst_U87 ( .A(
        round_inst_S_15__sbox_inst_n5), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n503), .S(
        round_inst_S_15__sbox_inst_com_y_inst_n483), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n450) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U86 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n449), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n448), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n452) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U85 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n447), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n446), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n448) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U84 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n445), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n446) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U83 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n497), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n447) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U82 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n443), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n449) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U81 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n441), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n440), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n454) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U80 ( .A(
        round_inst_S_15__sbox_inst_n1), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n440) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U79 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n478), .B(round_inst_n69), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n467) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U78 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n503), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n478) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U77 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n514), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n469) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U76 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n465), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n438), .Z(
        round_inst_srout2_y[63]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U75 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n437), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n436), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n438) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U74 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n483), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n510), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n436) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U73 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n435), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n434), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n510) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U72 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n433), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n432), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n434) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U71 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n445), .A2(round_inst_sin_w[63]), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n432) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U70 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n455), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n431), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n445) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U69 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n483), .A2(bout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n431) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U68 ( .A1(
        round_inst_S_15__sbox_inst_n1), .A2(round_inst_sin_w[60]), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n455) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_y_inst_U67 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n443), .A2(bout[3]), .A3(
        round_inst_S_15__sbox_inst_n1), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n433) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U66 ( .A(round_inst_sin_w[60]), 
        .B(bout[0]), .Z(round_inst_S_15__sbox_inst_com_y_inst_n443) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U65 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n430), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n429), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n435) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U64 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n428), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n427), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n429) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U63 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n426), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n456), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n427) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U62 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n425), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n428) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U61 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n424), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n423), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n430) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U60 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n422), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n421), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n423) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U59 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n420), .A2(round_inst_sin_w[63]), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n421) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U58 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n456), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n444), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n420) );
  AND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U57 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n483), .A2(round_inst_sin_w[61]), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n456) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U56 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n473), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n419), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n422) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U55 ( .A(bout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n473) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U54 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n418), .A2(
        round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n424) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U53 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n425), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n417), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n418) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U52 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n444), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n416), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n417) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U51 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n415), .A2(round_inst_sin_w[60]), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n416) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U50 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n414), .B(bout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n415) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U49 ( .A(round_inst_sin_w[61]), .B(round_inst_S_15__sbox_inst_n1), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n414) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U48 ( .A1(
        round_inst_S_15__sbox_inst_n1), .A2(bout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n444) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U47 ( .A1(
        round_inst_S_15__sbox_inst_n1), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n483), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n425) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U46 ( .A(round_inst_sin_x[58]), 
        .B(round_inst_S_15__sbox_inst_com_y_inst_n513), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n437) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U45 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n413), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n412), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n513) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U44 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n496), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n411), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n412) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U43 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n410), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n409), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n411) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U42 ( .A(round_inst_sin_w[61]), 
        .B(bout[3]), .Z(round_inst_S_15__sbox_inst_com_y_inst_n409) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U41 ( .A(bout[1]), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n498), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n410) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U40 ( .A(round_inst_sin_w[63]), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n498) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U39 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n408), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n439), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n413) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U38 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n483), .B(round_inst_sin_w[60]), 
        .Z(round_inst_S_15__sbox_inst_com_y_inst_n439) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U37 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n496), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n483) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U36 ( .A(dout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n496) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U35 ( .A(
        round_inst_S_15__sbox_inst_n1), .B(round_inst_S_15__sbox_inst_n3), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n408) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U34 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n407), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n406), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n465) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U33 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n405), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n404), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n406) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U32 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n403), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n402), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n404) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U31 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n401), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n400), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n402) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U30 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n419), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n497), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n400) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U29 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n489), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n497) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U28 ( .A(
        round_inst_S_15__sbox_inst_n5), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n489) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U27 ( .A1(
        round_inst_sin_w[61]), .A2(round_inst_S_15__sbox_inst_n3), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n419) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U26 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n472), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n442), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n401) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U25 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n514), .A2(round_inst_sin_w[61]), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n442) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_y_inst_U24 ( .A1(
        round_inst_S_15__sbox_inst_n1), .A2(round_inst_sin_w[63]), .A3(
        round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n403) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U23 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n399), .A2(
        round_inst_S_15__sbox_inst_n1), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n405) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U22 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n398), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n397), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n399) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U21 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n396), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n397) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U20 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n504), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n394), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n398) );
  OR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U19 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n505), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n395), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n394) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U18 ( .A(
        round_inst_S_15__sbox_inst_n3), .B(round_inst_sin_w[63]), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n395) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U17 ( .A(
        round_inst_S_15__sbox_inst_n3), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n472), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n504) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U16 ( .A(round_inst_sin_w[63]), .B(bout[3]), .ZN(round_inst_S_15__sbox_inst_com_y_inst_n472) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U15 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n393), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n392), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n407) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U14 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n391), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n390), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n392) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_y_inst_U13 ( .A1(bout[1]), .A2(
        round_inst_sin_w[63]), .A3(round_inst_S_15__sbox_inst_com_y_inst_n514), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n390) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_y_inst_U12 ( .A1(
        round_inst_S_15__sbox_inst_n3), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n389), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n391) );
  MUX2_X1 round_inst_S_15__sbox_inst_com_y_inst_U11 ( .A(round_inst_sin_w[61]), 
        .B(bout[1]), .S(round_inst_S_15__sbox_inst_com_y_inst_n503), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n389) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U10 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n388), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n387), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n393) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_y_inst_U9 ( .A1(bout[1]), .A2(
        round_inst_S_15__sbox_inst_com_y_inst_n426), .A3(
        round_inst_S_15__sbox_inst_com_y_inst_n514), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n387) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U8 ( .A(
        round_inst_S_15__sbox_inst_n3), .B(bout[3]), .Z(
        round_inst_S_15__sbox_inst_com_y_inst_n426) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_y_inst_U7 ( .A1(
        round_inst_S_15__sbox_inst_com_y_inst_n386), .A2(
        round_inst_S_15__sbox_inst_n1), .A3(bout[3]), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n388) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U6 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n441), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n386) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_y_inst_U5 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n514), .B(
        round_inst_S_15__sbox_inst_com_y_inst_n503), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n441) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U4 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n396), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n503) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U3 ( .A(round_inst_sin_w[62]), 
        .ZN(round_inst_S_15__sbox_inst_com_y_inst_n396) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U2 ( .A(
        round_inst_S_15__sbox_inst_com_y_inst_n505), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n514) );
  INV_X1 round_inst_S_15__sbox_inst_com_y_inst_U1 ( .A(dout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_y_inst_n505) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U132 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n517), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n516), .ZN(round_inst_sout_z[60]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U131 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n515), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n514), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n516) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U130 ( .A(
        round_inst_sin_w[62]), .B(round_inst_sin_w[63]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n514) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U129 ( .A(round_inst_sin_x[56]), .B(round_inst_n59), .Z(round_inst_S_15__sbox_inst_com_z_inst_n515) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U128 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n512), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n517) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U127 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n513), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n511), .ZN(
        round_inst_srout2_z[62]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U126 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n510), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n509), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n511) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U125 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n508), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n507), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n509) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U124 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n506), .A2(cout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n507) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U123 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n505), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n504), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n508) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U122 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n503), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n502), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n504) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U121 ( .A(
        round_inst_sin_w[61]), .B(round_inst_sin_x[59]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n502) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U120 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n501), .B(round_inst_sin_y[59]), 
        .Z(round_inst_S_15__sbox_inst_com_z_inst_n503) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U119 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n500), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n499), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n501) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U118 ( .A1(cout[2]), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n498), .A3(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n499) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U117 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n496), .A2(bout[0]), .A3(
        round_inst_sin_w[63]), .ZN(round_inst_S_15__sbox_inst_com_z_inst_n500)
         );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U116 ( .A(
        round_inst_S_15__sbox_inst_n5), .B(cout[2]), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n496) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U115 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_15__sbox_inst_n5), .A3(bout[3]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n505) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U114 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n495), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n494), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n510) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U113 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n493), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n492), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n494) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U112 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n491), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n490), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n492) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U111 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n489), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n488), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n490) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U110 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n487), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n491) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U109 ( .A1(
        round_inst_sin_w[62]), .A2(bout[3]), .A3(cout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n493) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U108 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n485), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n486), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n513) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U107 ( .A1(
        round_inst_sin_w[62]), .A2(round_inst_S_15__sbox_inst_com_z_inst_n498), 
        .ZN(round_inst_S_15__sbox_inst_com_z_inst_n486) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U106 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n484), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n506), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n485) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U105 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n483), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n482), .Z(
        round_inst_srout2_z[60]) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U104 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n481), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n480), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n482) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U103 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n479), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n484), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n480) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U102 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n478), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n477), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n484) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U101 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n476), .A2(bout[0]), .A3(
        round_inst_sin_w[62]), .ZN(round_inst_S_15__sbox_inst_com_z_inst_n477)
         );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U100 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n475), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n474), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n478) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U99 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n473), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .A3(cout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n474) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U98 ( .A(round_inst_sin_w[61]), 
        .B(cout[1]), .Z(round_inst_S_15__sbox_inst_com_z_inst_n473) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U97 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n472), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n471), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n475) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U96 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n470), .A2(
        round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n471) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U95 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n469), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n468), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n472) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U94 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n467), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n466), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n468) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U93 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n465), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n464), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n466) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U92 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n463), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n462), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n464) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U91 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n461), .A2(cout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n462) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U90 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n460), .A2(
        round_inst_S_15__sbox_inst_n5), .A3(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n463) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U89 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n459), .A2(cout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n465) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U88 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n458), .A2(round_inst_sin_w[62]), 
        .ZN(round_inst_S_15__sbox_inst_com_z_inst_n467) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U87 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n457), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n469) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U86 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n455), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n454), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n457) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U85 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n453), .A2(cout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n454) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U84 ( .A(round_inst_sin_w[61]), .B(round_inst_S_15__sbox_inst_com_z_inst_n452), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n453) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U83 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n451), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n450), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n455) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U82 ( .A1(
        round_inst_sin_w[62]), .A2(bout[0]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n479) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U81 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n449), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n448), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n481) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U80 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n488), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n447), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n448) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U79 ( .A(round_inst_sin_y[57]), 
        .B(round_inst_n69), .Z(round_inst_S_15__sbox_inst_com_z_inst_n447) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U78 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n488) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U77 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n446), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n483) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U76 ( .A(round_inst_sin_w[62]), .B(cout[2]), .ZN(round_inst_S_15__sbox_inst_com_z_inst_n446) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U75 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n444), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n443), .ZN(
        round_inst_srout2_z[63]) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U74 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n495), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n512), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n443) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U73 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n442), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n441), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n512) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U72 ( .A1(bout[0]), .A2(
        round_inst_sin_w[63]), .ZN(round_inst_S_15__sbox_inst_com_z_inst_n441)
         );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U71 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n458), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n440), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n442) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U70 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n498), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n440) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U69 ( .A(round_inst_sin_w[63]), .B(round_inst_S_15__sbox_inst_com_z_inst_n439), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n498) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U68 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n438), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n437), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n495) );
  MUX2_X1 round_inst_S_15__sbox_inst_com_z_inst_U67 ( .A(bout[3]), .B(
        round_inst_sin_w[63]), .S(round_inst_S_15__sbox_inst_com_z_inst_n436), 
        .Z(round_inst_S_15__sbox_inst_com_z_inst_n437) );
  OR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U66 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n487), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n436) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U65 ( .A(bout[0]), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n487) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U64 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n434), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n433), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n438) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U63 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .A2(bout[3]), .A3(
        round_inst_S_15__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n433) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U62 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n432), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n431), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n434) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U61 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n430), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n429), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n431) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U60 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n428), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n427), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n429) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U59 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n426), .A2(round_inst_sin_w[63]), 
        .ZN(round_inst_S_15__sbox_inst_com_z_inst_n427) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U58 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n425), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n424), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n426) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U57 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n423), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n422), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n424) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U56 ( .A1(bout[0]), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n460), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n422) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U55 ( .A1(cout[1]), .A2(
        bout[0]), .ZN(round_inst_S_15__sbox_inst_com_z_inst_n425) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U54 ( .A1(cout[0]), .A2(
        bout[3]), .A3(round_inst_sin_w[61]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n428) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U53 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n458), .A2(cout[3]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n430) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U52 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n421), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n470), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n458) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U51 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n461), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n423), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n470) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U50 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .A2(cout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n423) );
  AND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U49 ( .A1(round_inst_sin_w[61]), .A2(bout[0]), .ZN(round_inst_S_15__sbox_inst_com_z_inst_n461) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U48 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n452), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n420), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n421) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U47 ( .A1(
        round_inst_sin_w[61]), .A2(round_inst_S_15__sbox_inst_com_z_inst_n497), 
        .ZN(round_inst_S_15__sbox_inst_com_z_inst_n420) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U46 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n460), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n452) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U45 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n419), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n418), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n432) );
  INV_X1 round_inst_S_15__sbox_inst_com_z_inst_U44 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n451), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n419) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U43 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .B(cout[0]), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n451) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U42 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n417), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n416), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n444) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U41 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n497), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n449), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n416) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U40 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n415), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n414), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n449) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U39 ( .A1(
        round_inst_sin_w[63]), .A2(round_inst_S_15__sbox_inst_com_z_inst_n413), 
        .ZN(round_inst_S_15__sbox_inst_com_z_inst_n414) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U38 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n450), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n456), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n413) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U37 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n412), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n411), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n415) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U36 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n410), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n409), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n411) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U35 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n506), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n460), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n409) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U34 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n408), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n407), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n410) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U33 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n406), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n405), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n407) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U32 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n404), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n405) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U31 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n403), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n402), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n404) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U30 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n506), .A2(cout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n402) );
  AND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U29 ( .A1(
        round_inst_S_15__sbox_inst_n5), .A2(round_inst_sin_w[63]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n506) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U28 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n401), .A2(cout[2]), .A3(
        round_inst_sin_w[61]), .ZN(round_inst_S_15__sbox_inst_com_z_inst_n403)
         );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U27 ( .A(round_inst_sin_w[63]), 
        .B(bout[3]), .Z(round_inst_S_15__sbox_inst_com_z_inst_n401) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U26 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n400), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n399), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n406) );
  MUX2_X1 round_inst_S_15__sbox_inst_com_z_inst_U25 ( .A(cout[3]), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n398), .S(
        round_inst_S_15__sbox_inst_com_z_inst_n450), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n399) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U24 ( .A1(
        round_inst_sin_w[61]), .A2(round_inst_S_15__sbox_inst_n5), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n450) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U23 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n397), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n398) );
  INV_X1 round_inst_S_15__sbox_inst_com_z_inst_U22 ( .A(bout[3]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n397) );
  NOR3_X1 round_inst_S_15__sbox_inst_com_z_inst_U21 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n396), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n489), .A3(
        round_inst_S_15__sbox_inst_com_z_inst_n395), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n400) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U20 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n394), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n395) );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U19 ( .A(round_inst_sin_w[63]), .B(cout[3]), .ZN(round_inst_S_15__sbox_inst_com_z_inst_n489) );
  AND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U18 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n435), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n459), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n396) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U17 ( .A1(
        round_inst_sin_w[62]), .A2(round_inst_S_15__sbox_inst_com_z_inst_n460), 
        .ZN(round_inst_S_15__sbox_inst_com_z_inst_n459) );
  INV_X1 round_inst_S_15__sbox_inst_com_z_inst_U16 ( .A(round_inst_sin_w[61]), 
        .ZN(round_inst_S_15__sbox_inst_com_z_inst_n435) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U15 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n393), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n392), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n408) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U14 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n391), .A2(cout[2]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n392) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U13 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n418), .B(
        round_inst_S_15__sbox_inst_com_z_inst_n390), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n391) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U12 ( .A1(
        round_inst_sin_w[61]), .A2(cout[3]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n390) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U11 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n460), .A2(round_inst_sin_w[63]), 
        .ZN(round_inst_S_15__sbox_inst_com_z_inst_n418) );
  NOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U10 ( .A1(
        round_inst_S_15__sbox_inst_com_z_inst_n439), .A2(
        round_inst_S_15__sbox_inst_com_z_inst_n456), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n393) );
  NAND2_X1 round_inst_S_15__sbox_inst_com_z_inst_U9 ( .A1(round_inst_sin_w[62]), .A2(round_inst_sin_w[61]), .ZN(round_inst_S_15__sbox_inst_com_z_inst_n456)
         );
  XNOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U8 ( .A(bout[3]), .B(cout[3]), 
        .ZN(round_inst_S_15__sbox_inst_com_z_inst_n439) );
  NAND3_X1 round_inst_S_15__sbox_inst_com_z_inst_U7 ( .A1(round_inst_sin_w[62]), .A2(bout[3]), .A3(round_inst_S_15__sbox_inst_com_z_inst_n476), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n412) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U6 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n460), .B(cout[1]), .Z(
        round_inst_S_15__sbox_inst_com_z_inst_n476) );
  INV_X1 round_inst_S_15__sbox_inst_com_z_inst_U5 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n394), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n460) );
  INV_X1 round_inst_S_15__sbox_inst_com_z_inst_U4 ( .A(bout[1]), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n394) );
  INV_X1 round_inst_S_15__sbox_inst_com_z_inst_U3 ( .A(
        round_inst_S_15__sbox_inst_com_z_inst_n445), .ZN(
        round_inst_S_15__sbox_inst_com_z_inst_n497) );
  INV_X1 round_inst_S_15__sbox_inst_com_z_inst_U2 ( .A(round_inst_sin_w[60]), 
        .ZN(round_inst_S_15__sbox_inst_com_z_inst_n445) );
  XOR2_X1 round_inst_S_15__sbox_inst_com_z_inst_U1 ( .A(round_inst_n60), .B(
        round_inst_sin_x[58]), .Z(round_inst_S_15__sbox_inst_com_z_inst_n417)
         );
  XNOR2_X1 round_inst_A2_0__aw2_U4 ( .A(round_inst_A2_0__aw2_n5), .B(
        round_inst_sout_w[0]), .ZN(round_inst_xin_w[1]) );
  XNOR2_X1 round_inst_A2_0__aw2_U3 ( .A(round_inst_sout_w[1]), .B(
        round_inst_xin_w[3]), .ZN(round_inst_A2_0__aw2_n5) );
  INV_X1 round_inst_A2_0__aw2_U2 ( .A(round_inst_sout_w[3]), .ZN(
        round_inst_xin_w[2]) );
  INV_X1 round_inst_A2_0__aw2_U1 ( .A(round_inst_sout_w[1]), .ZN(
        round_inst_xin_w[0]) );
  XNOR2_X1 round_inst_A2_0__ax2_U2 ( .A(round_inst_A2_0__ax2_n3), .B(
        round_inst_sout_x[0]), .ZN(round_inst_srout2_x[17]) );
  XNOR2_X1 round_inst_A2_0__ax2_U1 ( .A(round_inst_srout2_x[16]), .B(
        round_inst_srout2_x[19]), .ZN(round_inst_A2_0__ax2_n3) );
  XNOR2_X1 round_inst_A2_0__ay2_U2 ( .A(round_inst_A2_0__ay2_n3), .B(
        round_inst_sout_y[0]), .ZN(round_inst_srout2_y[17]) );
  XNOR2_X1 round_inst_A2_0__ay2_U1 ( .A(round_inst_srout2_y[16]), .B(
        round_inst_srout2_y[19]), .ZN(round_inst_A2_0__ay2_n3) );
  XNOR2_X1 round_inst_A2_0__az2_U2 ( .A(round_inst_A2_0__az2_n3), .B(
        round_inst_sout_z[0]), .ZN(round_inst_srout2_z[17]) );
  XNOR2_X1 round_inst_A2_0__az2_U1 ( .A(round_inst_srout2_z[16]), .B(
        round_inst_srout2_z[19]), .ZN(round_inst_A2_0__az2_n3) );
  XNOR2_X1 round_inst_A2_1__aw2_U4 ( .A(round_inst_A2_1__aw2_n5), .B(
        round_inst_sout_w[4]), .ZN(round_inst_xin_w[5]) );
  XNOR2_X1 round_inst_A2_1__aw2_U3 ( .A(round_inst_sout_w[5]), .B(
        round_inst_xin_w[7]), .ZN(round_inst_A2_1__aw2_n5) );
  INV_X1 round_inst_A2_1__aw2_U2 ( .A(round_inst_sout_w[7]), .ZN(
        round_inst_xin_w[6]) );
  INV_X1 round_inst_A2_1__aw2_U1 ( .A(round_inst_sout_w[5]), .ZN(
        round_inst_xin_w[4]) );
  XNOR2_X1 round_inst_A2_1__ax2_U2 ( .A(round_inst_A2_1__ax2_n3), .B(
        round_inst_sout_x[4]), .ZN(round_inst_srout2_x[37]) );
  XNOR2_X1 round_inst_A2_1__ax2_U1 ( .A(round_inst_srout2_x[36]), .B(
        round_inst_srout2_x[39]), .ZN(round_inst_A2_1__ax2_n3) );
  XNOR2_X1 round_inst_A2_1__ay2_U2 ( .A(round_inst_A2_1__ay2_n3), .B(
        round_inst_sout_y[4]), .ZN(round_inst_srout2_y[37]) );
  XNOR2_X1 round_inst_A2_1__ay2_U1 ( .A(round_inst_srout2_y[36]), .B(
        round_inst_srout2_y[39]), .ZN(round_inst_A2_1__ay2_n3) );
  XNOR2_X1 round_inst_A2_1__az2_U2 ( .A(round_inst_A2_1__az2_n3), .B(
        round_inst_sout_z[4]), .ZN(round_inst_srout2_z[37]) );
  XNOR2_X1 round_inst_A2_1__az2_U1 ( .A(round_inst_srout2_z[36]), .B(
        round_inst_srout2_z[39]), .ZN(round_inst_A2_1__az2_n3) );
  XNOR2_X1 round_inst_A2_2__aw2_U4 ( .A(round_inst_A2_2__aw2_n5), .B(
        round_inst_sout_w[8]), .ZN(round_inst_xin_w[9]) );
  XNOR2_X1 round_inst_A2_2__aw2_U3 ( .A(round_inst_sout_w[9]), .B(
        round_inst_xin_w[11]), .ZN(round_inst_A2_2__aw2_n5) );
  INV_X1 round_inst_A2_2__aw2_U2 ( .A(round_inst_sout_w[11]), .ZN(
        round_inst_xin_w[10]) );
  INV_X1 round_inst_A2_2__aw2_U1 ( .A(round_inst_sout_w[9]), .ZN(
        round_inst_xin_w[8]) );
  XNOR2_X1 round_inst_A2_2__ax2_U2 ( .A(round_inst_A2_2__ax2_n3), .B(
        round_inst_sout_x[8]), .ZN(round_inst_srout2_x[57]) );
  XNOR2_X1 round_inst_A2_2__ax2_U1 ( .A(round_inst_srout2_x[56]), .B(
        round_inst_srout2_x[59]), .ZN(round_inst_A2_2__ax2_n3) );
  XNOR2_X1 round_inst_A2_2__ay2_U2 ( .A(round_inst_A2_2__ay2_n3), .B(
        round_inst_sout_y[8]), .ZN(round_inst_srout2_y[57]) );
  XNOR2_X1 round_inst_A2_2__ay2_U1 ( .A(round_inst_srout2_y[56]), .B(
        round_inst_srout2_y[59]), .ZN(round_inst_A2_2__ay2_n3) );
  XNOR2_X1 round_inst_A2_2__az2_U2 ( .A(round_inst_A2_2__az2_n3), .B(
        round_inst_sout_z[8]), .ZN(round_inst_srout2_z[57]) );
  XNOR2_X1 round_inst_A2_2__az2_U1 ( .A(round_inst_srout2_z[56]), .B(
        round_inst_srout2_z[59]), .ZN(round_inst_A2_2__az2_n3) );
  XNOR2_X1 round_inst_A2_3__aw2_U4 ( .A(round_inst_A2_3__aw2_n5), .B(
        round_inst_sout_w[12]), .ZN(round_inst_xin_w[13]) );
  XNOR2_X1 round_inst_A2_3__aw2_U3 ( .A(round_inst_sout_w[13]), .B(
        round_inst_xin_w[15]), .ZN(round_inst_A2_3__aw2_n5) );
  INV_X1 round_inst_A2_3__aw2_U2 ( .A(round_inst_sout_w[15]), .ZN(
        round_inst_xin_w[14]) );
  INV_X1 round_inst_A2_3__aw2_U1 ( .A(round_inst_sout_w[13]), .ZN(
        round_inst_xin_w[12]) );
  XNOR2_X1 round_inst_A2_3__ax2_U2 ( .A(round_inst_A2_3__ax2_n3), .B(
        round_inst_sout_x[12]), .ZN(round_inst_srout2_x[13]) );
  XNOR2_X1 round_inst_A2_3__ax2_U1 ( .A(round_inst_srout2_x[12]), .B(
        round_inst_srout2_x[15]), .ZN(round_inst_A2_3__ax2_n3) );
  XNOR2_X1 round_inst_A2_3__ay2_U2 ( .A(round_inst_A2_3__ay2_n3), .B(
        round_inst_sout_y[12]), .ZN(round_inst_srout2_y[13]) );
  XNOR2_X1 round_inst_A2_3__ay2_U1 ( .A(round_inst_srout2_y[12]), .B(
        round_inst_srout2_y[15]), .ZN(round_inst_A2_3__ay2_n3) );
  XNOR2_X1 round_inst_A2_3__az2_U2 ( .A(round_inst_A2_3__az2_n3), .B(
        round_inst_sout_z[12]), .ZN(round_inst_srout2_z[13]) );
  XNOR2_X1 round_inst_A2_3__az2_U1 ( .A(round_inst_srout2_z[12]), .B(
        round_inst_srout2_z[15]), .ZN(round_inst_A2_3__az2_n3) );
  XNOR2_X1 round_inst_A2_4__aw2_U4 ( .A(round_inst_A2_4__aw2_n5), .B(
        round_inst_sout_w[16]), .ZN(round_inst_xin_w[17]) );
  XNOR2_X1 round_inst_A2_4__aw2_U3 ( .A(round_inst_sout_w[17]), .B(
        round_inst_xin_w[19]), .ZN(round_inst_A2_4__aw2_n5) );
  INV_X1 round_inst_A2_4__aw2_U2 ( .A(round_inst_sout_w[19]), .ZN(
        round_inst_xin_w[18]) );
  INV_X1 round_inst_A2_4__aw2_U1 ( .A(round_inst_sout_w[17]), .ZN(
        round_inst_xin_w[16]) );
  XNOR2_X1 round_inst_A2_4__ax2_U2 ( .A(round_inst_A2_4__ax2_n3), .B(
        round_inst_sout_x[16]), .ZN(round_inst_srout2_x[33]) );
  XNOR2_X1 round_inst_A2_4__ax2_U1 ( .A(round_inst_srout2_x[32]), .B(
        round_inst_srout2_x[35]), .ZN(round_inst_A2_4__ax2_n3) );
  XNOR2_X1 round_inst_A2_4__ay2_U2 ( .A(round_inst_A2_4__ay2_n3), .B(
        round_inst_sout_y[16]), .ZN(round_inst_srout2_y[33]) );
  XNOR2_X1 round_inst_A2_4__ay2_U1 ( .A(round_inst_srout2_y[32]), .B(
        round_inst_srout2_y[35]), .ZN(round_inst_A2_4__ay2_n3) );
  XNOR2_X1 round_inst_A2_4__az2_U2 ( .A(round_inst_A2_4__az2_n3), .B(
        round_inst_sout_z[16]), .ZN(round_inst_srout2_z[33]) );
  XNOR2_X1 round_inst_A2_4__az2_U1 ( .A(round_inst_srout2_z[32]), .B(
        round_inst_srout2_z[35]), .ZN(round_inst_A2_4__az2_n3) );
  XNOR2_X1 round_inst_A2_5__aw2_U4 ( .A(round_inst_A2_5__aw2_n5), .B(
        round_inst_sout_w[20]), .ZN(round_inst_xin_w[21]) );
  XNOR2_X1 round_inst_A2_5__aw2_U3 ( .A(round_inst_sout_w[21]), .B(
        round_inst_xin_w[23]), .ZN(round_inst_A2_5__aw2_n5) );
  INV_X1 round_inst_A2_5__aw2_U2 ( .A(round_inst_sout_w[23]), .ZN(
        round_inst_xin_w[22]) );
  INV_X1 round_inst_A2_5__aw2_U1 ( .A(round_inst_sout_w[21]), .ZN(
        round_inst_xin_w[20]) );
  XNOR2_X1 round_inst_A2_5__ax2_U2 ( .A(round_inst_A2_5__ax2_n3), .B(
        round_inst_sout_x[20]), .ZN(round_inst_srout2_x[53]) );
  XNOR2_X1 round_inst_A2_5__ax2_U1 ( .A(round_inst_srout2_x[52]), .B(
        round_inst_srout2_x[55]), .ZN(round_inst_A2_5__ax2_n3) );
  XNOR2_X1 round_inst_A2_5__ay2_U2 ( .A(round_inst_A2_5__ay2_n3), .B(
        round_inst_sout_y[20]), .ZN(round_inst_srout2_y[53]) );
  XNOR2_X1 round_inst_A2_5__ay2_U1 ( .A(round_inst_srout2_y[52]), .B(
        round_inst_srout2_y[55]), .ZN(round_inst_A2_5__ay2_n3) );
  XNOR2_X1 round_inst_A2_5__az2_U2 ( .A(round_inst_A2_5__az2_n3), .B(
        round_inst_sout_z[20]), .ZN(round_inst_srout2_z[53]) );
  XNOR2_X1 round_inst_A2_5__az2_U1 ( .A(round_inst_srout2_z[52]), .B(
        round_inst_srout2_z[55]), .ZN(round_inst_A2_5__az2_n3) );
  XNOR2_X1 round_inst_A2_6__aw2_U4 ( .A(round_inst_A2_6__aw2_n5), .B(
        round_inst_sout_w[24]), .ZN(round_inst_xin_w[25]) );
  XNOR2_X1 round_inst_A2_6__aw2_U3 ( .A(round_inst_sout_w[25]), .B(
        round_inst_xin_w[27]), .ZN(round_inst_A2_6__aw2_n5) );
  INV_X1 round_inst_A2_6__aw2_U2 ( .A(round_inst_sout_w[27]), .ZN(
        round_inst_xin_w[26]) );
  INV_X1 round_inst_A2_6__aw2_U1 ( .A(round_inst_sout_w[25]), .ZN(
        round_inst_xin_w[24]) );
  XNOR2_X1 round_inst_A2_6__ax2_U2 ( .A(round_inst_A2_6__ax2_n3), .B(
        round_inst_sout_x[24]), .ZN(round_inst_srout2_x[9]) );
  XNOR2_X1 round_inst_A2_6__ax2_U1 ( .A(round_inst_srout2_x[8]), .B(
        round_inst_srout2_x[11]), .ZN(round_inst_A2_6__ax2_n3) );
  XNOR2_X1 round_inst_A2_6__ay2_U2 ( .A(round_inst_A2_6__ay2_n3), .B(
        round_inst_sout_y[24]), .ZN(round_inst_srout2_y[9]) );
  XNOR2_X1 round_inst_A2_6__ay2_U1 ( .A(round_inst_srout2_y[8]), .B(
        round_inst_srout2_y[11]), .ZN(round_inst_A2_6__ay2_n3) );
  XNOR2_X1 round_inst_A2_6__az2_U2 ( .A(round_inst_A2_6__az2_n3), .B(
        round_inst_sout_z[24]), .ZN(round_inst_srout2_z[9]) );
  XNOR2_X1 round_inst_A2_6__az2_U1 ( .A(round_inst_srout2_z[8]), .B(
        round_inst_srout2_z[11]), .ZN(round_inst_A2_6__az2_n3) );
  XNOR2_X1 round_inst_A2_7__aw2_U4 ( .A(round_inst_A2_7__aw2_n5), .B(
        round_inst_sout_w[28]), .ZN(round_inst_xin_w[29]) );
  XNOR2_X1 round_inst_A2_7__aw2_U3 ( .A(round_inst_sout_w[29]), .B(
        round_inst_xin_w[31]), .ZN(round_inst_A2_7__aw2_n5) );
  INV_X1 round_inst_A2_7__aw2_U2 ( .A(round_inst_sout_w[31]), .ZN(
        round_inst_xin_w[30]) );
  INV_X1 round_inst_A2_7__aw2_U1 ( .A(round_inst_sout_w[29]), .ZN(
        round_inst_xin_w[28]) );
  XNOR2_X1 round_inst_A2_7__ax2_U2 ( .A(round_inst_A2_7__ax2_n3), .B(
        round_inst_sout_x[28]), .ZN(round_inst_srout2_x[29]) );
  XNOR2_X1 round_inst_A2_7__ax2_U1 ( .A(round_inst_srout2_x[28]), .B(
        round_inst_srout2_x[31]), .ZN(round_inst_A2_7__ax2_n3) );
  XNOR2_X1 round_inst_A2_7__ay2_U2 ( .A(round_inst_A2_7__ay2_n3), .B(
        round_inst_sout_y[28]), .ZN(round_inst_srout2_y[29]) );
  XNOR2_X1 round_inst_A2_7__ay2_U1 ( .A(round_inst_srout2_y[28]), .B(
        round_inst_srout2_y[31]), .ZN(round_inst_A2_7__ay2_n3) );
  XNOR2_X1 round_inst_A2_7__az2_U2 ( .A(round_inst_A2_7__az2_n3), .B(
        round_inst_sout_z[28]), .ZN(round_inst_srout2_z[29]) );
  XNOR2_X1 round_inst_A2_7__az2_U1 ( .A(round_inst_srout2_z[28]), .B(
        round_inst_srout2_z[31]), .ZN(round_inst_A2_7__az2_n3) );
  XNOR2_X1 round_inst_A2_8__aw2_U4 ( .A(round_inst_A2_8__aw2_n5), .B(
        round_inst_sout_w[32]), .ZN(round_inst_xin_w[33]) );
  XNOR2_X1 round_inst_A2_8__aw2_U3 ( .A(round_inst_sout_w[33]), .B(
        round_inst_xin_w[35]), .ZN(round_inst_A2_8__aw2_n5) );
  INV_X1 round_inst_A2_8__aw2_U2 ( .A(round_inst_sout_w[35]), .ZN(
        round_inst_xin_w[34]) );
  INV_X1 round_inst_A2_8__aw2_U1 ( .A(round_inst_sout_w[33]), .ZN(
        round_inst_xin_w[32]) );
  XNOR2_X1 round_inst_A2_8__ax2_U2 ( .A(round_inst_A2_8__ax2_n3), .B(
        round_inst_sout_x[32]), .ZN(round_inst_srout2_x[49]) );
  XNOR2_X1 round_inst_A2_8__ax2_U1 ( .A(round_inst_srout2_x[48]), .B(
        round_inst_srout2_x[51]), .ZN(round_inst_A2_8__ax2_n3) );
  XNOR2_X1 round_inst_A2_8__ay2_U2 ( .A(round_inst_A2_8__ay2_n3), .B(
        round_inst_sout_y[32]), .ZN(round_inst_srout2_y[49]) );
  XNOR2_X1 round_inst_A2_8__ay2_U1 ( .A(round_inst_srout2_y[48]), .B(
        round_inst_srout2_y[51]), .ZN(round_inst_A2_8__ay2_n3) );
  XNOR2_X1 round_inst_A2_8__az2_U2 ( .A(round_inst_A2_8__az2_n3), .B(
        round_inst_sout_z[32]), .ZN(round_inst_srout2_z[49]) );
  XNOR2_X1 round_inst_A2_8__az2_U1 ( .A(round_inst_srout2_z[48]), .B(
        round_inst_srout2_z[51]), .ZN(round_inst_A2_8__az2_n3) );
  XNOR2_X1 round_inst_A2_9__aw2_U4 ( .A(round_inst_A2_9__aw2_n5), .B(
        round_inst_sout_w[36]), .ZN(round_inst_xin_w[37]) );
  XNOR2_X1 round_inst_A2_9__aw2_U3 ( .A(round_inst_sout_w[37]), .B(
        round_inst_xin_w[39]), .ZN(round_inst_A2_9__aw2_n5) );
  INV_X1 round_inst_A2_9__aw2_U2 ( .A(round_inst_sout_w[39]), .ZN(
        round_inst_xin_w[38]) );
  INV_X1 round_inst_A2_9__aw2_U1 ( .A(round_inst_sout_w[37]), .ZN(
        round_inst_xin_w[36]) );
  XNOR2_X1 round_inst_A2_9__ax2_U2 ( .A(round_inst_A2_9__ax2_n3), .B(
        round_inst_sout_x[36]), .ZN(round_inst_srout2_x[5]) );
  XNOR2_X1 round_inst_A2_9__ax2_U1 ( .A(round_inst_srout2_x[4]), .B(
        round_inst_srout2_x[7]), .ZN(round_inst_A2_9__ax2_n3) );
  XNOR2_X1 round_inst_A2_9__ay2_U2 ( .A(round_inst_A2_9__ay2_n3), .B(
        round_inst_sout_y[36]), .ZN(round_inst_srout2_y[5]) );
  XNOR2_X1 round_inst_A2_9__ay2_U1 ( .A(round_inst_srout2_y[4]), .B(
        round_inst_srout2_y[7]), .ZN(round_inst_A2_9__ay2_n3) );
  XNOR2_X1 round_inst_A2_9__az2_U2 ( .A(round_inst_A2_9__az2_n3), .B(
        round_inst_sout_z[36]), .ZN(round_inst_srout2_z[5]) );
  XNOR2_X1 round_inst_A2_9__az2_U1 ( .A(round_inst_srout2_z[4]), .B(
        round_inst_srout2_z[7]), .ZN(round_inst_A2_9__az2_n3) );
  XNOR2_X1 round_inst_A2_10__aw2_U4 ( .A(round_inst_A2_10__aw2_n5), .B(
        round_inst_sout_w[40]), .ZN(round_inst_xin_w[41]) );
  XNOR2_X1 round_inst_A2_10__aw2_U3 ( .A(round_inst_sout_w[41]), .B(
        round_inst_xin_w[43]), .ZN(round_inst_A2_10__aw2_n5) );
  INV_X1 round_inst_A2_10__aw2_U2 ( .A(round_inst_sout_w[43]), .ZN(
        round_inst_xin_w[42]) );
  INV_X1 round_inst_A2_10__aw2_U1 ( .A(round_inst_sout_w[41]), .ZN(
        round_inst_xin_w[40]) );
  XNOR2_X1 round_inst_A2_10__ax2_U2 ( .A(round_inst_A2_10__ax2_n3), .B(
        round_inst_sout_x[40]), .ZN(round_inst_srout2_x[25]) );
  XNOR2_X1 round_inst_A2_10__ax2_U1 ( .A(round_inst_srout2_x[24]), .B(
        round_inst_srout2_x[27]), .ZN(round_inst_A2_10__ax2_n3) );
  XNOR2_X1 round_inst_A2_10__ay2_U2 ( .A(round_inst_A2_10__ay2_n3), .B(
        round_inst_sout_y[40]), .ZN(round_inst_srout2_y[25]) );
  XNOR2_X1 round_inst_A2_10__ay2_U1 ( .A(round_inst_srout2_y[24]), .B(
        round_inst_srout2_y[27]), .ZN(round_inst_A2_10__ay2_n3) );
  XNOR2_X1 round_inst_A2_10__az2_U2 ( .A(round_inst_A2_10__az2_n3), .B(
        round_inst_sout_z[40]), .ZN(round_inst_srout2_z[25]) );
  XNOR2_X1 round_inst_A2_10__az2_U1 ( .A(round_inst_srout2_z[24]), .B(
        round_inst_srout2_z[27]), .ZN(round_inst_A2_10__az2_n3) );
  XNOR2_X1 round_inst_A2_11__aw2_U4 ( .A(round_inst_A2_11__aw2_n5), .B(
        round_inst_sout_w[44]), .ZN(round_inst_xin_w[45]) );
  XNOR2_X1 round_inst_A2_11__aw2_U3 ( .A(round_inst_sout_w[45]), .B(
        round_inst_xin_w[47]), .ZN(round_inst_A2_11__aw2_n5) );
  INV_X1 round_inst_A2_11__aw2_U2 ( .A(round_inst_sout_w[47]), .ZN(
        round_inst_xin_w[46]) );
  INV_X1 round_inst_A2_11__aw2_U1 ( .A(round_inst_sout_w[45]), .ZN(
        round_inst_xin_w[44]) );
  XNOR2_X1 round_inst_A2_11__ax2_U2 ( .A(round_inst_A2_11__ax2_n3), .B(
        round_inst_sout_x[44]), .ZN(round_inst_srout2_x[45]) );
  XNOR2_X1 round_inst_A2_11__ax2_U1 ( .A(round_inst_srout2_x[44]), .B(
        round_inst_srout2_x[47]), .ZN(round_inst_A2_11__ax2_n3) );
  XNOR2_X1 round_inst_A2_11__ay2_U2 ( .A(round_inst_A2_11__ay2_n3), .B(
        round_inst_sout_y[44]), .ZN(round_inst_srout2_y[45]) );
  XNOR2_X1 round_inst_A2_11__ay2_U1 ( .A(round_inst_srout2_y[44]), .B(
        round_inst_srout2_y[47]), .ZN(round_inst_A2_11__ay2_n3) );
  XNOR2_X1 round_inst_A2_11__az2_U2 ( .A(round_inst_A2_11__az2_n3), .B(
        round_inst_sout_z[44]), .ZN(round_inst_srout2_z[45]) );
  XNOR2_X1 round_inst_A2_11__az2_U1 ( .A(round_inst_srout2_z[44]), .B(
        round_inst_srout2_z[47]), .ZN(round_inst_A2_11__az2_n3) );
  XNOR2_X1 round_inst_A2_12__aw2_U4 ( .A(round_inst_A2_12__aw2_n5), .B(
        round_inst_sout_w[48]), .ZN(round_inst_xin_w[49]) );
  XNOR2_X1 round_inst_A2_12__aw2_U3 ( .A(round_inst_sout_w[49]), .B(
        round_inst_xin_w[51]), .ZN(round_inst_A2_12__aw2_n5) );
  INV_X1 round_inst_A2_12__aw2_U2 ( .A(round_inst_sout_w[51]), .ZN(
        round_inst_xin_w[50]) );
  INV_X1 round_inst_A2_12__aw2_U1 ( .A(round_inst_sout_w[49]), .ZN(
        round_inst_xin_w[48]) );
  XNOR2_X1 round_inst_A2_12__ax2_U2 ( .A(round_inst_A2_12__ax2_n3), .B(
        round_inst_sout_x[48]), .ZN(round_inst_srout2_x[1]) );
  XNOR2_X1 round_inst_A2_12__ax2_U1 ( .A(round_inst_srout2_x[0]), .B(
        round_inst_srout2_x[3]), .ZN(round_inst_A2_12__ax2_n3) );
  XNOR2_X1 round_inst_A2_12__ay2_U2 ( .A(round_inst_A2_12__ay2_n3), .B(
        round_inst_sout_y[48]), .ZN(round_inst_srout2_y[1]) );
  XNOR2_X1 round_inst_A2_12__ay2_U1 ( .A(round_inst_srout2_y[0]), .B(
        round_inst_srout2_y[3]), .ZN(round_inst_A2_12__ay2_n3) );
  XNOR2_X1 round_inst_A2_12__az2_U2 ( .A(round_inst_A2_12__az2_n3), .B(
        round_inst_sout_z[48]), .ZN(round_inst_srout2_z[1]) );
  XNOR2_X1 round_inst_A2_12__az2_U1 ( .A(round_inst_srout2_z[0]), .B(
        round_inst_srout2_z[3]), .ZN(round_inst_A2_12__az2_n3) );
  XNOR2_X1 round_inst_A2_13__aw2_U4 ( .A(round_inst_A2_13__aw2_n5), .B(
        round_inst_sout_w[52]), .ZN(round_inst_xin_w[53]) );
  XNOR2_X1 round_inst_A2_13__aw2_U3 ( .A(round_inst_sout_w[53]), .B(
        round_inst_xin_w[55]), .ZN(round_inst_A2_13__aw2_n5) );
  INV_X1 round_inst_A2_13__aw2_U2 ( .A(round_inst_sout_w[55]), .ZN(
        round_inst_xin_w[54]) );
  INV_X1 round_inst_A2_13__aw2_U1 ( .A(round_inst_sout_w[53]), .ZN(
        round_inst_xin_w[52]) );
  XNOR2_X1 round_inst_A2_13__ax2_U2 ( .A(round_inst_A2_13__ax2_n3), .B(
        round_inst_sout_x[52]), .ZN(round_inst_srout2_x[21]) );
  XNOR2_X1 round_inst_A2_13__ax2_U1 ( .A(round_inst_srout2_x[20]), .B(
        round_inst_srout2_x[23]), .ZN(round_inst_A2_13__ax2_n3) );
  XNOR2_X1 round_inst_A2_13__ay2_U2 ( .A(round_inst_A2_13__ay2_n3), .B(
        round_inst_sout_y[52]), .ZN(round_inst_srout2_y[21]) );
  XNOR2_X1 round_inst_A2_13__ay2_U1 ( .A(round_inst_srout2_y[20]), .B(
        round_inst_srout2_y[23]), .ZN(round_inst_A2_13__ay2_n3) );
  XNOR2_X1 round_inst_A2_13__az2_U2 ( .A(round_inst_A2_13__az2_n3), .B(
        round_inst_sout_z[52]), .ZN(round_inst_srout2_z[21]) );
  XNOR2_X1 round_inst_A2_13__az2_U1 ( .A(round_inst_srout2_z[20]), .B(
        round_inst_srout2_z[23]), .ZN(round_inst_A2_13__az2_n3) );
  XNOR2_X1 round_inst_A2_14__aw2_U4 ( .A(round_inst_A2_14__aw2_n5), .B(
        round_inst_sout_w[56]), .ZN(round_inst_xin_w[57]) );
  XNOR2_X1 round_inst_A2_14__aw2_U3 ( .A(round_inst_sout_w[57]), .B(
        round_inst_xin_w[59]), .ZN(round_inst_A2_14__aw2_n5) );
  INV_X1 round_inst_A2_14__aw2_U2 ( .A(round_inst_sout_w[59]), .ZN(
        round_inst_xin_w[58]) );
  INV_X1 round_inst_A2_14__aw2_U1 ( .A(round_inst_sout_w[57]), .ZN(
        round_inst_xin_w[56]) );
  XNOR2_X1 round_inst_A2_14__ax2_U2 ( .A(round_inst_A2_14__ax2_n3), .B(
        round_inst_sout_x[56]), .ZN(round_inst_srout2_x[41]) );
  XNOR2_X1 round_inst_A2_14__ax2_U1 ( .A(round_inst_srout2_x[40]), .B(
        round_inst_srout2_x[43]), .ZN(round_inst_A2_14__ax2_n3) );
  XNOR2_X1 round_inst_A2_14__ay2_U2 ( .A(round_inst_A2_14__ay2_n3), .B(
        round_inst_sout_y[56]), .ZN(round_inst_srout2_y[41]) );
  XNOR2_X1 round_inst_A2_14__ay2_U1 ( .A(round_inst_srout2_y[40]), .B(
        round_inst_srout2_y[43]), .ZN(round_inst_A2_14__ay2_n3) );
  XNOR2_X1 round_inst_A2_14__az2_U2 ( .A(round_inst_A2_14__az2_n3), .B(
        round_inst_sout_z[56]), .ZN(round_inst_srout2_z[41]) );
  XNOR2_X1 round_inst_A2_14__az2_U1 ( .A(round_inst_srout2_z[40]), .B(
        round_inst_srout2_z[43]), .ZN(round_inst_A2_14__az2_n3) );
  XNOR2_X1 round_inst_A2_15__aw2_U4 ( .A(round_inst_A2_15__aw2_n5), .B(
        round_inst_sout_w[60]), .ZN(round_inst_xin_w[61]) );
  XNOR2_X1 round_inst_A2_15__aw2_U3 ( .A(round_inst_sout_w[61]), .B(
        round_inst_xin_w[63]), .ZN(round_inst_A2_15__aw2_n5) );
  INV_X1 round_inst_A2_15__aw2_U2 ( .A(round_inst_sout_w[63]), .ZN(
        round_inst_xin_w[62]) );
  INV_X1 round_inst_A2_15__aw2_U1 ( .A(round_inst_sout_w[61]), .ZN(
        round_inst_xin_w[60]) );
  XNOR2_X1 round_inst_A2_15__ax2_U2 ( .A(round_inst_A2_15__ax2_n3), .B(
        round_inst_sout_x[60]), .ZN(round_inst_srout2_x[61]) );
  XNOR2_X1 round_inst_A2_15__ax2_U1 ( .A(round_inst_srout2_x[60]), .B(
        round_inst_srout2_x[63]), .ZN(round_inst_A2_15__ax2_n3) );
  XNOR2_X1 round_inst_A2_15__ay2_U2 ( .A(round_inst_A2_15__ay2_n3), .B(
        round_inst_sout_y[60]), .ZN(round_inst_srout2_y[61]) );
  XNOR2_X1 round_inst_A2_15__ay2_U1 ( .A(round_inst_srout2_y[60]), .B(
        round_inst_srout2_y[63]), .ZN(round_inst_A2_15__ay2_n3) );
  XNOR2_X1 round_inst_A2_15__az2_U2 ( .A(round_inst_A2_15__az2_n3), .B(
        round_inst_sout_z[60]), .ZN(round_inst_srout2_z[61]) );
  XNOR2_X1 round_inst_A2_15__az2_U1 ( .A(round_inst_srout2_z[60]), .B(
        round_inst_srout2_z[63]), .ZN(round_inst_A2_15__az2_n3) );
  MUX2_X1 round_inst_mux_inv_w2_U68 ( .A(round_inst_srout2_w[1]), .B(
        round_inst_sout_w[1]), .S(inv_sig), .Z(round_inst_min_w[1]) );
  MUX2_X1 round_inst_mux_inv_w2_U67 ( .A(round_inst_srout2_w[3]), .B(
        round_inst_sout_w[3]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[3]) );
  MUX2_X1 round_inst_mux_inv_w2_U66 ( .A(round_inst_srout2_w[2]), .B(
        round_inst_xin_w[3]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[2]) );
  MUX2_X1 round_inst_mux_inv_w2_U65 ( .A(round_inst_srout2_w[15]), .B(
        round_inst_sout_w[15]), .S(inv_sig), .Z(round_inst_min_w[15]) );
  MUX2_X1 round_inst_mux_inv_w2_U64 ( .A(round_inst_srout2_w[51]), .B(
        round_inst_sout_w[51]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[51]) );
  MUX2_X1 round_inst_mux_inv_w2_U63 ( .A(round_inst_srout2_w[11]), .B(
        round_inst_sout_w[11]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[11]) );
  MUX2_X1 round_inst_mux_inv_w2_U62 ( .A(round_inst_srout2_w[55]), .B(
        round_inst_sout_w[55]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[55]) );
  MUX2_X1 round_inst_mux_inv_w2_U61 ( .A(round_inst_srout2_w[57]), .B(
        round_inst_sout_w[57]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[57]) );
  MUX2_X1 round_inst_mux_inv_w2_U60 ( .A(round_inst_srout2_w[49]), .B(
        round_inst_sout_w[49]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[49]) );
  MUX2_X1 round_inst_mux_inv_w2_U59 ( .A(round_inst_srout2_w[37]), .B(
        round_inst_sout_w[37]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[37]) );
  MUX2_X1 round_inst_mux_inv_w2_U58 ( .A(round_inst_srout2_w[33]), .B(
        round_inst_sout_w[33]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[33]) );
  MUX2_X1 round_inst_mux_inv_w2_U57 ( .A(round_inst_srout2_w[17]), .B(
        round_inst_sout_w[17]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[17]) );
  MUX2_X1 round_inst_mux_inv_w2_U56 ( .A(round_inst_srout2_w[25]), .B(
        round_inst_sout_w[25]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[25]) );
  MUX2_X1 round_inst_mux_inv_w2_U55 ( .A(round_inst_srout2_w[13]), .B(
        round_inst_sout_w[13]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[13]) );
  MUX2_X1 round_inst_mux_inv_w2_U54 ( .A(round_inst_srout2_w[50]), .B(
        round_inst_xin_w[51]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[50]) );
  MUX2_X1 round_inst_mux_inv_w2_U53 ( .A(round_inst_srout2_w[52]), .B(
        round_inst_sout_w[52]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[52]) );
  INV_X1 round_inst_mux_inv_w2_U52 ( .A(round_inst_mux_inv_w2_n263), .ZN(
        round_inst_mux_inv_w2_n266) );
  MUX2_X1 round_inst_mux_inv_w2_U51 ( .A(round_inst_srout2_w[54]), .B(
        round_inst_xin_w[55]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[54]) );
  MUX2_X1 round_inst_mux_inv_w2_U50 ( .A(round_inst_srout2_w[48]), .B(
        round_inst_sout_w[48]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[48]) );
  MUX2_X1 round_inst_mux_inv_w2_U49 ( .A(round_inst_srout2_w[34]), .B(
        round_inst_xin_w[35]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[34]) );
  MUX2_X1 round_inst_mux_inv_w2_U48 ( .A(round_inst_srout2_w[40]), .B(
        round_inst_sout_w[40]), .S(inv_sig), .Z(round_inst_min_w[40]) );
  MUX2_X1 round_inst_mux_inv_w2_U47 ( .A(round_inst_srout2_w[38]), .B(
        round_inst_xin_w[39]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[38]) );
  MUX2_X1 round_inst_mux_inv_w2_U46 ( .A(round_inst_srout2_w[32]), .B(
        round_inst_sout_w[32]), .S(inv_sig), .Z(round_inst_min_w[32]) );
  MUX2_X1 round_inst_mux_inv_w2_U45 ( .A(round_inst_srout2_w[16]), .B(
        round_inst_sout_w[16]), .S(inv_sig), .Z(round_inst_min_w[16]) );
  MUX2_X1 round_inst_mux_inv_w2_U44 ( .A(round_inst_srout2_w[26]), .B(
        round_inst_xin_w[27]), .S(inv_sig), .Z(round_inst_min_w[26]) );
  MUX2_X1 round_inst_mux_inv_w2_U43 ( .A(round_inst_srout2_w[20]), .B(
        round_inst_sout_w[20]), .S(round_inst_mux_inv_w2_n266), .Z(
        round_inst_min_w[20]) );
  MUX2_X1 round_inst_mux_inv_w2_U42 ( .A(round_inst_srout2_w[14]), .B(
        round_inst_xin_w[15]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[14]) );
  MUX2_X1 round_inst_mux_inv_w2_U41 ( .A(round_inst_srout2_w[12]), .B(
        round_inst_sout_w[12]), .S(inv_sig), .Z(round_inst_min_w[12]) );
  MUX2_X1 round_inst_mux_inv_w2_U40 ( .A(round_inst_srout2_w[10]), .B(
        round_inst_xin_w[11]), .S(inv_sig), .Z(round_inst_min_w[10]) );
  MUX2_X1 round_inst_mux_inv_w2_U39 ( .A(round_inst_srout2_w[0]), .B(
        round_inst_sout_w[0]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[0]) );
  MUX2_X1 round_inst_mux_inv_w2_U38 ( .A(round_inst_srout2_w[63]), .B(
        round_inst_sout_w[63]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[63]) );
  MUX2_X1 round_inst_mux_inv_w2_U37 ( .A(round_inst_srout2_w[47]), .B(
        round_inst_sout_w[47]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[47]) );
  MUX2_X1 round_inst_mux_inv_w2_U36 ( .A(round_inst_srout2_w[7]), .B(
        round_inst_sout_w[7]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[7]) );
  MUX2_X1 round_inst_mux_inv_w2_U35 ( .A(round_inst_srout2_w[59]), .B(
        round_inst_sout_w[59]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[59]) );
  MUX2_X1 round_inst_mux_inv_w2_U34 ( .A(round_inst_srout2_w[61]), .B(
        round_inst_sout_w[61]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[61]) );
  MUX2_X1 round_inst_mux_inv_w2_U33 ( .A(round_inst_srout2_w[53]), .B(
        round_inst_sout_w[53]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[53]) );
  MUX2_X1 round_inst_mux_inv_w2_U32 ( .A(round_inst_srout2_w[45]), .B(
        round_inst_sout_w[45]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[45]) );
  MUX2_X1 round_inst_mux_inv_w2_U31 ( .A(round_inst_srout2_w[41]), .B(
        round_inst_sout_w[41]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[41]) );
  MUX2_X1 round_inst_mux_inv_w2_U30 ( .A(round_inst_srout2_w[21]), .B(
        round_inst_sout_w[21]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[21]) );
  MUX2_X1 round_inst_mux_inv_w2_U29 ( .A(round_inst_srout2_w[29]), .B(
        round_inst_sout_w[29]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[29]) );
  MUX2_X1 round_inst_mux_inv_w2_U28 ( .A(round_inst_srout2_w[9]), .B(
        round_inst_sout_w[9]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[9]) );
  MUX2_X1 round_inst_mux_inv_w2_U27 ( .A(round_inst_srout2_w[5]), .B(
        round_inst_sout_w[5]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[5]) );
  MUX2_X1 round_inst_mux_inv_w2_U26 ( .A(round_inst_srout2_w[62]), .B(
        round_inst_xin_w[63]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[62]) );
  MUX2_X1 round_inst_mux_inv_w2_U25 ( .A(round_inst_srout2_w[58]), .B(
        round_inst_xin_w[59]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[58]) );
  MUX2_X1 round_inst_mux_inv_w2_U24 ( .A(round_inst_srout2_w[56]), .B(
        round_inst_sout_w[56]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[56]) );
  MUX2_X1 round_inst_mux_inv_w2_U23 ( .A(round_inst_srout2_w[42]), .B(
        round_inst_xin_w[43]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[42]) );
  MUX2_X1 round_inst_mux_inv_w2_U22 ( .A(round_inst_srout2_w[46]), .B(
        round_inst_xin_w[47]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[46]) );
  MUX2_X1 round_inst_mux_inv_w2_U21 ( .A(round_inst_srout2_w[22]), .B(
        round_inst_xin_w[23]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[22]) );
  MUX2_X1 round_inst_mux_inv_w2_U20 ( .A(round_inst_srout2_w[28]), .B(
        round_inst_sout_w[28]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[28]) );
  MUX2_X1 round_inst_mux_inv_w2_U19 ( .A(round_inst_srout2_w[24]), .B(
        round_inst_sout_w[24]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[24]) );
  MUX2_X1 round_inst_mux_inv_w2_U18 ( .A(round_inst_srout2_w[8]), .B(
        round_inst_sout_w[8]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[8]) );
  MUX2_X1 round_inst_mux_inv_w2_U17 ( .A(round_inst_srout2_w[4]), .B(
        round_inst_sout_w[4]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[4]) );
  MUX2_X1 round_inst_mux_inv_w2_U16 ( .A(round_inst_srout2_w[60]), .B(
        round_inst_sout_w[60]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[60]) );
  MUX2_X1 round_inst_mux_inv_w2_U15 ( .A(round_inst_srout2_w[44]), .B(
        round_inst_sout_w[44]), .S(inv_sig), .Z(round_inst_min_w[44]) );
  MUX2_X1 round_inst_mux_inv_w2_U14 ( .A(round_inst_srout2_w[36]), .B(
        round_inst_sout_w[36]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[36]) );
  MUX2_X1 round_inst_mux_inv_w2_U13 ( .A(round_inst_srout2_w[30]), .B(
        round_inst_xin_w[31]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[30]) );
  MUX2_X1 round_inst_mux_inv_w2_U12 ( .A(round_inst_srout2_w[6]), .B(
        round_inst_xin_w[7]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[6]) );
  MUX2_X1 round_inst_mux_inv_w2_U11 ( .A(round_inst_srout2_w[18]), .B(
        round_inst_xin_w[19]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[18]) );
  MUX2_X1 round_inst_mux_inv_w2_U10 ( .A(round_inst_srout2_w[39]), .B(
        round_inst_sout_w[39]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[39]) );
  MUX2_X1 round_inst_mux_inv_w2_U9 ( .A(round_inst_srout2_w[43]), .B(
        round_inst_sout_w[43]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[43]) );
  MUX2_X1 round_inst_mux_inv_w2_U8 ( .A(round_inst_srout2_w[35]), .B(
        round_inst_sout_w[35]), .S(inv_sig), .Z(round_inst_min_w[35]) );
  MUX2_X1 round_inst_mux_inv_w2_U7 ( .A(round_inst_srout2_w[23]), .B(
        round_inst_sout_w[23]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[23]) );
  MUX2_X1 round_inst_mux_inv_w2_U6 ( .A(round_inst_srout2_w[27]), .B(
        round_inst_sout_w[27]), .S(round_inst_mux_inv_w2_n264), .Z(
        round_inst_min_w[27]) );
  INV_X1 round_inst_mux_inv_w2_U5 ( .A(round_inst_mux_inv_w2_n263), .ZN(
        round_inst_mux_inv_w2_n264) );
  MUX2_X1 round_inst_mux_inv_w2_U4 ( .A(round_inst_srout2_w[19]), .B(
        round_inst_sout_w[19]), .S(inv_sig), .Z(round_inst_min_w[19]) );
  MUX2_X1 round_inst_mux_inv_w2_U3 ( .A(round_inst_srout2_w[31]), .B(
        round_inst_sout_w[31]), .S(round_inst_mux_inv_w2_n265), .Z(
        round_inst_min_w[31]) );
  INV_X1 round_inst_mux_inv_w2_U2 ( .A(round_inst_mux_inv_w2_n263), .ZN(
        round_inst_mux_inv_w2_n265) );
  INV_X1 round_inst_mux_inv_w2_U1 ( .A(inv_sig), .ZN(
        round_inst_mux_inv_w2_n263) );
  MUX2_X1 round_inst_mux_inv_x2_U69 ( .A(round_inst_srout2_x[18]), .B(
        round_inst_srout2_x[35]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[18]) );
  MUX2_X1 round_inst_mux_inv_x2_U68 ( .A(round_inst_srout2_x[2]), .B(
        round_inst_srout2_x[19]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[2]) );
  MUX2_X1 round_inst_mux_inv_x2_U67 ( .A(round_inst_srout2_x[3]), .B(
        round_inst_srout2_x[18]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[3]) );
  MUX2_X1 round_inst_mux_inv_x2_U66 ( .A(round_inst_srout2_x[19]), .B(
        round_inst_srout2_x[34]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[19]) );
  MUX2_X1 round_inst_mux_inv_x2_U65 ( .A(round_inst_srout2_x[1]), .B(
        round_inst_srout2_x[16]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[1]) );
  MUX2_X1 round_inst_mux_inv_x2_U64 ( .A(round_inst_srout2_x[17]), .B(
        round_inst_srout2_x[32]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[17]) );
  MUX2_X1 round_inst_mux_inv_x2_U63 ( .A(round_inst_srout2_x[50]), .B(
        round_inst_srout2_x[3]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[50]) );
  MUX2_X1 round_inst_mux_inv_x2_U62 ( .A(round_inst_srout2_x[54]), .B(
        round_inst_srout2_x[23]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[54]) );
  MUX2_X1 round_inst_mux_inv_x2_U61 ( .A(round_inst_srout2_x[34]), .B(
        round_inst_srout2_x[51]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[34]) );
  MUX2_X1 round_inst_mux_inv_x2_U60 ( .A(round_inst_srout2_x[38]), .B(
        round_inst_srout2_x[7]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[38]) );
  MUX2_X1 round_inst_mux_inv_x2_U59 ( .A(round_inst_srout2_x[26]), .B(
        round_inst_srout2_x[11]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[26]) );
  MUX2_X1 round_inst_mux_inv_x2_U58 ( .A(round_inst_srout2_x[14]), .B(
        round_inst_srout2_x[15]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[14]) );
  MUX2_X1 round_inst_mux_inv_x2_U57 ( .A(round_inst_srout2_x[10]), .B(
        round_inst_srout2_x[59]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[10]) );
  MUX2_X1 round_inst_mux_inv_x2_U56 ( .A(round_inst_srout2_x[62]), .B(
        round_inst_srout2_x[63]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[62]) );
  MUX2_X1 round_inst_mux_inv_x2_U55 ( .A(round_inst_srout2_x[58]), .B(
        round_inst_srout2_x[43]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[58]) );
  MUX2_X1 round_inst_mux_inv_x2_U54 ( .A(round_inst_srout2_x[42]), .B(
        round_inst_srout2_x[27]), .S(round_inst_mux_inv_x2_n267), .Z(
        round_inst_min_x[42]) );
  INV_X1 round_inst_mux_inv_x2_U53 ( .A(round_inst_mux_inv_x2_n265), .ZN(
        round_inst_mux_inv_x2_n267) );
  MUX2_X1 round_inst_mux_inv_x2_U52 ( .A(round_inst_srout2_x[46]), .B(
        round_inst_srout2_x[47]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[46]) );
  MUX2_X1 round_inst_mux_inv_x2_U51 ( .A(round_inst_srout2_x[22]), .B(
        round_inst_srout2_x[55]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[22]) );
  MUX2_X1 round_inst_mux_inv_x2_U50 ( .A(round_inst_srout2_x[30]), .B(
        round_inst_srout2_x[31]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[30]) );
  MUX2_X1 round_inst_mux_inv_x2_U49 ( .A(round_inst_srout2_x[6]), .B(
        round_inst_srout2_x[39]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[6]) );
  MUX2_X1 round_inst_mux_inv_x2_U48 ( .A(round_inst_srout2_x[51]), .B(
        round_inst_srout2_x[2]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[51]) );
  MUX2_X1 round_inst_mux_inv_x2_U47 ( .A(round_inst_srout2_x[39]), .B(
        round_inst_srout2_x[6]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[39]) );
  MUX2_X1 round_inst_mux_inv_x2_U46 ( .A(round_inst_srout2_x[23]), .B(
        round_inst_srout2_x[54]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[23]) );
  MUX2_X1 round_inst_mux_inv_x2_U45 ( .A(round_inst_srout2_x[15]), .B(
        round_inst_srout2_x[14]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[15]) );
  MUX2_X1 round_inst_mux_inv_x2_U44 ( .A(round_inst_srout2_x[16]), .B(
        round_inst_sout_x[16]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[16]) );
  MUX2_X1 round_inst_mux_inv_x2_U43 ( .A(round_inst_srout2_x[52]), .B(
        round_inst_sout_x[52]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[52]) );
  MUX2_X1 round_inst_mux_inv_x2_U42 ( .A(round_inst_srout2_x[48]), .B(
        round_inst_sout_x[48]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[48]) );
  MUX2_X1 round_inst_mux_inv_x2_U41 ( .A(round_inst_srout2_x[40]), .B(
        round_inst_sout_x[40]), .S(round_inst_mux_inv_x2_n266), .Z(
        round_inst_min_x[40]) );
  INV_X1 round_inst_mux_inv_x2_U40 ( .A(round_inst_mux_inv_x2_n265), .ZN(
        round_inst_mux_inv_x2_n266) );
  INV_X1 round_inst_mux_inv_x2_U39 ( .A(inv_sig), .ZN(
        round_inst_mux_inv_x2_n265) );
  MUX2_X1 round_inst_mux_inv_x2_U38 ( .A(round_inst_srout2_x[32]), .B(
        round_inst_sout_x[32]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[32]) );
  MUX2_X1 round_inst_mux_inv_x2_U37 ( .A(round_inst_srout2_x[20]), .B(
        round_inst_sout_x[20]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[20]) );
  MUX2_X1 round_inst_mux_inv_x2_U36 ( .A(round_inst_srout2_x[12]), .B(
        round_inst_sout_x[12]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[12]) );
  MUX2_X1 round_inst_mux_inv_x2_U35 ( .A(round_inst_srout2_x[0]), .B(
        round_inst_sout_x[0]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[0]) );
  MUX2_X1 round_inst_mux_inv_x2_U34 ( .A(round_inst_srout2_x[59]), .B(
        round_inst_srout2_x[42]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[59]) );
  MUX2_X1 round_inst_mux_inv_x2_U33 ( .A(round_inst_srout2_x[63]), .B(
        round_inst_srout2_x[62]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[63]) );
  MUX2_X1 round_inst_mux_inv_x2_U32 ( .A(round_inst_srout2_x[43]), .B(
        round_inst_srout2_x[26]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[43]) );
  MUX2_X1 round_inst_mux_inv_x2_U31 ( .A(round_inst_srout2_x[47]), .B(
        round_inst_srout2_x[46]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[47]) );
  MUX2_X1 round_inst_mux_inv_x2_U30 ( .A(round_inst_srout2_x[27]), .B(
        round_inst_srout2_x[10]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[27]) );
  MUX2_X1 round_inst_mux_inv_x2_U29 ( .A(round_inst_srout2_x[31]), .B(
        round_inst_srout2_x[30]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[31]) );
  MUX2_X1 round_inst_mux_inv_x2_U28 ( .A(round_inst_srout2_x[7]), .B(
        round_inst_srout2_x[38]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[7]) );
  MUX2_X1 round_inst_mux_inv_x2_U27 ( .A(round_inst_srout2_x[60]), .B(
        round_inst_sout_x[60]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[60]) );
  MUX2_X1 round_inst_mux_inv_x2_U26 ( .A(round_inst_srout2_x[56]), .B(
        round_inst_sout_x[56]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[56]) );
  MUX2_X1 round_inst_mux_inv_x2_U25 ( .A(round_inst_srout2_x[44]), .B(
        round_inst_sout_x[44]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[44]) );
  MUX2_X1 round_inst_mux_inv_x2_U24 ( .A(round_inst_srout2_x[36]), .B(
        round_inst_sout_x[36]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[36]) );
  MUX2_X1 round_inst_mux_inv_x2_U23 ( .A(round_inst_srout2_x[28]), .B(
        round_inst_sout_x[28]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[28]) );
  MUX2_X1 round_inst_mux_inv_x2_U22 ( .A(round_inst_srout2_x[24]), .B(
        round_inst_sout_x[24]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[24]) );
  MUX2_X1 round_inst_mux_inv_x2_U21 ( .A(round_inst_srout2_x[8]), .B(
        round_inst_sout_x[8]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[8]) );
  MUX2_X1 round_inst_mux_inv_x2_U20 ( .A(round_inst_srout2_x[4]), .B(
        round_inst_sout_x[4]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[4]) );
  MUX2_X1 round_inst_mux_inv_x2_U19 ( .A(round_inst_srout2_x[55]), .B(
        round_inst_srout2_x[22]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[55]) );
  MUX2_X1 round_inst_mux_inv_x2_U18 ( .A(round_inst_srout2_x[35]), .B(
        round_inst_srout2_x[50]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[35]) );
  MUX2_X1 round_inst_mux_inv_x2_U17 ( .A(round_inst_srout2_x[11]), .B(
        round_inst_srout2_x[58]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[11]) );
  MUX2_X1 round_inst_mux_inv_x2_U16 ( .A(round_inst_srout2_x[57]), .B(
        round_inst_srout2_x[40]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[57]) );
  MUX2_X1 round_inst_mux_inv_x2_U15 ( .A(round_inst_srout2_x[49]), .B(
        round_inst_srout2_x[0]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[49]) );
  MUX2_X1 round_inst_mux_inv_x2_U14 ( .A(round_inst_srout2_x[37]), .B(
        round_inst_srout2_x[4]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[37]) );
  MUX2_X1 round_inst_mux_inv_x2_U13 ( .A(round_inst_srout2_x[33]), .B(
        round_inst_srout2_x[48]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[33]) );
  MUX2_X1 round_inst_mux_inv_x2_U12 ( .A(round_inst_srout2_x[25]), .B(
        round_inst_srout2_x[8]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[25]) );
  MUX2_X1 round_inst_mux_inv_x2_U11 ( .A(round_inst_srout2_x[13]), .B(
        round_inst_srout2_x[12]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[13]) );
  MUX2_X1 round_inst_mux_inv_x2_U10 ( .A(round_inst_srout2_x[61]), .B(
        round_inst_srout2_x[60]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[61]) );
  MUX2_X1 round_inst_mux_inv_x2_U9 ( .A(round_inst_srout2_x[53]), .B(
        round_inst_srout2_x[20]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[53]) );
  MUX2_X1 round_inst_mux_inv_x2_U8 ( .A(round_inst_srout2_x[45]), .B(
        round_inst_srout2_x[44]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[45]) );
  MUX2_X1 round_inst_mux_inv_x2_U7 ( .A(round_inst_srout2_x[41]), .B(
        round_inst_srout2_x[24]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[41]) );
  MUX2_X1 round_inst_mux_inv_x2_U6 ( .A(round_inst_srout2_x[21]), .B(
        round_inst_srout2_x[52]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[21]) );
  MUX2_X1 round_inst_mux_inv_x2_U5 ( .A(round_inst_srout2_x[29]), .B(
        round_inst_srout2_x[28]), .S(round_inst_mux_inv_x2_n263), .Z(
        round_inst_min_x[29]) );
  INV_X1 round_inst_mux_inv_x2_U4 ( .A(round_inst_mux_inv_x2_n265), .ZN(
        round_inst_mux_inv_x2_n263) );
  MUX2_X1 round_inst_mux_inv_x2_U3 ( .A(round_inst_srout2_x[9]), .B(
        round_inst_srout2_x[56]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[9]) );
  MUX2_X1 round_inst_mux_inv_x2_U2 ( .A(round_inst_srout2_x[5]), .B(
        round_inst_srout2_x[36]), .S(round_inst_mux_inv_x2_n264), .Z(
        round_inst_min_x[5]) );
  INV_X1 round_inst_mux_inv_x2_U1 ( .A(round_inst_mux_inv_x2_n265), .ZN(
        round_inst_mux_inv_x2_n264) );
  MUX2_X1 round_inst_mux_inv_y2_U69 ( .A(round_inst_srout2_y[18]), .B(
        round_inst_srout2_y[35]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[18]) );
  MUX2_X1 round_inst_mux_inv_y2_U68 ( .A(round_inst_srout2_y[2]), .B(
        round_inst_srout2_y[19]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[2]) );
  MUX2_X1 round_inst_mux_inv_y2_U67 ( .A(round_inst_srout2_y[19]), .B(
        round_inst_srout2_y[34]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[19]) );
  MUX2_X1 round_inst_mux_inv_y2_U66 ( .A(round_inst_srout2_y[3]), .B(
        round_inst_srout2_y[18]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[3]) );
  MUX2_X1 round_inst_mux_inv_y2_U65 ( .A(round_inst_srout2_y[1]), .B(
        round_inst_srout2_y[16]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[1]) );
  MUX2_X1 round_inst_mux_inv_y2_U64 ( .A(round_inst_srout2_y[57]), .B(
        round_inst_srout2_y[40]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[57]) );
  MUX2_X1 round_inst_mux_inv_y2_U63 ( .A(round_inst_srout2_y[49]), .B(
        round_inst_srout2_y[0]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[49]) );
  MUX2_X1 round_inst_mux_inv_y2_U62 ( .A(round_inst_srout2_y[33]), .B(
        round_inst_srout2_y[48]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[33]) );
  MUX2_X1 round_inst_mux_inv_y2_U61 ( .A(round_inst_srout2_y[17]), .B(
        round_inst_srout2_y[32]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[17]) );
  MUX2_X1 round_inst_mux_inv_y2_U60 ( .A(round_inst_srout2_y[25]), .B(
        round_inst_srout2_y[8]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[25]) );
  MUX2_X1 round_inst_mux_inv_y2_U59 ( .A(round_inst_srout2_y[45]), .B(
        round_inst_srout2_y[44]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[45]) );
  MUX2_X1 round_inst_mux_inv_y2_U58 ( .A(round_inst_srout2_y[29]), .B(
        round_inst_srout2_y[28]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[29]) );
  MUX2_X1 round_inst_mux_inv_y2_U57 ( .A(round_inst_srout2_y[5]), .B(
        round_inst_srout2_y[36]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[5]) );
  MUX2_X1 round_inst_mux_inv_y2_U56 ( .A(round_inst_srout2_y[50]), .B(
        round_inst_srout2_y[3]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[50]) );
  MUX2_X1 round_inst_mux_inv_y2_U55 ( .A(round_inst_srout2_y[54]), .B(
        round_inst_srout2_y[23]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[54]) );
  MUX2_X1 round_inst_mux_inv_y2_U54 ( .A(round_inst_srout2_y[34]), .B(
        round_inst_srout2_y[51]), .S(round_inst_mux_inv_y2_n267), .Z(
        round_inst_min_y[34]) );
  INV_X1 round_inst_mux_inv_y2_U53 ( .A(round_inst_mux_inv_y2_n263), .ZN(
        round_inst_mux_inv_y2_n267) );
  MUX2_X1 round_inst_mux_inv_y2_U52 ( .A(round_inst_srout2_y[38]), .B(
        round_inst_srout2_y[7]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[38]) );
  MUX2_X1 round_inst_mux_inv_y2_U51 ( .A(round_inst_srout2_y[26]), .B(
        round_inst_srout2_y[11]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[26]) );
  MUX2_X1 round_inst_mux_inv_y2_U50 ( .A(round_inst_srout2_y[14]), .B(
        round_inst_srout2_y[15]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[14]) );
  MUX2_X1 round_inst_mux_inv_y2_U49 ( .A(round_inst_srout2_y[10]), .B(
        round_inst_srout2_y[59]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[10]) );
  MUX2_X1 round_inst_mux_inv_y2_U48 ( .A(round_inst_srout2_y[62]), .B(
        round_inst_srout2_y[63]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[62]) );
  MUX2_X1 round_inst_mux_inv_y2_U47 ( .A(round_inst_srout2_y[58]), .B(
        round_inst_srout2_y[43]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[58]) );
  MUX2_X1 round_inst_mux_inv_y2_U46 ( .A(round_inst_srout2_y[42]), .B(
        round_inst_srout2_y[27]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[42]) );
  MUX2_X1 round_inst_mux_inv_y2_U45 ( .A(round_inst_srout2_y[46]), .B(
        round_inst_srout2_y[47]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[46]) );
  MUX2_X1 round_inst_mux_inv_y2_U44 ( .A(round_inst_srout2_y[22]), .B(
        round_inst_srout2_y[55]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[22]) );
  MUX2_X1 round_inst_mux_inv_y2_U43 ( .A(round_inst_srout2_y[30]), .B(
        round_inst_srout2_y[31]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[30]) );
  MUX2_X1 round_inst_mux_inv_y2_U42 ( .A(round_inst_srout2_y[6]), .B(
        round_inst_srout2_y[39]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[6]) );
  MUX2_X1 round_inst_mux_inv_y2_U41 ( .A(round_inst_srout2_y[55]), .B(
        round_inst_srout2_y[22]), .S(round_inst_mux_inv_y2_n266), .Z(
        round_inst_min_y[55]) );
  INV_X1 round_inst_mux_inv_y2_U40 ( .A(round_inst_mux_inv_y2_n263), .ZN(
        round_inst_mux_inv_y2_n266) );
  MUX2_X1 round_inst_mux_inv_y2_U39 ( .A(round_inst_srout2_y[35]), .B(
        round_inst_srout2_y[50]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[35]) );
  MUX2_X1 round_inst_mux_inv_y2_U38 ( .A(round_inst_srout2_y[11]), .B(
        round_inst_srout2_y[58]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[11]) );
  MUX2_X1 round_inst_mux_inv_y2_U37 ( .A(round_inst_srout2_y[16]), .B(
        round_inst_sout_y[16]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[16]) );
  MUX2_X1 round_inst_mux_inv_y2_U36 ( .A(round_inst_srout2_y[52]), .B(
        round_inst_sout_y[52]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[52]) );
  MUX2_X1 round_inst_mux_inv_y2_U35 ( .A(round_inst_srout2_y[48]), .B(
        round_inst_sout_y[48]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[48]) );
  MUX2_X1 round_inst_mux_inv_y2_U34 ( .A(round_inst_srout2_y[40]), .B(
        round_inst_sout_y[40]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[40]) );
  MUX2_X1 round_inst_mux_inv_y2_U33 ( .A(round_inst_srout2_y[32]), .B(
        round_inst_sout_y[32]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[32]) );
  MUX2_X1 round_inst_mux_inv_y2_U32 ( .A(round_inst_srout2_y[20]), .B(
        round_inst_sout_y[20]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[20]) );
  MUX2_X1 round_inst_mux_inv_y2_U31 ( .A(round_inst_srout2_y[12]), .B(
        round_inst_sout_y[12]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[12]) );
  MUX2_X1 round_inst_mux_inv_y2_U30 ( .A(round_inst_srout2_y[0]), .B(
        round_inst_sout_y[0]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[0]) );
  MUX2_X1 round_inst_mux_inv_y2_U29 ( .A(round_inst_srout2_y[59]), .B(
        round_inst_srout2_y[42]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[59]) );
  MUX2_X1 round_inst_mux_inv_y2_U28 ( .A(round_inst_srout2_y[63]), .B(
        round_inst_srout2_y[62]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[63]) );
  MUX2_X1 round_inst_mux_inv_y2_U27 ( .A(round_inst_srout2_y[43]), .B(
        round_inst_srout2_y[26]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[43]) );
  MUX2_X1 round_inst_mux_inv_y2_U26 ( .A(round_inst_srout2_y[47]), .B(
        round_inst_srout2_y[46]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[47]) );
  MUX2_X1 round_inst_mux_inv_y2_U25 ( .A(round_inst_srout2_y[27]), .B(
        round_inst_srout2_y[10]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[27]) );
  MUX2_X1 round_inst_mux_inv_y2_U24 ( .A(round_inst_srout2_y[31]), .B(
        round_inst_srout2_y[30]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[31]) );
  MUX2_X1 round_inst_mux_inv_y2_U23 ( .A(round_inst_srout2_y[7]), .B(
        round_inst_srout2_y[38]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[7]) );
  MUX2_X1 round_inst_mux_inv_y2_U22 ( .A(round_inst_srout2_y[60]), .B(
        round_inst_sout_y[60]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[60]) );
  MUX2_X1 round_inst_mux_inv_y2_U21 ( .A(round_inst_srout2_y[56]), .B(
        round_inst_sout_y[56]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[56]) );
  MUX2_X1 round_inst_mux_inv_y2_U20 ( .A(round_inst_srout2_y[44]), .B(
        round_inst_sout_y[44]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[44]) );
  MUX2_X1 round_inst_mux_inv_y2_U19 ( .A(round_inst_srout2_y[36]), .B(
        round_inst_sout_y[36]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[36]) );
  MUX2_X1 round_inst_mux_inv_y2_U18 ( .A(round_inst_srout2_y[28]), .B(
        round_inst_sout_y[28]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[28]) );
  MUX2_X1 round_inst_mux_inv_y2_U17 ( .A(round_inst_srout2_y[24]), .B(
        round_inst_sout_y[24]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[24]) );
  MUX2_X1 round_inst_mux_inv_y2_U16 ( .A(round_inst_srout2_y[8]), .B(
        round_inst_sout_y[8]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[8]) );
  MUX2_X1 round_inst_mux_inv_y2_U15 ( .A(round_inst_srout2_y[4]), .B(
        round_inst_sout_y[4]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[4]) );
  MUX2_X1 round_inst_mux_inv_y2_U14 ( .A(round_inst_srout2_y[51]), .B(
        round_inst_srout2_y[2]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[51]) );
  MUX2_X1 round_inst_mux_inv_y2_U13 ( .A(round_inst_srout2_y[39]), .B(
        round_inst_srout2_y[6]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[39]) );
  MUX2_X1 round_inst_mux_inv_y2_U12 ( .A(round_inst_srout2_y[23]), .B(
        round_inst_srout2_y[54]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[23]) );
  MUX2_X1 round_inst_mux_inv_y2_U11 ( .A(round_inst_srout2_y[15]), .B(
        round_inst_srout2_y[14]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[15]) );
  MUX2_X1 round_inst_mux_inv_y2_U10 ( .A(round_inst_srout2_y[37]), .B(
        round_inst_srout2_y[4]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[37]) );
  MUX2_X1 round_inst_mux_inv_y2_U9 ( .A(round_inst_srout2_y[13]), .B(
        round_inst_srout2_y[12]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[13]) );
  MUX2_X1 round_inst_mux_inv_y2_U8 ( .A(round_inst_srout2_y[61]), .B(
        round_inst_srout2_y[60]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[61]) );
  MUX2_X1 round_inst_mux_inv_y2_U7 ( .A(round_inst_srout2_y[53]), .B(
        round_inst_srout2_y[20]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[53]) );
  MUX2_X1 round_inst_mux_inv_y2_U6 ( .A(round_inst_srout2_y[41]), .B(
        round_inst_srout2_y[24]), .S(round_inst_mux_inv_y2_n264), .Z(
        round_inst_min_y[41]) );
  INV_X1 round_inst_mux_inv_y2_U5 ( .A(round_inst_mux_inv_y2_n263), .ZN(
        round_inst_mux_inv_y2_n264) );
  MUX2_X1 round_inst_mux_inv_y2_U4 ( .A(round_inst_srout2_y[21]), .B(
        round_inst_srout2_y[52]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[21]) );
  MUX2_X1 round_inst_mux_inv_y2_U3 ( .A(round_inst_srout2_y[9]), .B(
        round_inst_srout2_y[56]), .S(round_inst_mux_inv_y2_n265), .Z(
        round_inst_min_y[9]) );
  INV_X1 round_inst_mux_inv_y2_U2 ( .A(round_inst_mux_inv_y2_n263), .ZN(
        round_inst_mux_inv_y2_n265) );
  INV_X1 round_inst_mux_inv_y2_U1 ( .A(inv_sig), .ZN(
        round_inst_mux_inv_y2_n263) );
  MUX2_X1 round_inst_mux_inv_z2_U69 ( .A(round_inst_srout2_z[1]), .B(
        round_inst_srout2_z[16]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[1]) );
  MUX2_X1 round_inst_mux_inv_z2_U68 ( .A(round_inst_srout2_z[2]), .B(
        round_inst_srout2_z[19]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[2]) );
  MUX2_X1 round_inst_mux_inv_z2_U67 ( .A(round_inst_srout2_z[19]), .B(
        round_inst_srout2_z[34]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[19]) );
  MUX2_X1 round_inst_mux_inv_z2_U66 ( .A(round_inst_srout2_z[16]), .B(
        round_inst_sout_z[16]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[16]) );
  MUX2_X1 round_inst_mux_inv_z2_U65 ( .A(round_inst_srout2_z[57]), .B(
        round_inst_srout2_z[40]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[57]) );
  MUX2_X1 round_inst_mux_inv_z2_U64 ( .A(round_inst_srout2_z[49]), .B(
        round_inst_srout2_z[0]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[49]) );
  MUX2_X1 round_inst_mux_inv_z2_U63 ( .A(round_inst_srout2_z[37]), .B(
        round_inst_srout2_z[4]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[37]) );
  MUX2_X1 round_inst_mux_inv_z2_U62 ( .A(round_inst_srout2_z[33]), .B(
        round_inst_srout2_z[48]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[33]) );
  MUX2_X1 round_inst_mux_inv_z2_U61 ( .A(round_inst_srout2_z[17]), .B(
        round_inst_srout2_z[32]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[17]) );
  MUX2_X1 round_inst_mux_inv_z2_U60 ( .A(round_inst_srout2_z[25]), .B(
        round_inst_srout2_z[8]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[25]) );
  MUX2_X1 round_inst_mux_inv_z2_U59 ( .A(round_inst_srout2_z[13]), .B(
        round_inst_srout2_z[12]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[13]) );
  MUX2_X1 round_inst_mux_inv_z2_U58 ( .A(round_inst_srout2_z[61]), .B(
        round_inst_srout2_z[60]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[61]) );
  MUX2_X1 round_inst_mux_inv_z2_U57 ( .A(round_inst_srout2_z[53]), .B(
        round_inst_srout2_z[20]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[53]) );
  MUX2_X1 round_inst_mux_inv_z2_U56 ( .A(round_inst_srout2_z[45]), .B(
        round_inst_srout2_z[44]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[45]) );
  MUX2_X1 round_inst_mux_inv_z2_U55 ( .A(round_inst_srout2_z[41]), .B(
        round_inst_srout2_z[24]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[41]) );
  MUX2_X1 round_inst_mux_inv_z2_U54 ( .A(round_inst_srout2_z[21]), .B(
        round_inst_srout2_z[52]), .S(round_inst_mux_inv_z2_n266), .Z(
        round_inst_min_z[21]) );
  INV_X1 round_inst_mux_inv_z2_U53 ( .A(round_inst_mux_inv_z2_n265), .ZN(
        round_inst_mux_inv_z2_n266) );
  MUX2_X1 round_inst_mux_inv_z2_U52 ( .A(round_inst_srout2_z[29]), .B(
        round_inst_srout2_z[28]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[29]) );
  MUX2_X1 round_inst_mux_inv_z2_U51 ( .A(round_inst_srout2_z[9]), .B(
        round_inst_srout2_z[56]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[9]) );
  MUX2_X1 round_inst_mux_inv_z2_U50 ( .A(round_inst_srout2_z[5]), .B(
        round_inst_srout2_z[36]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[5]) );
  MUX2_X1 round_inst_mux_inv_z2_U49 ( .A(round_inst_srout2_z[50]), .B(
        round_inst_srout2_z[3]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[50]) );
  MUX2_X1 round_inst_mux_inv_z2_U48 ( .A(round_inst_srout2_z[54]), .B(
        round_inst_srout2_z[23]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[54]) );
  MUX2_X1 round_inst_mux_inv_z2_U47 ( .A(round_inst_srout2_z[34]), .B(
        round_inst_srout2_z[51]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[34]) );
  MUX2_X1 round_inst_mux_inv_z2_U46 ( .A(round_inst_srout2_z[38]), .B(
        round_inst_srout2_z[7]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[38]) );
  MUX2_X1 round_inst_mux_inv_z2_U45 ( .A(round_inst_srout2_z[18]), .B(
        round_inst_srout2_z[35]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[18]) );
  MUX2_X1 round_inst_mux_inv_z2_U44 ( .A(round_inst_srout2_z[26]), .B(
        round_inst_srout2_z[11]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[26]) );
  MUX2_X1 round_inst_mux_inv_z2_U43 ( .A(round_inst_srout2_z[14]), .B(
        round_inst_srout2_z[15]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[14]) );
  MUX2_X1 round_inst_mux_inv_z2_U42 ( .A(round_inst_srout2_z[10]), .B(
        round_inst_srout2_z[59]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[10]) );
  MUX2_X1 round_inst_mux_inv_z2_U41 ( .A(round_inst_srout2_z[62]), .B(
        round_inst_srout2_z[63]), .S(round_inst_mux_inv_z2_n267), .Z(
        round_inst_min_z[62]) );
  INV_X1 round_inst_mux_inv_z2_U40 ( .A(round_inst_mux_inv_z2_n265), .ZN(
        round_inst_mux_inv_z2_n267) );
  INV_X1 round_inst_mux_inv_z2_U39 ( .A(inv_sig), .ZN(
        round_inst_mux_inv_z2_n265) );
  MUX2_X1 round_inst_mux_inv_z2_U38 ( .A(round_inst_srout2_z[58]), .B(
        round_inst_srout2_z[43]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[58]) );
  MUX2_X1 round_inst_mux_inv_z2_U37 ( .A(round_inst_srout2_z[42]), .B(
        round_inst_srout2_z[27]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[42]) );
  MUX2_X1 round_inst_mux_inv_z2_U36 ( .A(round_inst_srout2_z[22]), .B(
        round_inst_srout2_z[55]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[22]) );
  MUX2_X1 round_inst_mux_inv_z2_U35 ( .A(round_inst_srout2_z[30]), .B(
        round_inst_srout2_z[31]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[30]) );
  MUX2_X1 round_inst_mux_inv_z2_U34 ( .A(round_inst_srout2_z[6]), .B(
        round_inst_srout2_z[39]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[6]) );
  MUX2_X1 round_inst_mux_inv_z2_U33 ( .A(round_inst_srout2_z[55]), .B(
        round_inst_srout2_z[22]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[55]) );
  MUX2_X1 round_inst_mux_inv_z2_U32 ( .A(round_inst_srout2_z[51]), .B(
        round_inst_srout2_z[2]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[51]) );
  MUX2_X1 round_inst_mux_inv_z2_U31 ( .A(round_inst_srout2_z[39]), .B(
        round_inst_srout2_z[6]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[39]) );
  MUX2_X1 round_inst_mux_inv_z2_U30 ( .A(round_inst_srout2_z[35]), .B(
        round_inst_srout2_z[50]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[35]) );
  MUX2_X1 round_inst_mux_inv_z2_U29 ( .A(round_inst_srout2_z[23]), .B(
        round_inst_srout2_z[54]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[23]) );
  MUX2_X1 round_inst_mux_inv_z2_U28 ( .A(round_inst_srout2_z[11]), .B(
        round_inst_srout2_z[58]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[11]) );
  MUX2_X1 round_inst_mux_inv_z2_U27 ( .A(round_inst_srout2_z[15]), .B(
        round_inst_srout2_z[14]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[15]) );
  MUX2_X1 round_inst_mux_inv_z2_U26 ( .A(round_inst_srout2_z[52]), .B(
        round_inst_sout_z[52]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[52]) );
  MUX2_X1 round_inst_mux_inv_z2_U25 ( .A(round_inst_srout2_z[48]), .B(
        round_inst_sout_z[48]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[48]) );
  MUX2_X1 round_inst_mux_inv_z2_U24 ( .A(round_inst_srout2_z[40]), .B(
        round_inst_sout_z[40]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[40]) );
  MUX2_X1 round_inst_mux_inv_z2_U23 ( .A(round_inst_srout2_z[32]), .B(
        round_inst_sout_z[32]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[32]) );
  MUX2_X1 round_inst_mux_inv_z2_U22 ( .A(round_inst_srout2_z[20]), .B(
        round_inst_sout_z[20]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[20]) );
  MUX2_X1 round_inst_mux_inv_z2_U21 ( .A(round_inst_srout2_z[12]), .B(
        round_inst_sout_z[12]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[12]) );
  MUX2_X1 round_inst_mux_inv_z2_U20 ( .A(round_inst_srout2_z[0]), .B(
        round_inst_sout_z[0]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[0]) );
  MUX2_X1 round_inst_mux_inv_z2_U19 ( .A(round_inst_srout2_z[59]), .B(
        round_inst_srout2_z[42]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[59]) );
  MUX2_X1 round_inst_mux_inv_z2_U18 ( .A(round_inst_srout2_z[63]), .B(
        round_inst_srout2_z[62]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[63]) );
  MUX2_X1 round_inst_mux_inv_z2_U17 ( .A(round_inst_srout2_z[43]), .B(
        round_inst_srout2_z[26]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[43]) );
  MUX2_X1 round_inst_mux_inv_z2_U16 ( .A(round_inst_srout2_z[47]), .B(
        round_inst_srout2_z[46]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[47]) );
  MUX2_X1 round_inst_mux_inv_z2_U15 ( .A(round_inst_srout2_z[27]), .B(
        round_inst_srout2_z[10]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[27]) );
  MUX2_X1 round_inst_mux_inv_z2_U14 ( .A(round_inst_srout2_z[31]), .B(
        round_inst_srout2_z[30]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[31]) );
  MUX2_X1 round_inst_mux_inv_z2_U13 ( .A(round_inst_srout2_z[7]), .B(
        round_inst_srout2_z[38]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[7]) );
  MUX2_X1 round_inst_mux_inv_z2_U12 ( .A(round_inst_srout2_z[3]), .B(
        round_inst_srout2_z[18]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[3]) );
  MUX2_X1 round_inst_mux_inv_z2_U11 ( .A(round_inst_srout2_z[60]), .B(
        round_inst_sout_z[60]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[60]) );
  MUX2_X1 round_inst_mux_inv_z2_U10 ( .A(round_inst_srout2_z[56]), .B(
        round_inst_sout_z[56]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[56]) );
  MUX2_X1 round_inst_mux_inv_z2_U9 ( .A(round_inst_srout2_z[44]), .B(
        round_inst_sout_z[44]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[44]) );
  MUX2_X1 round_inst_mux_inv_z2_U8 ( .A(round_inst_srout2_z[36]), .B(
        round_inst_sout_z[36]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[36]) );
  MUX2_X1 round_inst_mux_inv_z2_U7 ( .A(round_inst_srout2_z[28]), .B(
        round_inst_sout_z[28]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[28]) );
  MUX2_X1 round_inst_mux_inv_z2_U6 ( .A(round_inst_srout2_z[24]), .B(
        round_inst_sout_z[24]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[24]) );
  MUX2_X1 round_inst_mux_inv_z2_U5 ( .A(round_inst_srout2_z[8]), .B(
        round_inst_sout_z[8]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[8]) );
  MUX2_X1 round_inst_mux_inv_z2_U4 ( .A(round_inst_srout2_z[4]), .B(
        round_inst_sout_z[4]), .S(round_inst_mux_inv_z2_n263), .Z(
        round_inst_min_z[4]) );
  INV_X1 round_inst_mux_inv_z2_U3 ( .A(round_inst_mux_inv_z2_n265), .ZN(
        round_inst_mux_inv_z2_n263) );
  MUX2_X1 round_inst_mux_inv_z2_U2 ( .A(round_inst_srout2_z[46]), .B(
        round_inst_srout2_z[47]), .S(round_inst_mux_inv_z2_n264), .Z(
        round_inst_min_z[46]) );
  INV_X1 round_inst_mux_inv_z2_U1 ( .A(round_inst_mux_inv_z2_n265), .ZN(
        round_inst_mux_inv_z2_n264) );
  XNOR2_X1 round_inst_mw_inst_U96 ( .A(round_inst_min_w[59]), .B(
        round_inst_mw_inst_n32), .ZN(rout_w[63]) );
  XNOR2_X1 round_inst_mw_inst_U95 ( .A(round_inst_min_w[63]), .B(
        round_inst_mw_inst_n32), .ZN(rout_w[51]) );
  XNOR2_X1 round_inst_mw_inst_U94 ( .A(round_inst_min_w[51]), .B(
        round_inst_min_w[55]), .ZN(round_inst_mw_inst_n32) );
  XNOR2_X1 round_inst_mw_inst_U93 ( .A(round_inst_min_w[62]), .B(
        round_inst_mw_inst_n31), .ZN(rout_w[62]) );
  XNOR2_X1 round_inst_mw_inst_U92 ( .A(round_inst_min_w[58]), .B(
        round_inst_mw_inst_n31), .ZN(rout_w[58]) );
  XNOR2_X1 round_inst_mw_inst_U91 ( .A(round_inst_min_w[50]), .B(
        round_inst_min_w[54]), .ZN(round_inst_mw_inst_n31) );
  XNOR2_X1 round_inst_mw_inst_U90 ( .A(round_inst_min_w[60]), .B(
        round_inst_mw_inst_n30), .ZN(rout_w[60]) );
  XNOR2_X1 round_inst_mw_inst_U89 ( .A(round_inst_min_w[48]), .B(
        round_inst_mw_inst_n30), .ZN(rout_w[48]) );
  XNOR2_X1 round_inst_mw_inst_U88 ( .A(round_inst_min_w[52]), .B(
        round_inst_min_w[56]), .ZN(round_inst_mw_inst_n30) );
  XNOR2_X1 round_inst_mw_inst_U87 ( .A(round_inst_min_w[42]), .B(
        round_inst_mw_inst_n29), .ZN(rout_w[46]) );
  XNOR2_X1 round_inst_mw_inst_U86 ( .A(round_inst_min_w[46]), .B(
        round_inst_mw_inst_n29), .ZN(rout_w[34]) );
  XNOR2_X1 round_inst_mw_inst_U85 ( .A(round_inst_min_w[34]), .B(
        round_inst_min_w[38]), .ZN(round_inst_mw_inst_n29) );
  XNOR2_X1 round_inst_mw_inst_U84 ( .A(round_inst_min_w[28]), .B(
        round_inst_mw_inst_n28), .ZN(rout_w[28]) );
  XNOR2_X1 round_inst_mw_inst_U83 ( .A(round_inst_min_w[20]), .B(
        round_inst_mw_inst_n28), .ZN(rout_w[20]) );
  XNOR2_X1 round_inst_mw_inst_U82 ( .A(round_inst_min_w[24]), .B(
        round_inst_min_w[16]), .ZN(round_inst_mw_inst_n28) );
  XNOR2_X1 round_inst_mw_inst_U81 ( .A(round_inst_min_w[31]), .B(
        round_inst_mw_inst_n27), .ZN(rout_w[27]) );
  XNOR2_X1 round_inst_mw_inst_U80 ( .A(round_inst_min_w[23]), .B(
        round_inst_mw_inst_n27), .ZN(rout_w[19]) );
  XNOR2_X1 round_inst_mw_inst_U79 ( .A(round_inst_min_w[19]), .B(
        round_inst_min_w[27]), .ZN(round_inst_mw_inst_n27) );
  XNOR2_X1 round_inst_mw_inst_U78 ( .A(round_inst_min_w[45]), .B(
        round_inst_mw_inst_n26), .ZN(rout_w[45]) );
  XNOR2_X1 round_inst_mw_inst_U77 ( .A(round_inst_min_w[41]), .B(
        round_inst_mw_inst_n26), .ZN(rout_w[41]) );
  XNOR2_X1 round_inst_mw_inst_U76 ( .A(round_inst_min_w[33]), .B(
        round_inst_min_w[37]), .ZN(round_inst_mw_inst_n26) );
  XNOR2_X1 round_inst_mw_inst_U75 ( .A(round_inst_min_w[22]), .B(
        round_inst_mw_inst_n25), .ZN(rout_w[26]) );
  XNOR2_X1 round_inst_mw_inst_U74 ( .A(round_inst_min_w[18]), .B(
        round_inst_mw_inst_n25), .ZN(rout_w[22]) );
  XNOR2_X1 round_inst_mw_inst_U73 ( .A(round_inst_min_w[30]), .B(
        round_inst_min_w[26]), .ZN(round_inst_mw_inst_n25) );
  XNOR2_X1 round_inst_mw_inst_U72 ( .A(round_inst_min_w[16]), .B(
        round_inst_mw_inst_n24), .ZN(rout_w[24]) );
  XNOR2_X1 round_inst_mw_inst_U71 ( .A(round_inst_min_w[24]), .B(
        round_inst_mw_inst_n24), .ZN(rout_w[16]) );
  XNOR2_X1 round_inst_mw_inst_U70 ( .A(round_inst_min_w[28]), .B(
        round_inst_min_w[20]), .ZN(round_inst_mw_inst_n24) );
  XNOR2_X1 round_inst_mw_inst_U69 ( .A(round_inst_min_w[55]), .B(
        round_inst_mw_inst_n23), .ZN(rout_w[59]) );
  XNOR2_X1 round_inst_mw_inst_U68 ( .A(round_inst_min_w[51]), .B(
        round_inst_mw_inst_n23), .ZN(rout_w[55]) );
  XNOR2_X1 round_inst_mw_inst_U67 ( .A(round_inst_min_w[59]), .B(
        round_inst_min_w[63]), .ZN(round_inst_mw_inst_n23) );
  XNOR2_X1 round_inst_mw_inst_U66 ( .A(round_inst_min_w[21]), .B(
        round_inst_mw_inst_n22), .ZN(rout_w[21]) );
  XNOR2_X1 round_inst_mw_inst_U65 ( .A(round_inst_min_w[17]), .B(
        round_inst_mw_inst_n22), .ZN(rout_w[17]) );
  XNOR2_X1 round_inst_mw_inst_U64 ( .A(round_inst_min_w[25]), .B(
        round_inst_min_w[29]), .ZN(round_inst_mw_inst_n22) );
  XNOR2_X1 round_inst_mw_inst_U63 ( .A(round_inst_min_w[7]), .B(
        round_inst_mw_inst_n21), .ZN(rout_w[15]) );
  XNOR2_X1 round_inst_mw_inst_U62 ( .A(round_inst_min_w[15]), .B(
        round_inst_mw_inst_n21), .ZN(rout_w[7]) );
  XNOR2_X1 round_inst_mw_inst_U61 ( .A(round_inst_min_w[3]), .B(
        round_inst_min_w[11]), .ZN(round_inst_mw_inst_n21) );
  XNOR2_X1 round_inst_mw_inst_U60 ( .A(round_inst_min_w[44]), .B(
        round_inst_mw_inst_n20), .ZN(rout_w[44]) );
  XNOR2_X1 round_inst_mw_inst_U59 ( .A(round_inst_min_w[36]), .B(
        round_inst_mw_inst_n20), .ZN(rout_w[36]) );
  XNOR2_X1 round_inst_mw_inst_U58 ( .A(round_inst_min_w[40]), .B(
        round_inst_min_w[32]), .ZN(round_inst_mw_inst_n20) );
  XNOR2_X1 round_inst_mw_inst_U57 ( .A(round_inst_min_w[11]), .B(
        round_inst_mw_inst_n19), .ZN(rout_w[11]) );
  XNOR2_X1 round_inst_mw_inst_U56 ( .A(round_inst_min_w[3]), .B(
        round_inst_mw_inst_n19), .ZN(rout_w[3]) );
  XNOR2_X1 round_inst_mw_inst_U55 ( .A(round_inst_min_w[7]), .B(
        round_inst_min_w[15]), .ZN(round_inst_mw_inst_n19) );
  XNOR2_X1 round_inst_mw_inst_U54 ( .A(round_inst_min_w[6]), .B(
        round_inst_mw_inst_n18), .ZN(rout_w[14]) );
  XNOR2_X1 round_inst_mw_inst_U53 ( .A(round_inst_min_w[10]), .B(
        round_inst_mw_inst_n18), .ZN(rout_w[2]) );
  XNOR2_X1 round_inst_mw_inst_U52 ( .A(round_inst_min_w[14]), .B(
        round_inst_min_w[2]), .ZN(round_inst_mw_inst_n18) );
  XNOR2_X1 round_inst_mw_inst_U51 ( .A(round_inst_min_w[61]), .B(
        round_inst_mw_inst_n17), .ZN(rout_w[61]) );
  XNOR2_X1 round_inst_mw_inst_U50 ( .A(round_inst_min_w[53]), .B(
        round_inst_mw_inst_n17), .ZN(rout_w[53]) );
  XNOR2_X1 round_inst_mw_inst_U49 ( .A(round_inst_min_w[57]), .B(
        round_inst_min_w[49]), .ZN(round_inst_mw_inst_n17) );
  XNOR2_X1 round_inst_mw_inst_U48 ( .A(round_inst_min_w[49]), .B(
        round_inst_mw_inst_n16), .ZN(rout_w[57]) );
  XNOR2_X1 round_inst_mw_inst_U47 ( .A(round_inst_min_w[57]), .B(
        round_inst_mw_inst_n16), .ZN(rout_w[49]) );
  XNOR2_X1 round_inst_mw_inst_U46 ( .A(round_inst_min_w[61]), .B(
        round_inst_min_w[53]), .ZN(round_inst_mw_inst_n16) );
  XNOR2_X1 round_inst_mw_inst_U45 ( .A(round_inst_min_w[2]), .B(
        round_inst_mw_inst_n15), .ZN(rout_w[10]) );
  XNOR2_X1 round_inst_mw_inst_U44 ( .A(round_inst_min_w[14]), .B(
        round_inst_mw_inst_n15), .ZN(rout_w[6]) );
  XNOR2_X1 round_inst_mw_inst_U43 ( .A(round_inst_min_w[6]), .B(
        round_inst_min_w[10]), .ZN(round_inst_mw_inst_n15) );
  XNOR2_X1 round_inst_mw_inst_U42 ( .A(round_inst_min_w[9]), .B(
        round_inst_mw_inst_n14), .ZN(rout_w[13]) );
  XNOR2_X1 round_inst_mw_inst_U41 ( .A(round_inst_min_w[5]), .B(
        round_inst_mw_inst_n14), .ZN(rout_w[9]) );
  XNOR2_X1 round_inst_mw_inst_U40 ( .A(round_inst_min_w[13]), .B(
        round_inst_min_w[1]), .ZN(round_inst_mw_inst_n14) );
  XNOR2_X1 round_inst_mw_inst_U39 ( .A(round_inst_min_w[47]), .B(
        round_inst_mw_inst_n13), .ZN(rout_w[43]) );
  XNOR2_X1 round_inst_mw_inst_U38 ( .A(round_inst_min_w[39]), .B(
        round_inst_mw_inst_n13), .ZN(rout_w[35]) );
  XNOR2_X1 round_inst_mw_inst_U37 ( .A(round_inst_min_w[35]), .B(
        round_inst_min_w[43]), .ZN(round_inst_mw_inst_n13) );
  XNOR2_X1 round_inst_mw_inst_U36 ( .A(round_inst_min_w[8]), .B(
        round_inst_mw_inst_n12), .ZN(rout_w[12]) );
  XNOR2_X1 round_inst_mw_inst_U35 ( .A(round_inst_min_w[0]), .B(
        round_inst_mw_inst_n12), .ZN(rout_w[4]) );
  XNOR2_X1 round_inst_mw_inst_U34 ( .A(round_inst_min_w[4]), .B(
        round_inst_min_w[12]), .ZN(round_inst_mw_inst_n12) );
  XNOR2_X1 round_inst_mw_inst_U33 ( .A(round_inst_min_w[56]), .B(
        round_inst_mw_inst_n11), .ZN(rout_w[56]) );
  XNOR2_X1 round_inst_mw_inst_U32 ( .A(round_inst_min_w[52]), .B(
        round_inst_mw_inst_n11), .ZN(rout_w[52]) );
  XNOR2_X1 round_inst_mw_inst_U31 ( .A(round_inst_min_w[60]), .B(
        round_inst_min_w[48]), .ZN(round_inst_mw_inst_n11) );
  XNOR2_X1 round_inst_mw_inst_U30 ( .A(round_inst_min_w[38]), .B(
        round_inst_mw_inst_n10), .ZN(rout_w[42]) );
  XNOR2_X1 round_inst_mw_inst_U29 ( .A(round_inst_min_w[34]), .B(
        round_inst_mw_inst_n10), .ZN(rout_w[38]) );
  XNOR2_X1 round_inst_mw_inst_U28 ( .A(round_inst_min_w[42]), .B(
        round_inst_min_w[46]), .ZN(round_inst_mw_inst_n10) );
  XNOR2_X1 round_inst_mw_inst_U27 ( .A(round_inst_min_w[32]), .B(
        round_inst_mw_inst_n9), .ZN(rout_w[40]) );
  XNOR2_X1 round_inst_mw_inst_U26 ( .A(round_inst_min_w[40]), .B(
        round_inst_mw_inst_n9), .ZN(rout_w[32]) );
  XNOR2_X1 round_inst_mw_inst_U25 ( .A(round_inst_min_w[44]), .B(
        round_inst_min_w[36]), .ZN(round_inst_mw_inst_n9) );
  XNOR2_X1 round_inst_mw_inst_U24 ( .A(round_inst_min_w[1]), .B(
        round_inst_mw_inst_n8), .ZN(rout_w[5]) );
  XNOR2_X1 round_inst_mw_inst_U23 ( .A(round_inst_min_w[13]), .B(
        round_inst_mw_inst_n8), .ZN(rout_w[1]) );
  XNOR2_X1 round_inst_mw_inst_U22 ( .A(round_inst_min_w[9]), .B(
        round_inst_min_w[5]), .ZN(round_inst_mw_inst_n8) );
  XNOR2_X1 round_inst_mw_inst_U21 ( .A(round_inst_min_w[12]), .B(
        round_inst_mw_inst_n7), .ZN(rout_w[8]) );
  XNOR2_X1 round_inst_mw_inst_U20 ( .A(round_inst_min_w[4]), .B(
        round_inst_mw_inst_n7), .ZN(rout_w[0]) );
  XNOR2_X1 round_inst_mw_inst_U19 ( .A(round_inst_min_w[8]), .B(
        round_inst_min_w[0]), .ZN(round_inst_mw_inst_n7) );
  XNOR2_X1 round_inst_mw_inst_U18 ( .A(round_inst_min_w[54]), .B(
        round_inst_mw_inst_n6), .ZN(rout_w[54]) );
  XNOR2_X1 round_inst_mw_inst_U17 ( .A(round_inst_min_w[50]), .B(
        round_inst_mw_inst_n6), .ZN(rout_w[50]) );
  XNOR2_X1 round_inst_mw_inst_U16 ( .A(round_inst_min_w[62]), .B(
        round_inst_min_w[58]), .ZN(round_inst_mw_inst_n6) );
  XNOR2_X1 round_inst_mw_inst_U15 ( .A(round_inst_min_w[37]), .B(
        round_inst_mw_inst_n5), .ZN(rout_w[37]) );
  XNOR2_X1 round_inst_mw_inst_U14 ( .A(round_inst_min_w[33]), .B(
        round_inst_mw_inst_n5), .ZN(rout_w[33]) );
  XNOR2_X1 round_inst_mw_inst_U13 ( .A(round_inst_min_w[45]), .B(
        round_inst_min_w[41]), .ZN(round_inst_mw_inst_n5) );
  XNOR2_X1 round_inst_mw_inst_U12 ( .A(round_inst_min_w[27]), .B(
        round_inst_mw_inst_n4), .ZN(rout_w[31]) );
  XNOR2_X1 round_inst_mw_inst_U11 ( .A(round_inst_min_w[19]), .B(
        round_inst_mw_inst_n4), .ZN(rout_w[23]) );
  XNOR2_X1 round_inst_mw_inst_U10 ( .A(round_inst_min_w[31]), .B(
        round_inst_min_w[23]), .ZN(round_inst_mw_inst_n4) );
  XNOR2_X1 round_inst_mw_inst_U9 ( .A(round_inst_min_w[43]), .B(
        round_inst_mw_inst_n3), .ZN(rout_w[47]) );
  XNOR2_X1 round_inst_mw_inst_U8 ( .A(round_inst_min_w[35]), .B(
        round_inst_mw_inst_n3), .ZN(rout_w[39]) );
  XNOR2_X1 round_inst_mw_inst_U7 ( .A(round_inst_min_w[47]), .B(
        round_inst_min_w[39]), .ZN(round_inst_mw_inst_n3) );
  XNOR2_X1 round_inst_mw_inst_U6 ( .A(round_inst_min_w[26]), .B(
        round_inst_mw_inst_n2), .ZN(rout_w[30]) );
  XNOR2_X1 round_inst_mw_inst_U5 ( .A(round_inst_min_w[30]), .B(
        round_inst_mw_inst_n2), .ZN(rout_w[18]) );
  XNOR2_X1 round_inst_mw_inst_U4 ( .A(round_inst_min_w[22]), .B(
        round_inst_min_w[18]), .ZN(round_inst_mw_inst_n2) );
  XNOR2_X1 round_inst_mw_inst_U3 ( .A(round_inst_min_w[29]), .B(
        round_inst_mw_inst_n1), .ZN(rout_w[29]) );
  XNOR2_X1 round_inst_mw_inst_U2 ( .A(round_inst_min_w[25]), .B(
        round_inst_mw_inst_n1), .ZN(rout_w[25]) );
  XNOR2_X1 round_inst_mw_inst_U1 ( .A(round_inst_min_w[21]), .B(
        round_inst_min_w[17]), .ZN(round_inst_mw_inst_n1) );
  XNOR2_X1 round_inst_mx_inst_U96 ( .A(round_inst_min_x[59]), .B(
        round_inst_mx_inst_n96), .ZN(rout_x[63]) );
  XNOR2_X1 round_inst_mx_inst_U95 ( .A(round_inst_min_x[63]), .B(
        round_inst_mx_inst_n96), .ZN(rout_x[51]) );
  XNOR2_X1 round_inst_mx_inst_U94 ( .A(round_inst_min_x[51]), .B(
        round_inst_min_x[55]), .ZN(round_inst_mx_inst_n96) );
  XNOR2_X1 round_inst_mx_inst_U93 ( .A(round_inst_min_x[62]), .B(
        round_inst_mx_inst_n95), .ZN(rout_x[62]) );
  XNOR2_X1 round_inst_mx_inst_U92 ( .A(round_inst_min_x[58]), .B(
        round_inst_mx_inst_n95), .ZN(rout_x[58]) );
  XNOR2_X1 round_inst_mx_inst_U91 ( .A(round_inst_min_x[50]), .B(
        round_inst_min_x[54]), .ZN(round_inst_mx_inst_n95) );
  XNOR2_X1 round_inst_mx_inst_U90 ( .A(round_inst_min_x[60]), .B(
        round_inst_mx_inst_n94), .ZN(rout_x[60]) );
  XNOR2_X1 round_inst_mx_inst_U89 ( .A(round_inst_min_x[48]), .B(
        round_inst_mx_inst_n94), .ZN(rout_x[48]) );
  XNOR2_X1 round_inst_mx_inst_U88 ( .A(round_inst_min_x[52]), .B(
        round_inst_min_x[56]), .ZN(round_inst_mx_inst_n94) );
  XNOR2_X1 round_inst_mx_inst_U87 ( .A(round_inst_min_x[42]), .B(
        round_inst_mx_inst_n93), .ZN(rout_x[46]) );
  XNOR2_X1 round_inst_mx_inst_U86 ( .A(round_inst_min_x[46]), .B(
        round_inst_mx_inst_n93), .ZN(rout_x[34]) );
  XNOR2_X1 round_inst_mx_inst_U85 ( .A(round_inst_min_x[34]), .B(
        round_inst_min_x[38]), .ZN(round_inst_mx_inst_n93) );
  XNOR2_X1 round_inst_mx_inst_U84 ( .A(round_inst_min_x[28]), .B(
        round_inst_mx_inst_n92), .ZN(rout_x[28]) );
  XNOR2_X1 round_inst_mx_inst_U83 ( .A(round_inst_min_x[20]), .B(
        round_inst_mx_inst_n92), .ZN(rout_x[20]) );
  XNOR2_X1 round_inst_mx_inst_U82 ( .A(round_inst_min_x[24]), .B(
        round_inst_min_x[16]), .ZN(round_inst_mx_inst_n92) );
  XNOR2_X1 round_inst_mx_inst_U81 ( .A(round_inst_min_x[31]), .B(
        round_inst_mx_inst_n91), .ZN(rout_x[27]) );
  XNOR2_X1 round_inst_mx_inst_U80 ( .A(round_inst_min_x[23]), .B(
        round_inst_mx_inst_n91), .ZN(rout_x[19]) );
  XNOR2_X1 round_inst_mx_inst_U79 ( .A(round_inst_min_x[19]), .B(
        round_inst_min_x[27]), .ZN(round_inst_mx_inst_n91) );
  XNOR2_X1 round_inst_mx_inst_U78 ( .A(round_inst_min_x[45]), .B(
        round_inst_mx_inst_n90), .ZN(rout_x[45]) );
  XNOR2_X1 round_inst_mx_inst_U77 ( .A(round_inst_min_x[41]), .B(
        round_inst_mx_inst_n90), .ZN(rout_x[41]) );
  XNOR2_X1 round_inst_mx_inst_U76 ( .A(round_inst_min_x[33]), .B(
        round_inst_min_x[37]), .ZN(round_inst_mx_inst_n90) );
  XNOR2_X1 round_inst_mx_inst_U75 ( .A(round_inst_min_x[22]), .B(
        round_inst_mx_inst_n89), .ZN(rout_x[26]) );
  XNOR2_X1 round_inst_mx_inst_U74 ( .A(round_inst_min_x[18]), .B(
        round_inst_mx_inst_n89), .ZN(rout_x[22]) );
  XNOR2_X1 round_inst_mx_inst_U73 ( .A(round_inst_min_x[30]), .B(
        round_inst_min_x[26]), .ZN(round_inst_mx_inst_n89) );
  XNOR2_X1 round_inst_mx_inst_U72 ( .A(round_inst_min_x[16]), .B(
        round_inst_mx_inst_n88), .ZN(rout_x[24]) );
  XNOR2_X1 round_inst_mx_inst_U71 ( .A(round_inst_min_x[24]), .B(
        round_inst_mx_inst_n88), .ZN(rout_x[16]) );
  XNOR2_X1 round_inst_mx_inst_U70 ( .A(round_inst_min_x[28]), .B(
        round_inst_min_x[20]), .ZN(round_inst_mx_inst_n88) );
  XNOR2_X1 round_inst_mx_inst_U69 ( .A(round_inst_min_x[55]), .B(
        round_inst_mx_inst_n87), .ZN(rout_x[59]) );
  XNOR2_X1 round_inst_mx_inst_U68 ( .A(round_inst_min_x[51]), .B(
        round_inst_mx_inst_n87), .ZN(rout_x[55]) );
  XNOR2_X1 round_inst_mx_inst_U67 ( .A(round_inst_min_x[59]), .B(
        round_inst_min_x[63]), .ZN(round_inst_mx_inst_n87) );
  XNOR2_X1 round_inst_mx_inst_U66 ( .A(round_inst_min_x[21]), .B(
        round_inst_mx_inst_n86), .ZN(rout_x[21]) );
  XNOR2_X1 round_inst_mx_inst_U65 ( .A(round_inst_min_x[17]), .B(
        round_inst_mx_inst_n86), .ZN(rout_x[17]) );
  XNOR2_X1 round_inst_mx_inst_U64 ( .A(round_inst_min_x[25]), .B(
        round_inst_min_x[29]), .ZN(round_inst_mx_inst_n86) );
  XNOR2_X1 round_inst_mx_inst_U63 ( .A(round_inst_min_x[7]), .B(
        round_inst_mx_inst_n85), .ZN(rout_x[15]) );
  XNOR2_X1 round_inst_mx_inst_U62 ( .A(round_inst_min_x[15]), .B(
        round_inst_mx_inst_n85), .ZN(rout_x[7]) );
  XNOR2_X1 round_inst_mx_inst_U61 ( .A(round_inst_min_x[3]), .B(
        round_inst_min_x[11]), .ZN(round_inst_mx_inst_n85) );
  XNOR2_X1 round_inst_mx_inst_U60 ( .A(round_inst_min_x[44]), .B(
        round_inst_mx_inst_n84), .ZN(rout_x[44]) );
  XNOR2_X1 round_inst_mx_inst_U59 ( .A(round_inst_min_x[36]), .B(
        round_inst_mx_inst_n84), .ZN(rout_x[36]) );
  XNOR2_X1 round_inst_mx_inst_U58 ( .A(round_inst_min_x[40]), .B(
        round_inst_min_x[32]), .ZN(round_inst_mx_inst_n84) );
  XNOR2_X1 round_inst_mx_inst_U57 ( .A(round_inst_min_x[11]), .B(
        round_inst_mx_inst_n83), .ZN(rout_x[11]) );
  XNOR2_X1 round_inst_mx_inst_U56 ( .A(round_inst_min_x[3]), .B(
        round_inst_mx_inst_n83), .ZN(rout_x[3]) );
  XNOR2_X1 round_inst_mx_inst_U55 ( .A(round_inst_min_x[7]), .B(
        round_inst_min_x[15]), .ZN(round_inst_mx_inst_n83) );
  XNOR2_X1 round_inst_mx_inst_U54 ( .A(round_inst_min_x[6]), .B(
        round_inst_mx_inst_n82), .ZN(rout_x[14]) );
  XNOR2_X1 round_inst_mx_inst_U53 ( .A(round_inst_min_x[10]), .B(
        round_inst_mx_inst_n82), .ZN(rout_x[2]) );
  XNOR2_X1 round_inst_mx_inst_U52 ( .A(round_inst_min_x[14]), .B(
        round_inst_min_x[2]), .ZN(round_inst_mx_inst_n82) );
  XNOR2_X1 round_inst_mx_inst_U51 ( .A(round_inst_min_x[61]), .B(
        round_inst_mx_inst_n81), .ZN(rout_x[61]) );
  XNOR2_X1 round_inst_mx_inst_U50 ( .A(round_inst_min_x[53]), .B(
        round_inst_mx_inst_n81), .ZN(rout_x[53]) );
  XNOR2_X1 round_inst_mx_inst_U49 ( .A(round_inst_min_x[57]), .B(
        round_inst_min_x[49]), .ZN(round_inst_mx_inst_n81) );
  XNOR2_X1 round_inst_mx_inst_U48 ( .A(round_inst_min_x[49]), .B(
        round_inst_mx_inst_n80), .ZN(rout_x[57]) );
  XNOR2_X1 round_inst_mx_inst_U47 ( .A(round_inst_min_x[57]), .B(
        round_inst_mx_inst_n80), .ZN(rout_x[49]) );
  XNOR2_X1 round_inst_mx_inst_U46 ( .A(round_inst_min_x[61]), .B(
        round_inst_min_x[53]), .ZN(round_inst_mx_inst_n80) );
  XNOR2_X1 round_inst_mx_inst_U45 ( .A(round_inst_min_x[2]), .B(
        round_inst_mx_inst_n79), .ZN(rout_x[10]) );
  XNOR2_X1 round_inst_mx_inst_U44 ( .A(round_inst_min_x[14]), .B(
        round_inst_mx_inst_n79), .ZN(rout_x[6]) );
  XNOR2_X1 round_inst_mx_inst_U43 ( .A(round_inst_min_x[6]), .B(
        round_inst_min_x[10]), .ZN(round_inst_mx_inst_n79) );
  XNOR2_X1 round_inst_mx_inst_U42 ( .A(round_inst_min_x[9]), .B(
        round_inst_mx_inst_n78), .ZN(rout_x[13]) );
  XNOR2_X1 round_inst_mx_inst_U41 ( .A(round_inst_min_x[5]), .B(
        round_inst_mx_inst_n78), .ZN(rout_x[9]) );
  XNOR2_X1 round_inst_mx_inst_U40 ( .A(round_inst_min_x[13]), .B(
        round_inst_min_x[1]), .ZN(round_inst_mx_inst_n78) );
  XNOR2_X1 round_inst_mx_inst_U39 ( .A(round_inst_min_x[47]), .B(
        round_inst_mx_inst_n77), .ZN(rout_x[43]) );
  XNOR2_X1 round_inst_mx_inst_U38 ( .A(round_inst_min_x[39]), .B(
        round_inst_mx_inst_n77), .ZN(rout_x[35]) );
  XNOR2_X1 round_inst_mx_inst_U37 ( .A(round_inst_min_x[35]), .B(
        round_inst_min_x[43]), .ZN(round_inst_mx_inst_n77) );
  XNOR2_X1 round_inst_mx_inst_U36 ( .A(round_inst_min_x[8]), .B(
        round_inst_mx_inst_n76), .ZN(rout_x[12]) );
  XNOR2_X1 round_inst_mx_inst_U35 ( .A(round_inst_min_x[0]), .B(
        round_inst_mx_inst_n76), .ZN(rout_x[4]) );
  XNOR2_X1 round_inst_mx_inst_U34 ( .A(round_inst_min_x[4]), .B(
        round_inst_min_x[12]), .ZN(round_inst_mx_inst_n76) );
  XNOR2_X1 round_inst_mx_inst_U33 ( .A(round_inst_min_x[56]), .B(
        round_inst_mx_inst_n75), .ZN(rout_x[56]) );
  XNOR2_X1 round_inst_mx_inst_U32 ( .A(round_inst_min_x[52]), .B(
        round_inst_mx_inst_n75), .ZN(rout_x[52]) );
  XNOR2_X1 round_inst_mx_inst_U31 ( .A(round_inst_min_x[60]), .B(
        round_inst_min_x[48]), .ZN(round_inst_mx_inst_n75) );
  XNOR2_X1 round_inst_mx_inst_U30 ( .A(round_inst_min_x[38]), .B(
        round_inst_mx_inst_n74), .ZN(rout_x[42]) );
  XNOR2_X1 round_inst_mx_inst_U29 ( .A(round_inst_min_x[34]), .B(
        round_inst_mx_inst_n74), .ZN(rout_x[38]) );
  XNOR2_X1 round_inst_mx_inst_U28 ( .A(round_inst_min_x[42]), .B(
        round_inst_min_x[46]), .ZN(round_inst_mx_inst_n74) );
  XNOR2_X1 round_inst_mx_inst_U27 ( .A(round_inst_min_x[32]), .B(
        round_inst_mx_inst_n73), .ZN(rout_x[40]) );
  XNOR2_X1 round_inst_mx_inst_U26 ( .A(round_inst_min_x[40]), .B(
        round_inst_mx_inst_n73), .ZN(rout_x[32]) );
  XNOR2_X1 round_inst_mx_inst_U25 ( .A(round_inst_min_x[44]), .B(
        round_inst_min_x[36]), .ZN(round_inst_mx_inst_n73) );
  XNOR2_X1 round_inst_mx_inst_U24 ( .A(round_inst_min_x[1]), .B(
        round_inst_mx_inst_n72), .ZN(rout_x[5]) );
  XNOR2_X1 round_inst_mx_inst_U23 ( .A(round_inst_min_x[13]), .B(
        round_inst_mx_inst_n72), .ZN(rout_x[1]) );
  XNOR2_X1 round_inst_mx_inst_U22 ( .A(round_inst_min_x[9]), .B(
        round_inst_min_x[5]), .ZN(round_inst_mx_inst_n72) );
  XNOR2_X1 round_inst_mx_inst_U21 ( .A(round_inst_min_x[12]), .B(
        round_inst_mx_inst_n71), .ZN(rout_x[8]) );
  XNOR2_X1 round_inst_mx_inst_U20 ( .A(round_inst_min_x[4]), .B(
        round_inst_mx_inst_n71), .ZN(rout_x[0]) );
  XNOR2_X1 round_inst_mx_inst_U19 ( .A(round_inst_min_x[8]), .B(
        round_inst_min_x[0]), .ZN(round_inst_mx_inst_n71) );
  XNOR2_X1 round_inst_mx_inst_U18 ( .A(round_inst_min_x[54]), .B(
        round_inst_mx_inst_n70), .ZN(rout_x[54]) );
  XNOR2_X1 round_inst_mx_inst_U17 ( .A(round_inst_min_x[50]), .B(
        round_inst_mx_inst_n70), .ZN(rout_x[50]) );
  XNOR2_X1 round_inst_mx_inst_U16 ( .A(round_inst_min_x[62]), .B(
        round_inst_min_x[58]), .ZN(round_inst_mx_inst_n70) );
  XNOR2_X1 round_inst_mx_inst_U15 ( .A(round_inst_min_x[37]), .B(
        round_inst_mx_inst_n69), .ZN(rout_x[37]) );
  XNOR2_X1 round_inst_mx_inst_U14 ( .A(round_inst_min_x[33]), .B(
        round_inst_mx_inst_n69), .ZN(rout_x[33]) );
  XNOR2_X1 round_inst_mx_inst_U13 ( .A(round_inst_min_x[45]), .B(
        round_inst_min_x[41]), .ZN(round_inst_mx_inst_n69) );
  XNOR2_X1 round_inst_mx_inst_U12 ( .A(round_inst_min_x[27]), .B(
        round_inst_mx_inst_n68), .ZN(rout_x[31]) );
  XNOR2_X1 round_inst_mx_inst_U11 ( .A(round_inst_min_x[19]), .B(
        round_inst_mx_inst_n68), .ZN(rout_x[23]) );
  XNOR2_X1 round_inst_mx_inst_U10 ( .A(round_inst_min_x[31]), .B(
        round_inst_min_x[23]), .ZN(round_inst_mx_inst_n68) );
  XNOR2_X1 round_inst_mx_inst_U9 ( .A(round_inst_min_x[43]), .B(
        round_inst_mx_inst_n67), .ZN(rout_x[47]) );
  XNOR2_X1 round_inst_mx_inst_U8 ( .A(round_inst_min_x[35]), .B(
        round_inst_mx_inst_n67), .ZN(rout_x[39]) );
  XNOR2_X1 round_inst_mx_inst_U7 ( .A(round_inst_min_x[47]), .B(
        round_inst_min_x[39]), .ZN(round_inst_mx_inst_n67) );
  XNOR2_X1 round_inst_mx_inst_U6 ( .A(round_inst_min_x[26]), .B(
        round_inst_mx_inst_n66), .ZN(rout_x[30]) );
  XNOR2_X1 round_inst_mx_inst_U5 ( .A(round_inst_min_x[30]), .B(
        round_inst_mx_inst_n66), .ZN(rout_x[18]) );
  XNOR2_X1 round_inst_mx_inst_U4 ( .A(round_inst_min_x[22]), .B(
        round_inst_min_x[18]), .ZN(round_inst_mx_inst_n66) );
  XNOR2_X1 round_inst_mx_inst_U3 ( .A(round_inst_min_x[29]), .B(
        round_inst_mx_inst_n65), .ZN(rout_x[29]) );
  XNOR2_X1 round_inst_mx_inst_U2 ( .A(round_inst_min_x[25]), .B(
        round_inst_mx_inst_n65), .ZN(rout_x[25]) );
  XNOR2_X1 round_inst_mx_inst_U1 ( .A(round_inst_min_x[21]), .B(
        round_inst_min_x[17]), .ZN(round_inst_mx_inst_n65) );
  XNOR2_X1 round_inst_my_inst_U96 ( .A(round_inst_min_y[59]), .B(
        round_inst_my_inst_n96), .ZN(rout_y[63]) );
  XNOR2_X1 round_inst_my_inst_U95 ( .A(round_inst_min_y[63]), .B(
        round_inst_my_inst_n96), .ZN(rout_y[51]) );
  XNOR2_X1 round_inst_my_inst_U94 ( .A(round_inst_min_y[51]), .B(
        round_inst_min_y[55]), .ZN(round_inst_my_inst_n96) );
  XNOR2_X1 round_inst_my_inst_U93 ( .A(round_inst_min_y[62]), .B(
        round_inst_my_inst_n95), .ZN(rout_y[62]) );
  XNOR2_X1 round_inst_my_inst_U92 ( .A(round_inst_min_y[58]), .B(
        round_inst_my_inst_n95), .ZN(rout_y[58]) );
  XNOR2_X1 round_inst_my_inst_U91 ( .A(round_inst_min_y[50]), .B(
        round_inst_min_y[54]), .ZN(round_inst_my_inst_n95) );
  XNOR2_X1 round_inst_my_inst_U90 ( .A(round_inst_min_y[60]), .B(
        round_inst_my_inst_n94), .ZN(rout_y[60]) );
  XNOR2_X1 round_inst_my_inst_U89 ( .A(round_inst_min_y[48]), .B(
        round_inst_my_inst_n94), .ZN(rout_y[48]) );
  XNOR2_X1 round_inst_my_inst_U88 ( .A(round_inst_min_y[52]), .B(
        round_inst_min_y[56]), .ZN(round_inst_my_inst_n94) );
  XNOR2_X1 round_inst_my_inst_U87 ( .A(round_inst_min_y[42]), .B(
        round_inst_my_inst_n93), .ZN(rout_y[46]) );
  XNOR2_X1 round_inst_my_inst_U86 ( .A(round_inst_min_y[46]), .B(
        round_inst_my_inst_n93), .ZN(rout_y[34]) );
  XNOR2_X1 round_inst_my_inst_U85 ( .A(round_inst_min_y[34]), .B(
        round_inst_min_y[38]), .ZN(round_inst_my_inst_n93) );
  XNOR2_X1 round_inst_my_inst_U84 ( .A(round_inst_min_y[28]), .B(
        round_inst_my_inst_n92), .ZN(rout_y[28]) );
  XNOR2_X1 round_inst_my_inst_U83 ( .A(round_inst_min_y[20]), .B(
        round_inst_my_inst_n92), .ZN(rout_y[20]) );
  XNOR2_X1 round_inst_my_inst_U82 ( .A(round_inst_min_y[24]), .B(
        round_inst_min_y[16]), .ZN(round_inst_my_inst_n92) );
  XNOR2_X1 round_inst_my_inst_U81 ( .A(round_inst_min_y[31]), .B(
        round_inst_my_inst_n91), .ZN(rout_y[27]) );
  XNOR2_X1 round_inst_my_inst_U80 ( .A(round_inst_min_y[23]), .B(
        round_inst_my_inst_n91), .ZN(rout_y[19]) );
  XNOR2_X1 round_inst_my_inst_U79 ( .A(round_inst_min_y[19]), .B(
        round_inst_min_y[27]), .ZN(round_inst_my_inst_n91) );
  XNOR2_X1 round_inst_my_inst_U78 ( .A(round_inst_min_y[45]), .B(
        round_inst_my_inst_n90), .ZN(rout_y[45]) );
  XNOR2_X1 round_inst_my_inst_U77 ( .A(round_inst_min_y[41]), .B(
        round_inst_my_inst_n90), .ZN(rout_y[41]) );
  XNOR2_X1 round_inst_my_inst_U76 ( .A(round_inst_min_y[33]), .B(
        round_inst_min_y[37]), .ZN(round_inst_my_inst_n90) );
  XNOR2_X1 round_inst_my_inst_U75 ( .A(round_inst_min_y[22]), .B(
        round_inst_my_inst_n89), .ZN(rout_y[26]) );
  XNOR2_X1 round_inst_my_inst_U74 ( .A(round_inst_min_y[18]), .B(
        round_inst_my_inst_n89), .ZN(rout_y[22]) );
  XNOR2_X1 round_inst_my_inst_U73 ( .A(round_inst_min_y[30]), .B(
        round_inst_min_y[26]), .ZN(round_inst_my_inst_n89) );
  XNOR2_X1 round_inst_my_inst_U72 ( .A(round_inst_min_y[16]), .B(
        round_inst_my_inst_n88), .ZN(rout_y[24]) );
  XNOR2_X1 round_inst_my_inst_U71 ( .A(round_inst_min_y[24]), .B(
        round_inst_my_inst_n88), .ZN(rout_y[16]) );
  XNOR2_X1 round_inst_my_inst_U70 ( .A(round_inst_min_y[28]), .B(
        round_inst_min_y[20]), .ZN(round_inst_my_inst_n88) );
  XNOR2_X1 round_inst_my_inst_U69 ( .A(round_inst_min_y[55]), .B(
        round_inst_my_inst_n87), .ZN(rout_y[59]) );
  XNOR2_X1 round_inst_my_inst_U68 ( .A(round_inst_min_y[51]), .B(
        round_inst_my_inst_n87), .ZN(rout_y[55]) );
  XNOR2_X1 round_inst_my_inst_U67 ( .A(round_inst_min_y[59]), .B(
        round_inst_min_y[63]), .ZN(round_inst_my_inst_n87) );
  XNOR2_X1 round_inst_my_inst_U66 ( .A(round_inst_min_y[21]), .B(
        round_inst_my_inst_n86), .ZN(rout_y[21]) );
  XNOR2_X1 round_inst_my_inst_U65 ( .A(round_inst_min_y[17]), .B(
        round_inst_my_inst_n86), .ZN(rout_y[17]) );
  XNOR2_X1 round_inst_my_inst_U64 ( .A(round_inst_min_y[25]), .B(
        round_inst_min_y[29]), .ZN(round_inst_my_inst_n86) );
  XNOR2_X1 round_inst_my_inst_U63 ( .A(round_inst_min_y[7]), .B(
        round_inst_my_inst_n85), .ZN(rout_y[15]) );
  XNOR2_X1 round_inst_my_inst_U62 ( .A(round_inst_min_y[15]), .B(
        round_inst_my_inst_n85), .ZN(rout_y[7]) );
  XNOR2_X1 round_inst_my_inst_U61 ( .A(round_inst_min_y[3]), .B(
        round_inst_min_y[11]), .ZN(round_inst_my_inst_n85) );
  XNOR2_X1 round_inst_my_inst_U60 ( .A(round_inst_min_y[44]), .B(
        round_inst_my_inst_n84), .ZN(rout_y[44]) );
  XNOR2_X1 round_inst_my_inst_U59 ( .A(round_inst_min_y[36]), .B(
        round_inst_my_inst_n84), .ZN(rout_y[36]) );
  XNOR2_X1 round_inst_my_inst_U58 ( .A(round_inst_min_y[40]), .B(
        round_inst_min_y[32]), .ZN(round_inst_my_inst_n84) );
  XNOR2_X1 round_inst_my_inst_U57 ( .A(round_inst_min_y[11]), .B(
        round_inst_my_inst_n83), .ZN(rout_y[11]) );
  XNOR2_X1 round_inst_my_inst_U56 ( .A(round_inst_min_y[3]), .B(
        round_inst_my_inst_n83), .ZN(rout_y[3]) );
  XNOR2_X1 round_inst_my_inst_U55 ( .A(round_inst_min_y[7]), .B(
        round_inst_min_y[15]), .ZN(round_inst_my_inst_n83) );
  XNOR2_X1 round_inst_my_inst_U54 ( .A(round_inst_min_y[6]), .B(
        round_inst_my_inst_n82), .ZN(rout_y[14]) );
  XNOR2_X1 round_inst_my_inst_U53 ( .A(round_inst_min_y[10]), .B(
        round_inst_my_inst_n82), .ZN(rout_y[2]) );
  XNOR2_X1 round_inst_my_inst_U52 ( .A(round_inst_min_y[14]), .B(
        round_inst_min_y[2]), .ZN(round_inst_my_inst_n82) );
  XNOR2_X1 round_inst_my_inst_U51 ( .A(round_inst_min_y[61]), .B(
        round_inst_my_inst_n81), .ZN(rout_y[61]) );
  XNOR2_X1 round_inst_my_inst_U50 ( .A(round_inst_min_y[53]), .B(
        round_inst_my_inst_n81), .ZN(rout_y[53]) );
  XNOR2_X1 round_inst_my_inst_U49 ( .A(round_inst_min_y[57]), .B(
        round_inst_min_y[49]), .ZN(round_inst_my_inst_n81) );
  XNOR2_X1 round_inst_my_inst_U48 ( .A(round_inst_min_y[49]), .B(
        round_inst_my_inst_n80), .ZN(rout_y[57]) );
  XNOR2_X1 round_inst_my_inst_U47 ( .A(round_inst_min_y[57]), .B(
        round_inst_my_inst_n80), .ZN(rout_y[49]) );
  XNOR2_X1 round_inst_my_inst_U46 ( .A(round_inst_min_y[61]), .B(
        round_inst_min_y[53]), .ZN(round_inst_my_inst_n80) );
  XNOR2_X1 round_inst_my_inst_U45 ( .A(round_inst_min_y[2]), .B(
        round_inst_my_inst_n79), .ZN(rout_y[10]) );
  XNOR2_X1 round_inst_my_inst_U44 ( .A(round_inst_min_y[14]), .B(
        round_inst_my_inst_n79), .ZN(rout_y[6]) );
  XNOR2_X1 round_inst_my_inst_U43 ( .A(round_inst_min_y[6]), .B(
        round_inst_min_y[10]), .ZN(round_inst_my_inst_n79) );
  XNOR2_X1 round_inst_my_inst_U42 ( .A(round_inst_min_y[9]), .B(
        round_inst_my_inst_n78), .ZN(rout_y[13]) );
  XNOR2_X1 round_inst_my_inst_U41 ( .A(round_inst_min_y[5]), .B(
        round_inst_my_inst_n78), .ZN(rout_y[9]) );
  XNOR2_X1 round_inst_my_inst_U40 ( .A(round_inst_min_y[13]), .B(
        round_inst_min_y[1]), .ZN(round_inst_my_inst_n78) );
  XNOR2_X1 round_inst_my_inst_U39 ( .A(round_inst_min_y[47]), .B(
        round_inst_my_inst_n77), .ZN(rout_y[43]) );
  XNOR2_X1 round_inst_my_inst_U38 ( .A(round_inst_min_y[39]), .B(
        round_inst_my_inst_n77), .ZN(rout_y[35]) );
  XNOR2_X1 round_inst_my_inst_U37 ( .A(round_inst_min_y[35]), .B(
        round_inst_min_y[43]), .ZN(round_inst_my_inst_n77) );
  XNOR2_X1 round_inst_my_inst_U36 ( .A(round_inst_min_y[8]), .B(
        round_inst_my_inst_n76), .ZN(rout_y[12]) );
  XNOR2_X1 round_inst_my_inst_U35 ( .A(round_inst_min_y[0]), .B(
        round_inst_my_inst_n76), .ZN(rout_y[4]) );
  XNOR2_X1 round_inst_my_inst_U34 ( .A(round_inst_min_y[4]), .B(
        round_inst_min_y[12]), .ZN(round_inst_my_inst_n76) );
  XNOR2_X1 round_inst_my_inst_U33 ( .A(round_inst_min_y[56]), .B(
        round_inst_my_inst_n75), .ZN(rout_y[56]) );
  XNOR2_X1 round_inst_my_inst_U32 ( .A(round_inst_min_y[52]), .B(
        round_inst_my_inst_n75), .ZN(rout_y[52]) );
  XNOR2_X1 round_inst_my_inst_U31 ( .A(round_inst_min_y[60]), .B(
        round_inst_min_y[48]), .ZN(round_inst_my_inst_n75) );
  XNOR2_X1 round_inst_my_inst_U30 ( .A(round_inst_min_y[38]), .B(
        round_inst_my_inst_n74), .ZN(rout_y[42]) );
  XNOR2_X1 round_inst_my_inst_U29 ( .A(round_inst_min_y[34]), .B(
        round_inst_my_inst_n74), .ZN(rout_y[38]) );
  XNOR2_X1 round_inst_my_inst_U28 ( .A(round_inst_min_y[42]), .B(
        round_inst_min_y[46]), .ZN(round_inst_my_inst_n74) );
  XNOR2_X1 round_inst_my_inst_U27 ( .A(round_inst_min_y[32]), .B(
        round_inst_my_inst_n73), .ZN(rout_y[40]) );
  XNOR2_X1 round_inst_my_inst_U26 ( .A(round_inst_min_y[40]), .B(
        round_inst_my_inst_n73), .ZN(rout_y[32]) );
  XNOR2_X1 round_inst_my_inst_U25 ( .A(round_inst_min_y[44]), .B(
        round_inst_min_y[36]), .ZN(round_inst_my_inst_n73) );
  XNOR2_X1 round_inst_my_inst_U24 ( .A(round_inst_min_y[1]), .B(
        round_inst_my_inst_n72), .ZN(rout_y[5]) );
  XNOR2_X1 round_inst_my_inst_U23 ( .A(round_inst_min_y[13]), .B(
        round_inst_my_inst_n72), .ZN(rout_y[1]) );
  XNOR2_X1 round_inst_my_inst_U22 ( .A(round_inst_min_y[9]), .B(
        round_inst_min_y[5]), .ZN(round_inst_my_inst_n72) );
  XNOR2_X1 round_inst_my_inst_U21 ( .A(round_inst_min_y[12]), .B(
        round_inst_my_inst_n71), .ZN(rout_y[8]) );
  XNOR2_X1 round_inst_my_inst_U20 ( .A(round_inst_min_y[4]), .B(
        round_inst_my_inst_n71), .ZN(rout_y[0]) );
  XNOR2_X1 round_inst_my_inst_U19 ( .A(round_inst_min_y[8]), .B(
        round_inst_min_y[0]), .ZN(round_inst_my_inst_n71) );
  XNOR2_X1 round_inst_my_inst_U18 ( .A(round_inst_min_y[54]), .B(
        round_inst_my_inst_n70), .ZN(rout_y[54]) );
  XNOR2_X1 round_inst_my_inst_U17 ( .A(round_inst_min_y[50]), .B(
        round_inst_my_inst_n70), .ZN(rout_y[50]) );
  XNOR2_X1 round_inst_my_inst_U16 ( .A(round_inst_min_y[62]), .B(
        round_inst_min_y[58]), .ZN(round_inst_my_inst_n70) );
  XNOR2_X1 round_inst_my_inst_U15 ( .A(round_inst_min_y[37]), .B(
        round_inst_my_inst_n69), .ZN(rout_y[37]) );
  XNOR2_X1 round_inst_my_inst_U14 ( .A(round_inst_min_y[33]), .B(
        round_inst_my_inst_n69), .ZN(rout_y[33]) );
  XNOR2_X1 round_inst_my_inst_U13 ( .A(round_inst_min_y[45]), .B(
        round_inst_min_y[41]), .ZN(round_inst_my_inst_n69) );
  XNOR2_X1 round_inst_my_inst_U12 ( .A(round_inst_min_y[27]), .B(
        round_inst_my_inst_n68), .ZN(rout_y[31]) );
  XNOR2_X1 round_inst_my_inst_U11 ( .A(round_inst_min_y[19]), .B(
        round_inst_my_inst_n68), .ZN(rout_y[23]) );
  XNOR2_X1 round_inst_my_inst_U10 ( .A(round_inst_min_y[31]), .B(
        round_inst_min_y[23]), .ZN(round_inst_my_inst_n68) );
  XNOR2_X1 round_inst_my_inst_U9 ( .A(round_inst_min_y[43]), .B(
        round_inst_my_inst_n67), .ZN(rout_y[47]) );
  XNOR2_X1 round_inst_my_inst_U8 ( .A(round_inst_min_y[35]), .B(
        round_inst_my_inst_n67), .ZN(rout_y[39]) );
  XNOR2_X1 round_inst_my_inst_U7 ( .A(round_inst_min_y[47]), .B(
        round_inst_min_y[39]), .ZN(round_inst_my_inst_n67) );
  XNOR2_X1 round_inst_my_inst_U6 ( .A(round_inst_min_y[26]), .B(
        round_inst_my_inst_n66), .ZN(rout_y[30]) );
  XNOR2_X1 round_inst_my_inst_U5 ( .A(round_inst_min_y[30]), .B(
        round_inst_my_inst_n66), .ZN(rout_y[18]) );
  XNOR2_X1 round_inst_my_inst_U4 ( .A(round_inst_min_y[22]), .B(
        round_inst_min_y[18]), .ZN(round_inst_my_inst_n66) );
  XNOR2_X1 round_inst_my_inst_U3 ( .A(round_inst_min_y[29]), .B(
        round_inst_my_inst_n65), .ZN(rout_y[29]) );
  XNOR2_X1 round_inst_my_inst_U2 ( .A(round_inst_min_y[25]), .B(
        round_inst_my_inst_n65), .ZN(rout_y[25]) );
  XNOR2_X1 round_inst_my_inst_U1 ( .A(round_inst_min_y[21]), .B(
        round_inst_min_y[17]), .ZN(round_inst_my_inst_n65) );
  XNOR2_X1 round_inst_mz_inst_U96 ( .A(round_inst_min_z[59]), .B(
        round_inst_mz_inst_n96), .ZN(rout_z[63]) );
  XNOR2_X1 round_inst_mz_inst_U95 ( .A(round_inst_min_z[63]), .B(
        round_inst_mz_inst_n96), .ZN(rout_z[51]) );
  XNOR2_X1 round_inst_mz_inst_U94 ( .A(round_inst_min_z[51]), .B(
        round_inst_min_z[55]), .ZN(round_inst_mz_inst_n96) );
  XNOR2_X1 round_inst_mz_inst_U93 ( .A(round_inst_min_z[62]), .B(
        round_inst_mz_inst_n95), .ZN(rout_z[62]) );
  XNOR2_X1 round_inst_mz_inst_U92 ( .A(round_inst_min_z[58]), .B(
        round_inst_mz_inst_n95), .ZN(rout_z[58]) );
  XNOR2_X1 round_inst_mz_inst_U91 ( .A(round_inst_min_z[50]), .B(
        round_inst_min_z[54]), .ZN(round_inst_mz_inst_n95) );
  XNOR2_X1 round_inst_mz_inst_U90 ( .A(round_inst_min_z[60]), .B(
        round_inst_mz_inst_n94), .ZN(rout_z[60]) );
  XNOR2_X1 round_inst_mz_inst_U89 ( .A(round_inst_min_z[48]), .B(
        round_inst_mz_inst_n94), .ZN(rout_z[48]) );
  XNOR2_X1 round_inst_mz_inst_U88 ( .A(round_inst_min_z[52]), .B(
        round_inst_min_z[56]), .ZN(round_inst_mz_inst_n94) );
  XNOR2_X1 round_inst_mz_inst_U87 ( .A(round_inst_min_z[42]), .B(
        round_inst_mz_inst_n93), .ZN(rout_z[46]) );
  XNOR2_X1 round_inst_mz_inst_U86 ( .A(round_inst_min_z[46]), .B(
        round_inst_mz_inst_n93), .ZN(rout_z[34]) );
  XNOR2_X1 round_inst_mz_inst_U85 ( .A(round_inst_min_z[34]), .B(
        round_inst_min_z[38]), .ZN(round_inst_mz_inst_n93) );
  XNOR2_X1 round_inst_mz_inst_U84 ( .A(round_inst_min_z[28]), .B(
        round_inst_mz_inst_n92), .ZN(rout_z[28]) );
  XNOR2_X1 round_inst_mz_inst_U83 ( .A(round_inst_min_z[20]), .B(
        round_inst_mz_inst_n92), .ZN(rout_z[20]) );
  XNOR2_X1 round_inst_mz_inst_U82 ( .A(round_inst_min_z[24]), .B(
        round_inst_min_z[16]), .ZN(round_inst_mz_inst_n92) );
  XNOR2_X1 round_inst_mz_inst_U81 ( .A(round_inst_min_z[31]), .B(
        round_inst_mz_inst_n91), .ZN(rout_z[27]) );
  XNOR2_X1 round_inst_mz_inst_U80 ( .A(round_inst_min_z[23]), .B(
        round_inst_mz_inst_n91), .ZN(rout_z[19]) );
  XNOR2_X1 round_inst_mz_inst_U79 ( .A(round_inst_min_z[19]), .B(
        round_inst_min_z[27]), .ZN(round_inst_mz_inst_n91) );
  XNOR2_X1 round_inst_mz_inst_U78 ( .A(round_inst_min_z[45]), .B(
        round_inst_mz_inst_n90), .ZN(rout_z[45]) );
  XNOR2_X1 round_inst_mz_inst_U77 ( .A(round_inst_min_z[41]), .B(
        round_inst_mz_inst_n90), .ZN(rout_z[41]) );
  XNOR2_X1 round_inst_mz_inst_U76 ( .A(round_inst_min_z[33]), .B(
        round_inst_min_z[37]), .ZN(round_inst_mz_inst_n90) );
  XNOR2_X1 round_inst_mz_inst_U75 ( .A(round_inst_min_z[22]), .B(
        round_inst_mz_inst_n89), .ZN(rout_z[26]) );
  XNOR2_X1 round_inst_mz_inst_U74 ( .A(round_inst_min_z[18]), .B(
        round_inst_mz_inst_n89), .ZN(rout_z[22]) );
  XNOR2_X1 round_inst_mz_inst_U73 ( .A(round_inst_min_z[30]), .B(
        round_inst_min_z[26]), .ZN(round_inst_mz_inst_n89) );
  XNOR2_X1 round_inst_mz_inst_U72 ( .A(round_inst_min_z[16]), .B(
        round_inst_mz_inst_n88), .ZN(rout_z[24]) );
  XNOR2_X1 round_inst_mz_inst_U71 ( .A(round_inst_min_z[24]), .B(
        round_inst_mz_inst_n88), .ZN(rout_z[16]) );
  XNOR2_X1 round_inst_mz_inst_U70 ( .A(round_inst_min_z[28]), .B(
        round_inst_min_z[20]), .ZN(round_inst_mz_inst_n88) );
  XNOR2_X1 round_inst_mz_inst_U69 ( .A(round_inst_min_z[55]), .B(
        round_inst_mz_inst_n87), .ZN(rout_z[59]) );
  XNOR2_X1 round_inst_mz_inst_U68 ( .A(round_inst_min_z[51]), .B(
        round_inst_mz_inst_n87), .ZN(rout_z[55]) );
  XNOR2_X1 round_inst_mz_inst_U67 ( .A(round_inst_min_z[59]), .B(
        round_inst_min_z[63]), .ZN(round_inst_mz_inst_n87) );
  XNOR2_X1 round_inst_mz_inst_U66 ( .A(round_inst_min_z[21]), .B(
        round_inst_mz_inst_n86), .ZN(rout_z[21]) );
  XNOR2_X1 round_inst_mz_inst_U65 ( .A(round_inst_min_z[17]), .B(
        round_inst_mz_inst_n86), .ZN(rout_z[17]) );
  XNOR2_X1 round_inst_mz_inst_U64 ( .A(round_inst_min_z[25]), .B(
        round_inst_min_z[29]), .ZN(round_inst_mz_inst_n86) );
  XNOR2_X1 round_inst_mz_inst_U63 ( .A(round_inst_min_z[7]), .B(
        round_inst_mz_inst_n85), .ZN(rout_z[15]) );
  XNOR2_X1 round_inst_mz_inst_U62 ( .A(round_inst_min_z[15]), .B(
        round_inst_mz_inst_n85), .ZN(rout_z[7]) );
  XNOR2_X1 round_inst_mz_inst_U61 ( .A(round_inst_min_z[3]), .B(
        round_inst_min_z[11]), .ZN(round_inst_mz_inst_n85) );
  XNOR2_X1 round_inst_mz_inst_U60 ( .A(round_inst_min_z[44]), .B(
        round_inst_mz_inst_n84), .ZN(rout_z[44]) );
  XNOR2_X1 round_inst_mz_inst_U59 ( .A(round_inst_min_z[36]), .B(
        round_inst_mz_inst_n84), .ZN(rout_z[36]) );
  XNOR2_X1 round_inst_mz_inst_U58 ( .A(round_inst_min_z[40]), .B(
        round_inst_min_z[32]), .ZN(round_inst_mz_inst_n84) );
  XNOR2_X1 round_inst_mz_inst_U57 ( .A(round_inst_min_z[11]), .B(
        round_inst_mz_inst_n83), .ZN(rout_z[11]) );
  XNOR2_X1 round_inst_mz_inst_U56 ( .A(round_inst_min_z[3]), .B(
        round_inst_mz_inst_n83), .ZN(rout_z[3]) );
  XNOR2_X1 round_inst_mz_inst_U55 ( .A(round_inst_min_z[7]), .B(
        round_inst_min_z[15]), .ZN(round_inst_mz_inst_n83) );
  XNOR2_X1 round_inst_mz_inst_U54 ( .A(round_inst_min_z[6]), .B(
        round_inst_mz_inst_n82), .ZN(rout_z[14]) );
  XNOR2_X1 round_inst_mz_inst_U53 ( .A(round_inst_min_z[10]), .B(
        round_inst_mz_inst_n82), .ZN(rout_z[2]) );
  XNOR2_X1 round_inst_mz_inst_U52 ( .A(round_inst_min_z[14]), .B(
        round_inst_min_z[2]), .ZN(round_inst_mz_inst_n82) );
  XNOR2_X1 round_inst_mz_inst_U51 ( .A(round_inst_min_z[61]), .B(
        round_inst_mz_inst_n81), .ZN(rout_z[61]) );
  XNOR2_X1 round_inst_mz_inst_U50 ( .A(round_inst_min_z[53]), .B(
        round_inst_mz_inst_n81), .ZN(rout_z[53]) );
  XNOR2_X1 round_inst_mz_inst_U49 ( .A(round_inst_min_z[57]), .B(
        round_inst_min_z[49]), .ZN(round_inst_mz_inst_n81) );
  XNOR2_X1 round_inst_mz_inst_U48 ( .A(round_inst_min_z[49]), .B(
        round_inst_mz_inst_n80), .ZN(rout_z[57]) );
  XNOR2_X1 round_inst_mz_inst_U47 ( .A(round_inst_min_z[57]), .B(
        round_inst_mz_inst_n80), .ZN(rout_z[49]) );
  XNOR2_X1 round_inst_mz_inst_U46 ( .A(round_inst_min_z[61]), .B(
        round_inst_min_z[53]), .ZN(round_inst_mz_inst_n80) );
  XNOR2_X1 round_inst_mz_inst_U45 ( .A(round_inst_min_z[2]), .B(
        round_inst_mz_inst_n79), .ZN(rout_z[10]) );
  XNOR2_X1 round_inst_mz_inst_U44 ( .A(round_inst_min_z[14]), .B(
        round_inst_mz_inst_n79), .ZN(rout_z[6]) );
  XNOR2_X1 round_inst_mz_inst_U43 ( .A(round_inst_min_z[6]), .B(
        round_inst_min_z[10]), .ZN(round_inst_mz_inst_n79) );
  XNOR2_X1 round_inst_mz_inst_U42 ( .A(round_inst_min_z[9]), .B(
        round_inst_mz_inst_n78), .ZN(rout_z[13]) );
  XNOR2_X1 round_inst_mz_inst_U41 ( .A(round_inst_min_z[5]), .B(
        round_inst_mz_inst_n78), .ZN(rout_z[9]) );
  XNOR2_X1 round_inst_mz_inst_U40 ( .A(round_inst_min_z[13]), .B(
        round_inst_min_z[1]), .ZN(round_inst_mz_inst_n78) );
  XNOR2_X1 round_inst_mz_inst_U39 ( .A(round_inst_min_z[47]), .B(
        round_inst_mz_inst_n77), .ZN(rout_z[43]) );
  XNOR2_X1 round_inst_mz_inst_U38 ( .A(round_inst_min_z[39]), .B(
        round_inst_mz_inst_n77), .ZN(rout_z[35]) );
  XNOR2_X1 round_inst_mz_inst_U37 ( .A(round_inst_min_z[35]), .B(
        round_inst_min_z[43]), .ZN(round_inst_mz_inst_n77) );
  XNOR2_X1 round_inst_mz_inst_U36 ( .A(round_inst_min_z[8]), .B(
        round_inst_mz_inst_n76), .ZN(rout_z[12]) );
  XNOR2_X1 round_inst_mz_inst_U35 ( .A(round_inst_min_z[0]), .B(
        round_inst_mz_inst_n76), .ZN(rout_z[4]) );
  XNOR2_X1 round_inst_mz_inst_U34 ( .A(round_inst_min_z[4]), .B(
        round_inst_min_z[12]), .ZN(round_inst_mz_inst_n76) );
  XNOR2_X1 round_inst_mz_inst_U33 ( .A(round_inst_min_z[56]), .B(
        round_inst_mz_inst_n75), .ZN(rout_z[56]) );
  XNOR2_X1 round_inst_mz_inst_U32 ( .A(round_inst_min_z[52]), .B(
        round_inst_mz_inst_n75), .ZN(rout_z[52]) );
  XNOR2_X1 round_inst_mz_inst_U31 ( .A(round_inst_min_z[60]), .B(
        round_inst_min_z[48]), .ZN(round_inst_mz_inst_n75) );
  XNOR2_X1 round_inst_mz_inst_U30 ( .A(round_inst_min_z[38]), .B(
        round_inst_mz_inst_n74), .ZN(rout_z[42]) );
  XNOR2_X1 round_inst_mz_inst_U29 ( .A(round_inst_min_z[34]), .B(
        round_inst_mz_inst_n74), .ZN(rout_z[38]) );
  XNOR2_X1 round_inst_mz_inst_U28 ( .A(round_inst_min_z[42]), .B(
        round_inst_min_z[46]), .ZN(round_inst_mz_inst_n74) );
  XNOR2_X1 round_inst_mz_inst_U27 ( .A(round_inst_min_z[32]), .B(
        round_inst_mz_inst_n73), .ZN(rout_z[40]) );
  XNOR2_X1 round_inst_mz_inst_U26 ( .A(round_inst_min_z[40]), .B(
        round_inst_mz_inst_n73), .ZN(rout_z[32]) );
  XNOR2_X1 round_inst_mz_inst_U25 ( .A(round_inst_min_z[44]), .B(
        round_inst_min_z[36]), .ZN(round_inst_mz_inst_n73) );
  XNOR2_X1 round_inst_mz_inst_U24 ( .A(round_inst_min_z[1]), .B(
        round_inst_mz_inst_n72), .ZN(rout_z[5]) );
  XNOR2_X1 round_inst_mz_inst_U23 ( .A(round_inst_min_z[13]), .B(
        round_inst_mz_inst_n72), .ZN(rout_z[1]) );
  XNOR2_X1 round_inst_mz_inst_U22 ( .A(round_inst_min_z[9]), .B(
        round_inst_min_z[5]), .ZN(round_inst_mz_inst_n72) );
  XNOR2_X1 round_inst_mz_inst_U21 ( .A(round_inst_min_z[12]), .B(
        round_inst_mz_inst_n71), .ZN(rout_z[8]) );
  XNOR2_X1 round_inst_mz_inst_U20 ( .A(round_inst_min_z[4]), .B(
        round_inst_mz_inst_n71), .ZN(rout_z[0]) );
  XNOR2_X1 round_inst_mz_inst_U19 ( .A(round_inst_min_z[8]), .B(
        round_inst_min_z[0]), .ZN(round_inst_mz_inst_n71) );
  XNOR2_X1 round_inst_mz_inst_U18 ( .A(round_inst_min_z[54]), .B(
        round_inst_mz_inst_n70), .ZN(rout_z[54]) );
  XNOR2_X1 round_inst_mz_inst_U17 ( .A(round_inst_min_z[50]), .B(
        round_inst_mz_inst_n70), .ZN(rout_z[50]) );
  XNOR2_X1 round_inst_mz_inst_U16 ( .A(round_inst_min_z[62]), .B(
        round_inst_min_z[58]), .ZN(round_inst_mz_inst_n70) );
  XNOR2_X1 round_inst_mz_inst_U15 ( .A(round_inst_min_z[37]), .B(
        round_inst_mz_inst_n69), .ZN(rout_z[37]) );
  XNOR2_X1 round_inst_mz_inst_U14 ( .A(round_inst_min_z[33]), .B(
        round_inst_mz_inst_n69), .ZN(rout_z[33]) );
  XNOR2_X1 round_inst_mz_inst_U13 ( .A(round_inst_min_z[45]), .B(
        round_inst_min_z[41]), .ZN(round_inst_mz_inst_n69) );
  XNOR2_X1 round_inst_mz_inst_U12 ( .A(round_inst_min_z[27]), .B(
        round_inst_mz_inst_n68), .ZN(rout_z[31]) );
  XNOR2_X1 round_inst_mz_inst_U11 ( .A(round_inst_min_z[19]), .B(
        round_inst_mz_inst_n68), .ZN(rout_z[23]) );
  XNOR2_X1 round_inst_mz_inst_U10 ( .A(round_inst_min_z[31]), .B(
        round_inst_min_z[23]), .ZN(round_inst_mz_inst_n68) );
  XNOR2_X1 round_inst_mz_inst_U9 ( .A(round_inst_min_z[43]), .B(
        round_inst_mz_inst_n67), .ZN(rout_z[47]) );
  XNOR2_X1 round_inst_mz_inst_U8 ( .A(round_inst_min_z[35]), .B(
        round_inst_mz_inst_n67), .ZN(rout_z[39]) );
  XNOR2_X1 round_inst_mz_inst_U7 ( .A(round_inst_min_z[47]), .B(
        round_inst_min_z[39]), .ZN(round_inst_mz_inst_n67) );
  XNOR2_X1 round_inst_mz_inst_U6 ( .A(round_inst_min_z[26]), .B(
        round_inst_mz_inst_n66), .ZN(rout_z[30]) );
  XNOR2_X1 round_inst_mz_inst_U5 ( .A(round_inst_min_z[30]), .B(
        round_inst_mz_inst_n66), .ZN(rout_z[18]) );
  XNOR2_X1 round_inst_mz_inst_U4 ( .A(round_inst_min_z[22]), .B(
        round_inst_min_z[18]), .ZN(round_inst_mz_inst_n66) );
  XNOR2_X1 round_inst_mz_inst_U3 ( .A(round_inst_min_z[29]), .B(
        round_inst_mz_inst_n65), .ZN(rout_z[29]) );
  XNOR2_X1 round_inst_mz_inst_U2 ( .A(round_inst_min_z[25]), .B(
        round_inst_mz_inst_n65), .ZN(rout_z[25]) );
  XNOR2_X1 round_inst_mz_inst_U1 ( .A(round_inst_min_z[21]), .B(
        round_inst_min_z[17]), .ZN(round_inst_mz_inst_n65) );
  AND2_X1 mux_c0_U67 ( .A1(mux_c0_n265), .A2(final_w_k[0]), .ZN(c0[0]) );
  AND2_X1 mux_c0_U66 ( .A1(mux_c0_n265), .A2(final_w_k[1]), .ZN(c0[1]) );
  AND2_X1 mux_c0_U65 ( .A1(done), .A2(final_w_k[44]), .ZN(c0[44]) );
  AND2_X1 mux_c0_U64 ( .A1(mux_c0_n265), .A2(final_w_k[2]), .ZN(c0[2]) );
  AND2_X1 mux_c0_U63 ( .A1(mux_c0_n265), .A2(final_w_k[3]), .ZN(c0[3]) );
  AND2_X1 mux_c0_U62 ( .A1(mux_c0_n265), .A2(final_w_k[4]), .ZN(c0[4]) );
  AND2_X1 mux_c0_U61 ( .A1(mux_c0_n265), .A2(final_w_k[5]), .ZN(c0[5]) );
  AND2_X1 mux_c0_U60 ( .A1(mux_c0_n265), .A2(final_w_k[6]), .ZN(c0[6]) );
  AND2_X1 mux_c0_U59 ( .A1(mux_c0_n265), .A2(final_w_k[7]), .ZN(c0[7]) );
  AND2_X1 mux_c0_U58 ( .A1(mux_c0_n265), .A2(final_w_k[8]), .ZN(c0[8]) );
  AND2_X1 mux_c0_U57 ( .A1(mux_c0_n265), .A2(final_w_k[9]), .ZN(c0[9]) );
  AND2_X1 mux_c0_U56 ( .A1(mux_c0_n265), .A2(final_w_k[10]), .ZN(c0[10]) );
  AND2_X1 mux_c0_U55 ( .A1(mux_c0_n265), .A2(final_w_k[11]), .ZN(c0[11]) );
  AND2_X1 mux_c0_U54 ( .A1(mux_c0_n264), .A2(final_w_k[12]), .ZN(c0[12]) );
  AND2_X1 mux_c0_U53 ( .A1(done), .A2(final_w_k[13]), .ZN(c0[13]) );
  AND2_X1 mux_c0_U52 ( .A1(mux_c0_n265), .A2(final_w_k[14]), .ZN(c0[14]) );
  AND2_X1 mux_c0_U51 ( .A1(mux_c0_n264), .A2(final_w_k[15]), .ZN(c0[15]) );
  AND2_X1 mux_c0_U50 ( .A1(done), .A2(final_w_k[16]), .ZN(c0[16]) );
  AND2_X1 mux_c0_U49 ( .A1(mux_c0_n265), .A2(final_w_k[17]), .ZN(c0[17]) );
  AND2_X1 mux_c0_U48 ( .A1(mux_c0_n264), .A2(final_w_k[18]), .ZN(c0[18]) );
  AND2_X1 mux_c0_U47 ( .A1(done), .A2(final_w_k[19]), .ZN(c0[19]) );
  AND2_X1 mux_c0_U46 ( .A1(mux_c0_n265), .A2(final_w_k[20]), .ZN(c0[20]) );
  AND2_X1 mux_c0_U45 ( .A1(mux_c0_n264), .A2(final_w_k[21]), .ZN(c0[21]) );
  AND2_X1 mux_c0_U44 ( .A1(done), .A2(final_w_k[22]), .ZN(c0[22]) );
  AND2_X1 mux_c0_U43 ( .A1(mux_c0_n265), .A2(final_w_k[23]), .ZN(c0[23]) );
  AND2_X1 mux_c0_U42 ( .A1(mux_c0_n264), .A2(final_w_k[24]), .ZN(c0[24]) );
  AND2_X1 mux_c0_U41 ( .A1(done), .A2(final_w_k[25]), .ZN(c0[25]) );
  AND2_X1 mux_c0_U40 ( .A1(mux_c0_n265), .A2(final_w_k[26]), .ZN(c0[26]) );
  AND2_X1 mux_c0_U39 ( .A1(mux_c0_n265), .A2(final_w_k[27]), .ZN(c0[27]) );
  AND2_X1 mux_c0_U38 ( .A1(mux_c0_n264), .A2(final_w_k[28]), .ZN(c0[28]) );
  AND2_X1 mux_c0_U37 ( .A1(done), .A2(final_w_k[29]), .ZN(c0[29]) );
  AND2_X1 mux_c0_U36 ( .A1(mux_c0_n264), .A2(final_w_k[30]), .ZN(c0[30]) );
  AND2_X1 mux_c0_U35 ( .A1(mux_c0_n265), .A2(final_w_k[31]), .ZN(c0[31]) );
  AND2_X1 mux_c0_U34 ( .A1(mux_c0_n264), .A2(final_w_k[32]), .ZN(c0[32]) );
  AND2_X1 mux_c0_U33 ( .A1(mux_c0_n264), .A2(final_w_k[33]), .ZN(c0[33]) );
  AND2_X1 mux_c0_U32 ( .A1(done), .A2(final_w_k[34]), .ZN(c0[34]) );
  AND2_X1 mux_c0_U31 ( .A1(done), .A2(final_w_k[35]), .ZN(c0[35]) );
  AND2_X1 mux_c0_U30 ( .A1(done), .A2(final_w_k[36]), .ZN(c0[36]) );
  AND2_X1 mux_c0_U29 ( .A1(mux_c0_n265), .A2(final_w_k[37]), .ZN(c0[37]) );
  AND2_X1 mux_c0_U28 ( .A1(mux_c0_n264), .A2(final_w_k[38]), .ZN(c0[38]) );
  AND2_X1 mux_c0_U27 ( .A1(done), .A2(final_w_k[39]), .ZN(c0[39]) );
  AND2_X1 mux_c0_U26 ( .A1(mux_c0_n265), .A2(final_w_k[40]), .ZN(c0[40]) );
  AND2_X1 mux_c0_U25 ( .A1(mux_c0_n264), .A2(final_w_k[41]), .ZN(c0[41]) );
  AND2_X1 mux_c0_U24 ( .A1(mux_c0_n265), .A2(final_w_k[42]), .ZN(c0[42]) );
  AND2_X1 mux_c0_U23 ( .A1(mux_c0_n264), .A2(final_w_k[43]), .ZN(c0[43]) );
  AND2_X1 mux_c0_U22 ( .A1(done), .A2(final_w_k[45]), .ZN(c0[45]) );
  AND2_X1 mux_c0_U21 ( .A1(mux_c0_n265), .A2(final_w_k[46]), .ZN(c0[46]) );
  AND2_X1 mux_c0_U20 ( .A1(done), .A2(final_w_k[47]), .ZN(c0[47]) );
  AND2_X1 mux_c0_U19 ( .A1(mux_c0_n265), .A2(final_w_k[48]), .ZN(c0[48]) );
  AND2_X1 mux_c0_U18 ( .A1(mux_c0_n264), .A2(final_w_k[49]), .ZN(c0[49]) );
  AND2_X1 mux_c0_U17 ( .A1(done), .A2(final_w_k[50]), .ZN(c0[50]) );
  AND2_X1 mux_c0_U16 ( .A1(mux_c0_n264), .A2(final_w_k[51]), .ZN(c0[51]) );
  AND2_X1 mux_c0_U15 ( .A1(done), .A2(final_w_k[52]), .ZN(c0[52]) );
  AND2_X1 mux_c0_U14 ( .A1(mux_c0_n264), .A2(final_w_k[53]), .ZN(c0[53]) );
  AND2_X1 mux_c0_U13 ( .A1(done), .A2(final_w_k[54]), .ZN(c0[54]) );
  AND2_X1 mux_c0_U12 ( .A1(mux_c0_n264), .A2(final_w_k[55]), .ZN(c0[55]) );
  AND2_X1 mux_c0_U11 ( .A1(mux_c0_n264), .A2(final_w_k[56]), .ZN(c0[56]) );
  AND2_X1 mux_c0_U10 ( .A1(mux_c0_n264), .A2(final_w_k[57]), .ZN(c0[57]) );
  AND2_X1 mux_c0_U9 ( .A1(mux_c0_n264), .A2(final_w_k[58]), .ZN(c0[58]) );
  AND2_X1 mux_c0_U8 ( .A1(mux_c0_n264), .A2(final_w_k[59]), .ZN(c0[59]) );
  AND2_X1 mux_c0_U7 ( .A1(mux_c0_n264), .A2(final_w_k[60]), .ZN(c0[60]) );
  AND2_X1 mux_c0_U6 ( .A1(mux_c0_n264), .A2(final_w_k[61]), .ZN(c0[61]) );
  AND2_X1 mux_c0_U5 ( .A1(mux_c0_n264), .A2(final_w_k[62]), .ZN(c0[62]) );
  AND2_X1 mux_c0_U4 ( .A1(mux_c0_n264), .A2(final_w_k[63]), .ZN(c0[63]) );
  INV_X1 mux_c0_U3 ( .A(mux_c0_n263), .ZN(mux_c0_n264) );
  INV_X1 mux_c0_U2 ( .A(mux_c0_n263), .ZN(mux_c0_n265) );
  INV_X1 mux_c0_U1 ( .A(done), .ZN(mux_c0_n263) );
  AND2_X1 mux_c1_U67 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[56]), .ZN(
        c1[8]) );
  AND2_X1 mux_c1_U66 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[57]), .ZN(
        c1[9]) );
  AND2_X1 mux_c1_U65 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[58]), .ZN(
        c1[10]) );
  AND2_X1 mux_c1_U64 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[59]), .ZN(
        c1[11]) );
  AND2_X1 mux_c1_U63 ( .A1(done), .A2(round_inst_srout2_x[12]), .ZN(c1[12]) );
  AND2_X1 mux_c1_U62 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[13]), .ZN(
        c1[13]) );
  AND2_X1 mux_c1_U61 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[14]), .ZN(
        c1[14]) );
  AND2_X1 mux_c1_U60 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[15]), .ZN(
        c1[15]) );
  AND2_X1 mux_c1_U59 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[32]), .ZN(
        c1[16]) );
  AND2_X1 mux_c1_U58 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[33]), .ZN(
        c1[17]) );
  AND2_X1 mux_c1_U57 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[34]), .ZN(
        c1[18]) );
  AND2_X1 mux_c1_U56 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[35]), .ZN(
        c1[19]) );
  AND2_X1 mux_c1_U55 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[52]), .ZN(
        c1[20]) );
  AND2_X1 mux_c1_U54 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[53]), .ZN(
        c1[21]) );
  AND2_X1 mux_c1_U53 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[54]), .ZN(
        c1[22]) );
  AND2_X1 mux_c1_U52 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[55]), .ZN(
        c1[23]) );
  AND2_X1 mux_c1_U51 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[8]), .ZN(
        c1[24]) );
  AND2_X1 mux_c1_U50 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[9]), .ZN(
        c1[25]) );
  AND2_X1 mux_c1_U49 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[39]), .ZN(
        c1[7]) );
  AND2_X1 mux_c1_U48 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[10]), .ZN(
        c1[26]) );
  AND2_X1 mux_c1_U47 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[11]), .ZN(
        c1[27]) );
  AND2_X1 mux_c1_U46 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[28]), .ZN(
        c1[28]) );
  AND2_X1 mux_c1_U45 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[29]), .ZN(
        c1[29]) );
  AND2_X1 mux_c1_U44 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[30]), .ZN(
        c1[30]) );
  AND2_X1 mux_c1_U43 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[31]), .ZN(
        c1[31]) );
  AND2_X1 mux_c1_U42 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[48]), .ZN(
        c1[32]) );
  AND2_X1 mux_c1_U41 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[49]), .ZN(
        c1[33]) );
  AND2_X1 mux_c1_U40 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[50]), .ZN(
        c1[34]) );
  AND2_X1 mux_c1_U39 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[51]), .ZN(
        c1[35]) );
  AND2_X1 mux_c1_U38 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[4]), .ZN(
        c1[36]) );
  AND2_X1 mux_c1_U37 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[5]), .ZN(
        c1[37]) );
  AND2_X1 mux_c1_U36 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[6]), .ZN(
        c1[38]) );
  AND2_X1 mux_c1_U35 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[7]), .ZN(
        c1[39]) );
  AND2_X1 mux_c1_U34 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[24]), .ZN(
        c1[40]) );
  AND2_X1 mux_c1_U33 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[25]), .ZN(
        c1[41]) );
  AND2_X1 mux_c1_U32 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[26]), .ZN(
        c1[42]) );
  AND2_X1 mux_c1_U31 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[27]), .ZN(
        c1[43]) );
  AND2_X1 mux_c1_U30 ( .A1(done), .A2(round_inst_srout2_x[44]), .ZN(c1[44]) );
  AND2_X1 mux_c1_U29 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[45]), .ZN(
        c1[45]) );
  AND2_X1 mux_c1_U28 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[46]), .ZN(
        c1[46]) );
  AND2_X1 mux_c1_U27 ( .A1(done), .A2(round_inst_srout2_x[47]), .ZN(c1[47]) );
  AND2_X1 mux_c1_U26 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[0]), .ZN(
        c1[48]) );
  AND2_X1 mux_c1_U25 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[1]), .ZN(
        c1[49]) );
  AND2_X1 mux_c1_U24 ( .A1(done), .A2(round_inst_srout2_x[2]), .ZN(c1[50]) );
  AND2_X1 mux_c1_U23 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[3]), .ZN(
        c1[51]) );
  AND2_X1 mux_c1_U22 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[20]), .ZN(
        c1[52]) );
  AND2_X1 mux_c1_U21 ( .A1(done), .A2(round_inst_srout2_x[21]), .ZN(c1[53]) );
  AND2_X1 mux_c1_U20 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[22]), .ZN(
        c1[54]) );
  AND2_X1 mux_c1_U19 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[23]), .ZN(
        c1[55]) );
  AND2_X1 mux_c1_U18 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[40]), .ZN(
        c1[56]) );
  AND2_X1 mux_c1_U17 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[41]), .ZN(
        c1[57]) );
  AND2_X1 mux_c1_U16 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[42]), .ZN(
        c1[58]) );
  AND2_X1 mux_c1_U15 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[43]), .ZN(
        c1[59]) );
  AND2_X1 mux_c1_U14 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[60]), .ZN(
        c1[60]) );
  AND2_X1 mux_c1_U13 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[61]), .ZN(
        c1[61]) );
  AND2_X1 mux_c1_U12 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[62]), .ZN(
        c1[62]) );
  AND2_X1 mux_c1_U11 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[63]), .ZN(
        c1[63]) );
  AND2_X1 mux_c1_U10 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[38]), .ZN(
        c1[6]) );
  AND2_X1 mux_c1_U9 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[16]), .ZN(
        c1[0]) );
  AND2_X1 mux_c1_U8 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[17]), .ZN(
        c1[1]) );
  AND2_X1 mux_c1_U7 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[18]), .ZN(
        c1[2]) );
  AND2_X1 mux_c1_U6 ( .A1(mux_c1_n264), .A2(round_inst_srout2_x[19]), .ZN(
        c1[3]) );
  AND2_X1 mux_c1_U5 ( .A1(done), .A2(round_inst_srout2_x[36]), .ZN(c1[4]) );
  AND2_X1 mux_c1_U4 ( .A1(mux_c1_n265), .A2(round_inst_srout2_x[37]), .ZN(
        c1[5]) );
  INV_X1 mux_c1_U3 ( .A(mux_c1_n263), .ZN(mux_c1_n264) );
  INV_X1 mux_c1_U2 ( .A(mux_c1_n263), .ZN(mux_c1_n265) );
  INV_X1 mux_c1_U1 ( .A(done), .ZN(mux_c1_n263) );
  AND2_X1 mux_c2_U66 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[16]), .ZN(
        c2[0]) );
  AND2_X1 mux_c2_U65 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[17]), .ZN(
        c2[1]) );
  AND2_X1 mux_c2_U64 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[18]), .ZN(
        c2[2]) );
  AND2_X1 mux_c2_U63 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[19]), .ZN(
        c2[3]) );
  AND2_X1 mux_c2_U62 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[36]), .ZN(
        c2[4]) );
  AND2_X1 mux_c2_U61 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[37]), .ZN(
        c2[5]) );
  AND2_X1 mux_c2_U60 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[38]), .ZN(
        c2[6]) );
  AND2_X1 mux_c2_U59 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[39]), .ZN(
        c2[7]) );
  AND2_X1 mux_c2_U58 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[56]), .ZN(
        c2[8]) );
  AND2_X1 mux_c2_U57 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[57]), .ZN(
        c2[9]) );
  AND2_X1 mux_c2_U56 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[58]), .ZN(
        c2[10]) );
  AND2_X1 mux_c2_U55 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[59]), .ZN(
        c2[11]) );
  AND2_X1 mux_c2_U54 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[12]), .ZN(
        c2[12]) );
  AND2_X1 mux_c2_U53 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[13]), .ZN(
        c2[13]) );
  AND2_X1 mux_c2_U52 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[14]), .ZN(
        c2[14]) );
  AND2_X1 mux_c2_U51 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[15]), .ZN(
        c2[15]) );
  AND2_X1 mux_c2_U50 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[32]), .ZN(
        c2[16]) );
  AND2_X1 mux_c2_U49 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[33]), .ZN(
        c2[17]) );
  AND2_X1 mux_c2_U48 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[34]), .ZN(
        c2[18]) );
  AND2_X1 mux_c2_U47 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[35]), .ZN(
        c2[19]) );
  AND2_X1 mux_c2_U46 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[52]), .ZN(
        c2[20]) );
  AND2_X1 mux_c2_U45 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[53]), .ZN(
        c2[21]) );
  AND2_X1 mux_c2_U44 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[54]), .ZN(
        c2[22]) );
  AND2_X1 mux_c2_U43 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[55]), .ZN(
        c2[23]) );
  AND2_X1 mux_c2_U42 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[8]), .ZN(
        c2[24]) );
  AND2_X1 mux_c2_U41 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[9]), .ZN(
        c2[25]) );
  AND2_X1 mux_c2_U40 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[10]), .ZN(
        c2[26]) );
  AND2_X1 mux_c2_U39 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[11]), .ZN(
        c2[27]) );
  AND2_X1 mux_c2_U38 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[28]), .ZN(
        c2[28]) );
  AND2_X1 mux_c2_U37 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[29]), .ZN(
        c2[29]) );
  AND2_X1 mux_c2_U36 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[30]), .ZN(
        c2[30]) );
  AND2_X1 mux_c2_U35 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[31]), .ZN(
        c2[31]) );
  AND2_X1 mux_c2_U34 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[48]), .ZN(
        c2[32]) );
  AND2_X1 mux_c2_U33 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[49]), .ZN(
        c2[33]) );
  AND2_X1 mux_c2_U32 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[50]), .ZN(
        c2[34]) );
  AND2_X1 mux_c2_U31 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[51]), .ZN(
        c2[35]) );
  AND2_X1 mux_c2_U30 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[4]), .ZN(
        c2[36]) );
  AND2_X1 mux_c2_U29 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[5]), .ZN(
        c2[37]) );
  AND2_X1 mux_c2_U28 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[6]), .ZN(
        c2[38]) );
  AND2_X1 mux_c2_U27 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[7]), .ZN(
        c2[39]) );
  AND2_X1 mux_c2_U26 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[24]), .ZN(
        c2[40]) );
  AND2_X1 mux_c2_U25 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[25]), .ZN(
        c2[41]) );
  AND2_X1 mux_c2_U24 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[26]), .ZN(
        c2[42]) );
  AND2_X1 mux_c2_U23 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[27]), .ZN(
        c2[43]) );
  AND2_X1 mux_c2_U22 ( .A1(done), .A2(round_inst_srout2_y[44]), .ZN(c2[44]) );
  AND2_X1 mux_c2_U21 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[45]), .ZN(
        c2[45]) );
  AND2_X1 mux_c2_U20 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[46]), .ZN(
        c2[46]) );
  AND2_X1 mux_c2_U19 ( .A1(done), .A2(round_inst_srout2_y[47]), .ZN(c2[47]) );
  AND2_X1 mux_c2_U18 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[0]), .ZN(
        c2[48]) );
  AND2_X1 mux_c2_U17 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[1]), .ZN(
        c2[49]) );
  AND2_X1 mux_c2_U16 ( .A1(done), .A2(round_inst_srout2_y[2]), .ZN(c2[50]) );
  AND2_X1 mux_c2_U15 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[3]), .ZN(
        c2[51]) );
  AND2_X1 mux_c2_U14 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[20]), .ZN(
        c2[52]) );
  AND2_X1 mux_c2_U13 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[21]), .ZN(
        c2[53]) );
  AND2_X1 mux_c2_U12 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[22]), .ZN(
        c2[54]) );
  AND2_X1 mux_c2_U11 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[23]), .ZN(
        c2[55]) );
  AND2_X1 mux_c2_U10 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[40]), .ZN(
        c2[56]) );
  AND2_X1 mux_c2_U9 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[41]), .ZN(
        c2[57]) );
  AND2_X1 mux_c2_U8 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[42]), .ZN(
        c2[58]) );
  AND2_X1 mux_c2_U7 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[43]), .ZN(
        c2[59]) );
  AND2_X1 mux_c2_U6 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[60]), .ZN(
        c2[60]) );
  AND2_X1 mux_c2_U5 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[61]), .ZN(
        c2[61]) );
  AND2_X1 mux_c2_U4 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[62]), .ZN(
        c2[62]) );
  AND2_X1 mux_c2_U3 ( .A1(mux_c2_n264), .A2(round_inst_srout2_y[63]), .ZN(
        c2[63]) );
  INV_X2 mux_c2_U2 ( .A(mux_c2_n263), .ZN(mux_c2_n264) );
  INV_X1 mux_c2_U1 ( .A(done), .ZN(mux_c2_n263) );
  AND2_X1 mux_c3_U67 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[17]), .ZN(
        c3[1]) );
  AND2_X1 mux_c3_U66 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[18]), .ZN(
        c3[2]) );
  AND2_X1 mux_c3_U65 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[19]), .ZN(
        c3[3]) );
  AND2_X1 mux_c3_U64 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[36]), .ZN(
        c3[4]) );
  AND2_X1 mux_c3_U63 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[37]), .ZN(
        c3[5]) );
  AND2_X1 mux_c3_U62 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[38]), .ZN(
        c3[6]) );
  AND2_X1 mux_c3_U61 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[39]), .ZN(
        c3[7]) );
  AND2_X1 mux_c3_U60 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[56]), .ZN(
        c3[8]) );
  AND2_X1 mux_c3_U59 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[57]), .ZN(
        c3[9]) );
  AND2_X1 mux_c3_U58 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[58]), .ZN(
        c3[10]) );
  AND2_X1 mux_c3_U57 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[59]), .ZN(
        c3[11]) );
  AND2_X1 mux_c3_U56 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[12]), .ZN(
        c3[12]) );
  AND2_X1 mux_c3_U55 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[13]), .ZN(
        c3[13]) );
  AND2_X1 mux_c3_U54 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[14]), .ZN(
        c3[14]) );
  AND2_X1 mux_c3_U53 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[15]), .ZN(
        c3[15]) );
  AND2_X1 mux_c3_U52 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[32]), .ZN(
        c3[16]) );
  AND2_X1 mux_c3_U51 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[33]), .ZN(
        c3[17]) );
  AND2_X1 mux_c3_U50 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[34]), .ZN(
        c3[18]) );
  AND2_X1 mux_c3_U49 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[35]), .ZN(
        c3[19]) );
  AND2_X1 mux_c3_U48 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[52]), .ZN(
        c3[20]) );
  AND2_X1 mux_c3_U47 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[53]), .ZN(
        c3[21]) );
  AND2_X1 mux_c3_U46 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[54]), .ZN(
        c3[22]) );
  AND2_X1 mux_c3_U45 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[55]), .ZN(
        c3[23]) );
  AND2_X1 mux_c3_U44 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[8]), .ZN(
        c3[24]) );
  AND2_X1 mux_c3_U43 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[9]), .ZN(
        c3[25]) );
  AND2_X1 mux_c3_U42 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[10]), .ZN(
        c3[26]) );
  AND2_X1 mux_c3_U41 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[11]), .ZN(
        c3[27]) );
  AND2_X1 mux_c3_U40 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[28]), .ZN(
        c3[28]) );
  AND2_X1 mux_c3_U39 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[29]), .ZN(
        c3[29]) );
  AND2_X1 mux_c3_U38 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[30]), .ZN(
        c3[30]) );
  AND2_X1 mux_c3_U37 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[31]), .ZN(
        c3[31]) );
  AND2_X1 mux_c3_U36 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[48]), .ZN(
        c3[32]) );
  AND2_X1 mux_c3_U35 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[49]), .ZN(
        c3[33]) );
  AND2_X1 mux_c3_U34 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[50]), .ZN(
        c3[34]) );
  AND2_X1 mux_c3_U33 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[51]), .ZN(
        c3[35]) );
  AND2_X1 mux_c3_U32 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[4]), .ZN(
        c3[36]) );
  AND2_X1 mux_c3_U31 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[5]), .ZN(
        c3[37]) );
  AND2_X1 mux_c3_U30 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[6]), .ZN(
        c3[38]) );
  AND2_X1 mux_c3_U29 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[7]), .ZN(
        c3[39]) );
  AND2_X1 mux_c3_U28 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[24]), .ZN(
        c3[40]) );
  AND2_X1 mux_c3_U27 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[25]), .ZN(
        c3[41]) );
  AND2_X1 mux_c3_U26 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[26]), .ZN(
        c3[42]) );
  AND2_X1 mux_c3_U25 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[27]), .ZN(
        c3[43]) );
  AND2_X1 mux_c3_U24 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[44]), .ZN(
        c3[44]) );
  AND2_X1 mux_c3_U23 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[45]), .ZN(
        c3[45]) );
  AND2_X1 mux_c3_U22 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[46]), .ZN(
        c3[46]) );
  AND2_X1 mux_c3_U21 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[47]), .ZN(
        c3[47]) );
  AND2_X1 mux_c3_U20 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[0]), .ZN(
        c3[48]) );
  AND2_X1 mux_c3_U19 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[1]), .ZN(
        c3[49]) );
  AND2_X1 mux_c3_U18 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[2]), .ZN(
        c3[50]) );
  AND2_X1 mux_c3_U17 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[3]), .ZN(
        c3[51]) );
  AND2_X1 mux_c3_U16 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[20]), .ZN(
        c3[52]) );
  AND2_X1 mux_c3_U15 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[21]), .ZN(
        c3[53]) );
  AND2_X1 mux_c3_U14 ( .A1(mux_c3_n263), .A2(round_inst_srout2_z[22]), .ZN(
        c3[54]) );
  AND2_X1 mux_c3_U13 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[23]), .ZN(
        c3[55]) );
  AND2_X1 mux_c3_U12 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[40]), .ZN(
        c3[56]) );
  AND2_X1 mux_c3_U11 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[41]), .ZN(
        c3[57]) );
  AND2_X1 mux_c3_U10 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[42]), .ZN(
        c3[58]) );
  AND2_X1 mux_c3_U9 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[43]), .ZN(
        c3[59]) );
  AND2_X1 mux_c3_U8 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[60]), .ZN(
        c3[60]) );
  AND2_X1 mux_c3_U7 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[61]), .ZN(
        c3[61]) );
  AND2_X1 mux_c3_U6 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[62]), .ZN(
        c3[62]) );
  AND2_X1 mux_c3_U5 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[63]), .ZN(
        c3[63]) );
  AND2_X1 mux_c3_U4 ( .A1(mux_c3_n264), .A2(round_inst_srout2_z[16]), .ZN(
        c3[0]) );
  INV_X1 mux_c3_U3 ( .A(mux_c3_n262), .ZN(mux_c3_n264) );
  INV_X1 mux_c3_U2 ( .A(mux_c3_n262), .ZN(mux_c3_n263) );
  INV_X1 mux_c3_U1 ( .A(done), .ZN(mux_c3_n262) );
endmodule

