
module circuit ( clk, rst, input1, input2, key, output1, output2, Done );
  input [7:0] input1;
  input [7:0] input2;
  input [7:0] key;
  output [7:0] output1;
  output [7:0] output2;
  input clk, rst;
  output Done;
  wire   Output_Sel, done_internal, Corr_63_5_, output1_A_5_, output1_A_4_,
         output1_A_2_, output1_A_1_, ShowRcon, KeyScheduleRegisterEN,
         state_reg_hold, DoMC, DoSR, key_reg_hold, DoKeySbox,
         JustFirstColShift, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, Affine_OutInv1_n4, Affine_OutInv1_n3, Affine_OutInv1_n2,
         Affine_OutInv1_n1, OutputReg_n67, OutputReg_n66, OutputReg_n65,
         OutputReg_n64, OutputReg_n63, OutputReg_n62, OutputReg_n61,
         OutputReg_n60, OutputReg_n59, OutputReg_n58, OutputReg_n57,
         OutputReg_n56, OutputReg_n55, OutputReg_n54, OutputReg_n53,
         OutputReg_n52, OutputReg_n19, OutputReg_n18, OutputReg_n17,
         OutputReg_n51, OutputReg_n50, OutputReg_n49, OutputReg_n48,
         OutputReg_n47, OutputReg_n46, OutputReg_n45, OutputReg_n44,
         OutputReg_n43, OutputReg_n42, OutputReg_n41, OutputReg_n40,
         OutputReg_n39, OutputReg_n38, OutputReg_n37, OutputReg_n36,
         OutputReg_n35, OutputReg_n34, OutputReg_n33, OutputReg_n32,
         OutputReg_n31, OutputReg_n30, OutputReg_n29, OutputReg_n28,
         OutputReg_n27, OutputReg_n26, OutputReg_n25, OutputReg_n24,
         OutputReg_n23, OutputReg_n22, OutputReg_n21, OutputReg_n20,
         Affine_output_Inst_n12, Affine_output_Inst_n11,
         Affine_output_Inst_n10, Affine_outputC_Inst_n12,
         Affine_outputC_Inst_n11, Affine_outputC_Inst_n10,
         KeySchedule_Inst1_Affine_OutInv1_n4,
         KeySchedule_Inst1_Affine_OutInv1_n3,
         KeySchedule_Inst1_Affine_OutInv1_n2,
         KeySchedule_Inst1_Affine_OutInv1_n1, KeySchedule_Inst1_A1_n14,
         KeySchedule_Inst1_A1_n13, KeySchedule_Inst1_A1_n12,
         KeySchedule_Inst1_GEN_reg_n34, KeySchedule_Inst1_GEN_reg_n33,
         KeySchedule_Inst1_GEN_reg_n32, KeySchedule_Inst1_GEN_reg_n31,
         KeySchedule_Inst1_GEN_reg_n30, KeySchedule_Inst1_GEN_reg_n29,
         KeySchedule_Inst1_GEN_reg_n28, KeySchedule_Inst1_GEN_reg_n27,
         KeySchedule_Inst1_GEN_reg_n26, KeySchedule_Inst1_GEN_reg_n24,
         KeySchedule_Inst1_GEN_reg_n23, KeySchedule_Inst1_GEN_reg_n22,
         KeySchedule_Inst1_GEN_reg_n21, KeySchedule_Inst1_GEN_reg_n20,
         KeySchedule_Inst1_GEN_reg_n19, KeySchedule_Inst1_GEN_reg_n18,
         KeySchedule_Inst1_GEN_reg_n17, KeySchedule_Inst1_GEN_reg_n16,
         KeySchedule_Inst1_GEN_reg_n15, KeySchedule_Inst1_GEN_reg_n14,
         KeySchedule_Inst1_GEN_reg_n13, KeySchedule_Inst1_GEN_reg_n12,
         KeySchedule_Inst1_GEN_reg_n11, KeySchedule_Inst1_GEN_reg_n10,
         KeySchedule_Inst1_GEN_reg_n9, KeySchedule_Inst1_GEN_reg2_n57,
         KeySchedule_Inst1_GEN_reg2_n56, KeySchedule_Inst1_GEN_reg2_n55,
         KeySchedule_Inst1_GEN_reg2_n54, KeySchedule_Inst1_GEN_reg2_n53,
         KeySchedule_Inst1_GEN_reg2_n52, KeySchedule_Inst1_GEN_reg2_n51,
         KeySchedule_Inst1_GEN_reg2_n50, KeySchedule_Inst1_GEN_reg2_n49,
         KeySchedule_Inst1_GEN_reg2_n40, KeySchedule_Inst1_GEN_reg2_n39,
         KeySchedule_Inst1_GEN_reg2_n38, KeySchedule_Inst1_GEN_reg2_n37,
         KeySchedule_Inst1_GEN_reg2_n36, KeySchedule_Inst1_GEN_reg2_n35,
         KeySchedule_Inst1_GEN_reg2_n34, KeySchedule_Inst1_GEN_reg2_n33,
         KeySchedule_Inst1_GEN_reg2_n32, KeySchedule_Inst1_GEN_reg2_n31,
         KeySchedule_Inst1_GEN_reg2_n30, KeySchedule_Inst1_GEN_reg2_n29,
         KeySchedule_Inst1_GEN_reg2_n28, KeySchedule_Inst1_GEN_reg2_n27,
         KeySchedule_Inst1_GEN_reg2_n26, KeySchedule_Inst1_GEN_reg2_n25,
         DataPath_Registers_Inst1_n529, DataPath_Registers_Inst1_n528,
         DataPath_Registers_Inst1_n527, DataPath_Registers_Inst1_n526,
         DataPath_Registers_Inst1_n525, DataPath_Registers_Inst1_n524,
         DataPath_Registers_Inst1_n523, DataPath_Registers_Inst1_n522,
         DataPath_Registers_Inst1_n521, DataPath_Registers_Inst1_n520,
         DataPath_Registers_Inst1_n519, DataPath_Registers_Inst1_n518,
         DataPath_Registers_Inst1_n517, DataPath_Registers_Inst1_n516,
         DataPath_Registers_Inst1_n515, DataPath_Registers_Inst1_n514,
         DataPath_Registers_Inst1_n513, DataPath_Registers_Inst1_n512,
         DataPath_Registers_Inst1_n511, DataPath_Registers_Inst1_n510,
         DataPath_Registers_Inst1_n509, DataPath_Registers_Inst1_n508,
         DataPath_Registers_Inst1_n507, DataPath_Registers_Inst1_n506,
         DataPath_Registers_Inst1_n505, DataPath_Registers_Inst1_n504,
         DataPath_Registers_Inst1_n503, DataPath_Registers_Inst1_n502,
         DataPath_Registers_Inst1_n501, DataPath_Registers_Inst1_n500,
         DataPath_Registers_Inst1_n499, DataPath_Registers_Inst1_n498,
         DataPath_Registers_Inst1_n497, DataPath_Registers_Inst1_n496,
         DataPath_Registers_Inst1_n495, DataPath_Registers_Inst1_n494,
         DataPath_Registers_Inst1_n493, DataPath_Registers_Inst1_n492,
         DataPath_Registers_Inst1_n491, DataPath_Registers_Inst1_n490,
         DataPath_Registers_Inst1_n489, DataPath_Registers_Inst1_n488,
         DataPath_Registers_Inst1_n487, DataPath_Registers_Inst1_n486,
         DataPath_Registers_Inst1_n485, DataPath_Registers_Inst1_n484,
         DataPath_Registers_Inst1_n483, DataPath_Registers_Inst1_n482,
         DataPath_Registers_Inst1_n481, DataPath_Registers_Inst1_n480,
         DataPath_Registers_Inst1_n479, DataPath_Registers_Inst1_n478,
         DataPath_Registers_Inst1_n477, DataPath_Registers_Inst1_n476,
         DataPath_Registers_Inst1_n475, DataPath_Registers_Inst1_n474,
         DataPath_Registers_Inst1_n473, DataPath_Registers_Inst1_n472,
         DataPath_Registers_Inst1_n471, DataPath_Registers_Inst1_n470,
         DataPath_Registers_Inst1_n469, DataPath_Registers_Inst1_n468,
         DataPath_Registers_Inst1_n467, DataPath_Registers_Inst1_n466,
         DataPath_Registers_Inst1_n465, DataPath_Registers_Inst1_n464,
         DataPath_Registers_Inst1_n463, DataPath_Registers_Inst1_n462,
         DataPath_Registers_Inst1_n461, DataPath_Registers_Inst1_n460,
         DataPath_Registers_Inst1_n459, DataPath_Registers_Inst1_n458,
         DataPath_Registers_Inst1_n457, DataPath_Registers_Inst1_n456,
         DataPath_Registers_Inst1_n455, DataPath_Registers_Inst1_n454,
         DataPath_Registers_Inst1_n453, DataPath_Registers_Inst1_n452,
         DataPath_Registers_Inst1_n451, DataPath_Registers_Inst1_n450,
         DataPath_Registers_Inst1_n449, DataPath_Registers_Inst1_n448,
         DataPath_Registers_Inst1_n447, DataPath_Registers_Inst1_n446,
         DataPath_Registers_Inst1_n445, DataPath_Registers_Inst1_n444,
         DataPath_Registers_Inst1_n443, DataPath_Registers_Inst1_n442,
         DataPath_Registers_Inst1_n441, DataPath_Registers_Inst1_n440,
         DataPath_Registers_Inst1_n439, DataPath_Registers_Inst1_n438,
         DataPath_Registers_Inst1_n437, DataPath_Registers_Inst1_n436,
         DataPath_Registers_Inst1_n435, DataPath_Registers_Inst1_n434,
         DataPath_Registers_Inst1_n433, DataPath_Registers_Inst1_n432,
         DataPath_Registers_Inst1_n431, DataPath_Registers_Inst1_n430,
         DataPath_Registers_Inst1_n429, DataPath_Registers_Inst1_n428,
         DataPath_Registers_Inst1_n427, DataPath_Registers_Inst1_n426,
         DataPath_Registers_Inst1_n425, DataPath_Registers_Inst1_n424,
         DataPath_Registers_Inst1_n423, DataPath_Registers_Inst1_n422,
         DataPath_Registers_Inst1_n421, DataPath_Registers_Inst1_n420,
         DataPath_Registers_Inst1_n419, DataPath_Registers_Inst1_n418,
         DataPath_Registers_Inst1_n417, DataPath_Registers_Inst1_n416,
         DataPath_Registers_Inst1_n415, DataPath_Registers_Inst1_n414,
         DataPath_Registers_Inst1_n413, DataPath_Registers_Inst1_n412,
         DataPath_Registers_Inst1_n411, DataPath_Registers_Inst1_n410,
         DataPath_Registers_Inst1_n409, DataPath_Registers_Inst1_n408,
         DataPath_Registers_Inst1_n407, DataPath_Registers_Inst1_n406,
         DataPath_Registers_Inst1_n405, DataPath_Registers_Inst1_n404,
         DataPath_Registers_Inst1_n403, DataPath_Registers_Inst1_n402,
         DataPath_Registers_Inst1_n401, DataPath_Registers_Inst1_n400,
         DataPath_Registers_Inst1_n399, DataPath_Registers_Inst1_n398,
         DataPath_Registers_Inst1_n397, DataPath_Registers_Inst1_n396,
         DataPath_Registers_Inst1_n395, DataPath_Registers_Inst1_n394,
         DataPath_Registers_Inst1_n393, DataPath_Registers_Inst1_n392,
         DataPath_Registers_Inst1_n391, DataPath_Registers_Inst1_n390,
         DataPath_Registers_Inst1_n389, DataPath_Registers_Inst1_n388,
         DataPath_Registers_Inst1_n387, DataPath_Registers_Inst1_n386,
         DataPath_Registers_Inst1_n385, DataPath_Registers_Inst1_n384,
         DataPath_Registers_Inst1_n383, DataPath_Registers_Inst1_n382,
         DataPath_Registers_Inst1_n381, DataPath_Registers_Inst1_n380,
         DataPath_Registers_Inst1_n379, DataPath_Registers_Inst1_n378,
         DataPath_Registers_Inst1_n377, DataPath_Registers_Inst1_n376,
         DataPath_Registers_Inst1_n375, DataPath_Registers_Inst1_n374,
         DataPath_Registers_Inst1_n373, DataPath_Registers_Inst1_n372,
         DataPath_Registers_Inst1_n371, DataPath_Registers_Inst1_n370,
         DataPath_Registers_Inst1_n369, DataPath_Registers_Inst1_n368,
         DataPath_Registers_Inst1_n367, DataPath_Registers_Inst1_n366,
         DataPath_Registers_Inst1_n365, DataPath_Registers_Inst1_n364,
         DataPath_Registers_Inst1_n363, DataPath_Registers_Inst1_n362,
         DataPath_Registers_Inst1_n361, DataPath_Registers_Inst1_n360,
         DataPath_Registers_Inst1_n359, DataPath_Registers_Inst1_n358,
         DataPath_Registers_Inst1_n357, DataPath_Registers_Inst1_n356,
         DataPath_Registers_Inst1_n355, DataPath_Registers_Inst1_n354,
         DataPath_Registers_Inst1_n353, DataPath_Registers_Inst1_n352,
         DataPath_Registers_Inst1_n351, DataPath_Registers_Inst1_n350,
         DataPath_Registers_Inst1_n349, DataPath_Registers_Inst1_n348,
         DataPath_Registers_Inst1_n347, DataPath_Registers_Inst1_n346,
         DataPath_Registers_Inst1_n345, DataPath_Registers_Inst1_n344,
         DataPath_Registers_Inst1_n343, DataPath_Registers_Inst1_n342,
         DataPath_Registers_Inst1_n341, DataPath_Registers_Inst1_n340,
         DataPath_Registers_Inst1_n339, DataPath_Registers_Inst1_n338,
         DataPath_Registers_Inst1_n337, DataPath_Registers_Inst1_n212,
         DataPath_Registers_Inst1_n210, DataPath_Registers_Inst1_n208,
         DataPath_Registers_Inst1_n206, DataPath_Registers_Inst1_n204,
         DataPath_Registers_Inst1_n203, DataPath_Registers_Inst1_n202,
         DataPath_Registers_Inst1_n201, DataPath_Registers_Inst1_n6,
         DataPath_Registers_Inst1_n324, DataPath_Registers_Inst1_n323,
         DataPath_Registers_Inst1_n322, DataPath_Registers_Inst1_n321,
         DataPath_Registers_Inst1_n320, DataPath_Registers_Inst1_n319,
         DataPath_Registers_Inst1_n318, DataPath_Registers_Inst1_n317,
         DataPath_Registers_Inst1_n316, DataPath_Registers_Inst1_n315,
         DataPath_Registers_Inst1_n314, DataPath_Registers_Inst1_n313,
         DataPath_Registers_Inst1_n312, DataPath_Registers_Inst1_n311,
         DataPath_Registers_Inst1_n310, DataPath_Registers_Inst1_n309,
         DataPath_Registers_Inst1_n308, DataPath_Registers_Inst1_n307,
         DataPath_Registers_Inst1_n306, DataPath_Registers_Inst1_n305,
         DataPath_Registers_Inst1_n304, DataPath_Registers_Inst1_n303,
         DataPath_Registers_Inst1_n301, DataPath_Registers_Inst1_n300,
         DataPath_Registers_Inst1_n299, DataPath_Registers_Inst1_n298,
         DataPath_Registers_Inst1_n297, DataPath_Registers_Inst1_n296,
         DataPath_Registers_Inst1_n295, DataPath_Registers_Inst1_n294,
         DataPath_Registers_Inst1_n293, DataPath_Registers_Inst1_n292,
         DataPath_Registers_Inst1_n291, DataPath_Registers_Inst1_n290,
         DataPath_Registers_Inst1_n289, DataPath_Registers_Inst1_n288,
         DataPath_Registers_Inst1_n287, DataPath_Registers_Inst1_n286,
         DataPath_Registers_Inst1_n285, DataPath_Registers_Inst1_n284,
         DataPath_Registers_Inst1_n283, DataPath_Registers_Inst1_n282,
         DataPath_Registers_Inst1_n281, DataPath_Registers_Inst1_n280,
         DataPath_Registers_Inst1_n279, DataPath_Registers_Inst1_n278,
         DataPath_Registers_Inst1_n277, DataPath_Registers_Inst1_n276,
         DataPath_Registers_Inst1_n275, DataPath_Registers_Inst1_n274,
         DataPath_Registers_Inst1_n273, DataPath_Registers_Inst1_n272,
         DataPath_Registers_Inst1_n271, DataPath_Registers_Inst1_n270,
         DataPath_Registers_Inst1_n269, DataPath_Registers_Inst1_n268,
         DataPath_Registers_Inst1_n266, DataPath_Registers_Inst1_n264,
         DataPath_Registers_Inst1_n263, DataPath_Registers_Inst1_n262,
         DataPath_Registers_Inst1_n261, DataPath_Registers_Inst1_n260,
         DataPath_Registers_Inst1_n259, DataPath_Registers_Inst1_n258,
         DataPath_Registers_Inst1_n257, DataPath_Registers_Inst1_n256,
         DataPath_Registers_Inst1_n255, DataPath_Registers_Inst1_n254,
         DataPath_Registers_Inst1_n253, DataPath_Registers_Inst1_n252,
         DataPath_Registers_Inst1_n251, DataPath_Registers_Inst1_n250,
         DataPath_Registers_Inst1_n249, DataPath_Registers_Inst1_n248,
         DataPath_Registers_Inst1_n246, DataPath_Registers_Inst1_n245,
         DataPath_Registers_Inst1_n242, DataPath_Registers_Inst1_n241,
         DataPath_Registers_Inst1_n240, DataPath_Registers_Inst1_n236,
         DataPath_Registers_Inst1_n235, DataPath_Registers_Inst1_n232,
         DataPath_Registers_Inst1_n231, DataPath_Registers_Inst1_n230,
         DataPath_Registers_Inst1_n227, DataPath_Registers_Inst1_n225,
         DataPath_Registers_Inst1_n224, DataPath_Registers_Inst1_n220,
         DataPath_Registers_Inst1_n219, DataPath_Registers_Inst1_n215,
         DataPath_Registers_Inst1_in4_0_, DataPath_Registers_Inst1_in4_1_,
         DataPath_Registers_Inst1_in4_2_, DataPath_Registers_Inst1_in4_3_,
         DataPath_Registers_Inst1_in4_4_, DataPath_Registers_Inst1_in4_5_,
         DataPath_Registers_Inst1_in4_6_, DataPath_Registers_Inst1_in4_7_,
         DataPath_Registers_Inst1_in3_0_, DataPath_Registers_Inst1_in3_1_,
         DataPath_Registers_Inst1_in3_2_, DataPath_Registers_Inst1_in3_3_,
         DataPath_Registers_Inst1_in3_4_, DataPath_Registers_Inst1_in3_5_,
         DataPath_Registers_Inst1_in3_6_, DataPath_Registers_Inst1_in3_7_,
         DataPath_Registers_Inst1_in2_0_, DataPath_Registers_Inst1_in2_1_,
         DataPath_Registers_Inst1_in2_2_, DataPath_Registers_Inst1_in2_3_,
         DataPath_Registers_Inst1_in2_4_, DataPath_Registers_Inst1_in2_5_,
         DataPath_Registers_Inst1_in2_6_, DataPath_Registers_Inst1_in2_7_,
         DataPath_Registers_Inst1_in1_0_, DataPath_Registers_Inst1_in1_1_,
         DataPath_Registers_Inst1_in1_2_, DataPath_Registers_Inst1_in1_3_,
         DataPath_Registers_Inst1_in1_4_, DataPath_Registers_Inst1_in1_5_,
         DataPath_Registers_Inst1_in1_6_, DataPath_Registers_Inst1_in1_7_,
         DataPath_Registers_Inst1_S12_0_, DataPath_Registers_Inst1_S12_1_,
         DataPath_Registers_Inst1_S12_2_, DataPath_Registers_Inst1_S12_3_,
         DataPath_Registers_Inst1_S12_4_, DataPath_Registers_Inst1_S12_5_,
         DataPath_Registers_Inst1_S12_6_, DataPath_Registers_Inst1_S12_7_,
         DataPath_Registers_Inst1_S14_0_, DataPath_Registers_Inst1_S14_1_,
         DataPath_Registers_Inst1_S14_2_, DataPath_Registers_Inst1_S14_3_,
         DataPath_Registers_Inst1_S14_4_, DataPath_Registers_Inst1_S14_5_,
         DataPath_Registers_Inst1_S14_6_, DataPath_Registers_Inst1_S14_7_,
         DataPath_Registers_Inst1_S8_0_, DataPath_Registers_Inst1_S8_1_,
         DataPath_Registers_Inst1_S8_2_, DataPath_Registers_Inst1_S8_3_,
         DataPath_Registers_Inst1_S8_4_, DataPath_Registers_Inst1_S8_5_,
         DataPath_Registers_Inst1_S8_6_, DataPath_Registers_Inst1_S8_7_,
         DataPath_Registers_Inst1_S15_0_, DataPath_Registers_Inst1_S15_1_,
         DataPath_Registers_Inst1_S15_2_, DataPath_Registers_Inst1_S15_3_,
         DataPath_Registers_Inst1_S15_4_, DataPath_Registers_Inst1_S15_5_,
         DataPath_Registers_Inst1_S15_6_, DataPath_Registers_Inst1_S15_7_,
         DataPath_Registers_Inst1_S7_0_, DataPath_Registers_Inst1_S7_1_,
         DataPath_Registers_Inst1_S7_2_, DataPath_Registers_Inst1_S7_3_,
         DataPath_Registers_Inst1_S7_4_, DataPath_Registers_Inst1_S7_5_,
         DataPath_Registers_Inst1_S7_6_, DataPath_Registers_Inst1_S7_7_,
         DataPath_Registers_Inst1_S10_0_, DataPath_Registers_Inst1_S10_1_,
         DataPath_Registers_Inst1_S10_2_, DataPath_Registers_Inst1_S10_3_,
         DataPath_Registers_Inst1_S10_4_, DataPath_Registers_Inst1_S10_5_,
         DataPath_Registers_Inst1_S10_6_, DataPath_Registers_Inst1_S10_7_,
         DataPath_Registers_Inst1_S11_0_, DataPath_Registers_Inst1_S11_1_,
         DataPath_Registers_Inst1_S11_2_, DataPath_Registers_Inst1_S11_3_,
         DataPath_Registers_Inst1_S11_4_, DataPath_Registers_Inst1_S11_5_,
         DataPath_Registers_Inst1_S11_6_, DataPath_Registers_Inst1_S11_7_,
         DataPath_Registers_Inst1_S6_0_, DataPath_Registers_Inst1_S6_1_,
         DataPath_Registers_Inst1_S6_2_, DataPath_Registers_Inst1_S6_3_,
         DataPath_Registers_Inst1_S6_4_, DataPath_Registers_Inst1_S6_5_,
         DataPath_Registers_Inst1_S6_6_, DataPath_Registers_Inst1_S6_7_,
         DataPath_Registers_Inst1_S4_0_, DataPath_Registers_Inst1_S4_1_,
         DataPath_Registers_Inst1_S4_2_, DataPath_Registers_Inst1_S4_3_,
         DataPath_Registers_Inst1_S4_4_, DataPath_Registers_Inst1_S4_5_,
         DataPath_Registers_Inst1_S4_6_, DataPath_Registers_Inst1_S4_7_,
         DataPath_Registers_Inst1_S3_0_, DataPath_Registers_Inst1_S3_1_,
         DataPath_Registers_Inst1_S3_2_, DataPath_Registers_Inst1_S3_3_,
         DataPath_Registers_Inst1_S3_4_, DataPath_Registers_Inst1_S3_5_,
         DataPath_Registers_Inst1_S3_6_, DataPath_Registers_Inst1_S3_7_,
         DataPath_Registers_Inst1_S2_0_, DataPath_Registers_Inst1_S2_1_,
         DataPath_Registers_Inst1_S2_2_, DataPath_Registers_Inst1_S2_3_,
         DataPath_Registers_Inst1_S2_4_, DataPath_Registers_Inst1_S2_5_,
         DataPath_Registers_Inst1_S2_6_, DataPath_Registers_Inst1_S2_7_,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n10,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n9,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n7,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n6,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n11,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n10,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n8,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n7,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n10,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n9,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n7,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n6,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n10,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n9,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n7,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n6,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n10,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n9,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n7,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n6,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n10,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n9,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n7,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n6,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n10,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n9,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n7,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n6,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n10,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n9,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n7,
         DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n6,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n12,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n11,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n10,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n8,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n7,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n12,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n11,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n10,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n8,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n7,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n12,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n11,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n10,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n8,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n7,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n12,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n11,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n10,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n8,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n7,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n12,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n11,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n10,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n8,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n7,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n12,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n11,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n10,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n8,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n7,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n12,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n11,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n10,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n8,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n7,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n12,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n11,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n10,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n8,
         DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n7,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n12,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n11,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n10,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n8,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n7,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n12,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n11,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n10,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n8,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n7,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n12,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n11,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n10,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n8,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n7,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n11,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n10,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n8,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n7,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n11,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n10,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n9,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n7,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n6,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n11,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n10,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n9,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n7,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n6,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n11,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n10,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n9,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n7,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n6,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n11,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n10,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n9,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n7,
         DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n6,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n12,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n11,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n10,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n8,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n7,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n12,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n11,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n10,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n8,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n7,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n12,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n11,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n10,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n8,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n7,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n12,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n11,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n10,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n8,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n7,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n12,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n11,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n10,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n8,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n7,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n12,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n11,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n10,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n8,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n7,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n12,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n11,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n10,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n8,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n7,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n12,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n11,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n10,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n8,
         DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n7,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n11,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n10,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n8,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n7,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n11,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n10,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n8,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n7,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n11,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n10,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n8,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n7,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n11,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n10,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n8,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n7,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n11,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n10,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n8,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n7,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n11,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n10,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n9,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n7,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n6,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n11,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n10,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n9,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n7,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n6,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n11,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n10,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n9,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n7,
         DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n6,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n12,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n11,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n10,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n8,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n7,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n12,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n11,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n10,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n8,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n7,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n12,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n11,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n10,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n8,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n7,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n12,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n11,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n10,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n8,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n7,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n12,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n11,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n10,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n8,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n7,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n12,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n11,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n10,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n8,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n7,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n12,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n11,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n10,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n8,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n7,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n12,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n11,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n10,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n8,
         DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n7,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n12,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n11,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n10,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n8,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n7,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n12,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n11,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n10,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n8,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n7,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n11,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n10,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n8,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n7,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n11,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n10,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n8,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n7,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n11,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n10,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n8,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n7,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n11,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n10,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n9,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n7,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n6,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n11,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n10,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n9,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n7,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n6,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n11,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n10,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n9,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n7,
         DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n6,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n11,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n10,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n8,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n7,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n11,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n10,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n8,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n7,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n11,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n10,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n8,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n7,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n11,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n10,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n8,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n7,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n11,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n10,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n8,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n7,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n11,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n10,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n8,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n7,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n11,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n10,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n8,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n7,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n11,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n10,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n8,
         DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n7,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n11,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n10,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n8,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n7,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n11,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n10,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n8,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n7,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n11,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n10,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n8,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n7,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n11,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n10,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n8,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n7,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n11,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n10,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n8,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n7,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n11,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n10,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n9,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n7,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n6,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n11,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n10,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n9,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n7,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n6,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n11,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n10,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n9,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n7,
         DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n6,
         DataPath_Registers_Inst1_GEN_reg1_n134,
         DataPath_Registers_Inst1_GEN_reg1_n133,
         DataPath_Registers_Inst1_GEN_reg1_n132,
         DataPath_Registers_Inst1_GEN_reg1_n131,
         DataPath_Registers_Inst1_GEN_reg1_n130,
         DataPath_Registers_Inst1_GEN_reg1_n129,
         DataPath_Registers_Inst1_GEN_reg1_n128,
         DataPath_Registers_Inst1_GEN_reg1_n127,
         DataPath_Registers_Inst1_GEN_reg1_n126,
         DataPath_Registers_Inst1_GEN_reg1_n125,
         DataPath_Registers_Inst1_GEN_reg1_n124,
         DataPath_Registers_Inst1_GEN_reg1_n123,
         DataPath_Registers_Inst1_GEN_reg1_n122,
         DataPath_Registers_Inst1_GEN_reg1_n121,
         DataPath_Registers_Inst1_GEN_reg1_n120,
         DataPath_Registers_Inst1_GEN_reg1_n119,
         DataPath_Registers_Inst1_GEN_reg1_n118,
         DataPath_Registers_Inst1_GEN_reg1_n117,
         DataPath_Registers_Inst1_GEN_reg1_n116,
         DataPath_Registers_Inst1_GEN_reg1_n115,
         DataPath_Registers_Inst1_GEN_reg1_n114,
         DataPath_Registers_Inst1_GEN_reg1_n113,
         DataPath_Registers_Inst1_GEN_reg1_n112,
         DataPath_Registers_Inst1_GEN_reg1_n111,
         DataPath_Registers_Inst1_GEN_reg1_n110,
         DataPath_Registers_Inst1_GEN_reg1_n109,
         DataPath_Registers_Inst1_GEN_reg1_n108,
         DataPath_Registers_Inst1_GEN_reg1_n107,
         DataPath_Registers_Inst1_GEN_reg1_n106,
         DataPath_Registers_Inst1_GEN_reg1_n105,
         DataPath_Registers_Inst1_GEN_reg1_n104,
         DataPath_Registers_Inst1_GEN_reg1_n103,
         DataPath_Registers_Inst1_GEN_reg1_n102,
         DataPath_Registers_Inst1_GEN_reg1_n101,
         DataPath_Registers_Inst1_GEN_reg1_n100,
         DataPath_Registers_Inst1_GEN_reg1_n96,
         DataPath_Registers_Inst1_GEN_reg1_n95,
         DataPath_Registers_Inst1_GEN_reg1_n94,
         DataPath_Registers_Inst1_GEN_reg1_n93,
         DataPath_Registers_Inst1_GEN_reg1_n92,
         DataPath_Registers_Inst1_GEN_reg1_n91,
         DataPath_Registers_Inst1_GEN_reg1_n90,
         DataPath_Registers_Inst1_GEN_reg1_n89,
         DataPath_Registers_Inst1_GEN_reg1_n88,
         DataPath_Registers_Inst1_GEN_reg1_n87,
         DataPath_Registers_Inst1_GEN_reg1_n86,
         DataPath_Registers_Inst1_GEN_reg1_n85,
         DataPath_Registers_Inst1_GEN_reg1_n84,
         DataPath_Registers_Inst1_GEN_reg1_n83,
         DataPath_Registers_Inst1_GEN_reg1_n82,
         DataPath_Registers_Inst1_GEN_reg1_n81,
         DataPath_Registers_Inst1_GEN_reg1_n80,
         DataPath_Registers_Inst1_GEN_reg1_n79,
         DataPath_Registers_Inst1_GEN_reg1_n78,
         DataPath_Registers_Inst1_GEN_reg1_n77,
         DataPath_Registers_Inst1_GEN_reg1_n76,
         DataPath_Registers_Inst1_GEN_reg1_n75,
         DataPath_Registers_Inst1_GEN_reg1_n74,
         DataPath_Registers_Inst1_GEN_reg1_n73,
         DataPath_Registers_Inst1_GEN_reg1_n72,
         DataPath_Registers_Inst1_GEN_reg1_n71,
         DataPath_Registers_Inst1_GEN_reg1_n70,
         DataPath_Registers_Inst1_GEN_reg1_n69,
         DataPath_Registers_Inst1_GEN_reg1_n68,
         DataPath_Registers_Inst1_GEN_reg1_n67,
         DataPath_Registers_Inst1_GEN_reg1_n66,
         DataPath_Registers_Inst1_GEN_reg1_n65,
         DataPath_Registers_Inst1_GEN_reg1_n64,
         DataPath_Registers_Inst1_GEN_reg1_n63,
         DataPath_Registers_Inst1_GEN_reg1_n62,
         DataPath_Registers_Inst1_GEN_reg1_n61,
         DataPath_Registers_Inst1_GEN_reg1_n60,
         DataPath_Registers_Inst1_GEN_reg1_n59,
         DataPath_Registers_Inst1_GEN_reg1_n58,
         DataPath_Registers_Inst1_GEN_reg1_n57,
         DataPath_Registers_Inst1_GEN_reg1_n56,
         DataPath_Registers_Inst1_GEN_reg1_n55,
         DataPath_Registers_Inst1_GEN_reg1_n54,
         DataPath_Registers_Inst1_GEN_reg1_n53,
         DataPath_Registers_Inst1_GEN_reg1_n52,
         DataPath_Registers_Inst1_GEN_reg1_n51,
         DataPath_Registers_Inst1_GEN_reg1_n50,
         DataPath_Registers_Inst1_GEN_reg1_n49,
         DataPath_Registers_Inst1_GEN_reg1_n48,
         DataPath_Registers_Inst1_GEN_reg1_n47,
         DataPath_Registers_Inst1_GEN_reg1_n46,
         DataPath_Registers_Inst1_GEN_reg1_n45,
         DataPath_Registers_Inst1_GEN_reg1_n44,
         DataPath_Registers_Inst1_GEN_reg1_n43,
         DataPath_Registers_Inst1_GEN_reg1_n42,
         DataPath_Registers_Inst1_GEN_reg1_n41,
         DataPath_Registers_Inst1_GEN_reg1_n40,
         DataPath_Registers_Inst1_GEN_reg1_n39,
         DataPath_Registers_Inst1_GEN_reg1_n38,
         DataPath_Registers_Inst1_GEN_reg1_n37,
         DataPath_Registers_Inst1_GEN_reg1_n36,
         DataPath_Registers_Inst1_GEN_reg1_n35,
         DataPath_Registers_Inst1_GEN_reg1_n34,
         DataPath_Registers_Inst1_GEN_reg1_n33,
         DataPath_Registers_Inst1_A1_n14, DataPath_Registers_Inst1_A1_n13,
         DataPath_Registers_Inst1_A1_n12, DataPath_Registers_Inst1_A2_n14,
         DataPath_Registers_Inst1_A2_n13, DataPath_Registers_Inst1_A2_n12,
         DataPath_Registers_Inst1_A3_n14, DataPath_Registers_Inst1_A3_n13,
         DataPath_Registers_Inst1_A3_n12, DataPath_Registers_Inst1_A4_n14,
         DataPath_Registers_Inst1_A4_n13, DataPath_Registers_Inst1_A4_n12,
         DataPath_Registers_Inst2_n529, DataPath_Registers_Inst2_n528,
         DataPath_Registers_Inst2_n527, DataPath_Registers_Inst2_n526,
         DataPath_Registers_Inst2_n525, DataPath_Registers_Inst2_n524,
         DataPath_Registers_Inst2_n523, DataPath_Registers_Inst2_n522,
         DataPath_Registers_Inst2_n521, DataPath_Registers_Inst2_n520,
         DataPath_Registers_Inst2_n519, DataPath_Registers_Inst2_n518,
         DataPath_Registers_Inst2_n517, DataPath_Registers_Inst2_n516,
         DataPath_Registers_Inst2_n515, DataPath_Registers_Inst2_n514,
         DataPath_Registers_Inst2_n513, DataPath_Registers_Inst2_n512,
         DataPath_Registers_Inst2_n511, DataPath_Registers_Inst2_n510,
         DataPath_Registers_Inst2_n509, DataPath_Registers_Inst2_n508,
         DataPath_Registers_Inst2_n507, DataPath_Registers_Inst2_n506,
         DataPath_Registers_Inst2_n505, DataPath_Registers_Inst2_n504,
         DataPath_Registers_Inst2_n503, DataPath_Registers_Inst2_n502,
         DataPath_Registers_Inst2_n501, DataPath_Registers_Inst2_n500,
         DataPath_Registers_Inst2_n499, DataPath_Registers_Inst2_n498,
         DataPath_Registers_Inst2_n497, DataPath_Registers_Inst2_n496,
         DataPath_Registers_Inst2_n495, DataPath_Registers_Inst2_n494,
         DataPath_Registers_Inst2_n493, DataPath_Registers_Inst2_n492,
         DataPath_Registers_Inst2_n491, DataPath_Registers_Inst2_n490,
         DataPath_Registers_Inst2_n489, DataPath_Registers_Inst2_n488,
         DataPath_Registers_Inst2_n487, DataPath_Registers_Inst2_n486,
         DataPath_Registers_Inst2_n485, DataPath_Registers_Inst2_n484,
         DataPath_Registers_Inst2_n483, DataPath_Registers_Inst2_n482,
         DataPath_Registers_Inst2_n481, DataPath_Registers_Inst2_n480,
         DataPath_Registers_Inst2_n479, DataPath_Registers_Inst2_n478,
         DataPath_Registers_Inst2_n477, DataPath_Registers_Inst2_n476,
         DataPath_Registers_Inst2_n475, DataPath_Registers_Inst2_n474,
         DataPath_Registers_Inst2_n473, DataPath_Registers_Inst2_n472,
         DataPath_Registers_Inst2_n471, DataPath_Registers_Inst2_n470,
         DataPath_Registers_Inst2_n469, DataPath_Registers_Inst2_n468,
         DataPath_Registers_Inst2_n467, DataPath_Registers_Inst2_n466,
         DataPath_Registers_Inst2_n465, DataPath_Registers_Inst2_n464,
         DataPath_Registers_Inst2_n463, DataPath_Registers_Inst2_n462,
         DataPath_Registers_Inst2_n461, DataPath_Registers_Inst2_n460,
         DataPath_Registers_Inst2_n459, DataPath_Registers_Inst2_n458,
         DataPath_Registers_Inst2_n457, DataPath_Registers_Inst2_n456,
         DataPath_Registers_Inst2_n455, DataPath_Registers_Inst2_n454,
         DataPath_Registers_Inst2_n453, DataPath_Registers_Inst2_n452,
         DataPath_Registers_Inst2_n451, DataPath_Registers_Inst2_n450,
         DataPath_Registers_Inst2_n449, DataPath_Registers_Inst2_n448,
         DataPath_Registers_Inst2_n447, DataPath_Registers_Inst2_n446,
         DataPath_Registers_Inst2_n445, DataPath_Registers_Inst2_n444,
         DataPath_Registers_Inst2_n443, DataPath_Registers_Inst2_n442,
         DataPath_Registers_Inst2_n441, DataPath_Registers_Inst2_n440,
         DataPath_Registers_Inst2_n439, DataPath_Registers_Inst2_n438,
         DataPath_Registers_Inst2_n437, DataPath_Registers_Inst2_n436,
         DataPath_Registers_Inst2_n435, DataPath_Registers_Inst2_n434,
         DataPath_Registers_Inst2_n433, DataPath_Registers_Inst2_n432,
         DataPath_Registers_Inst2_n431, DataPath_Registers_Inst2_n430,
         DataPath_Registers_Inst2_n429, DataPath_Registers_Inst2_n428,
         DataPath_Registers_Inst2_n427, DataPath_Registers_Inst2_n426,
         DataPath_Registers_Inst2_n425, DataPath_Registers_Inst2_n424,
         DataPath_Registers_Inst2_n423, DataPath_Registers_Inst2_n422,
         DataPath_Registers_Inst2_n421, DataPath_Registers_Inst2_n420,
         DataPath_Registers_Inst2_n419, DataPath_Registers_Inst2_n418,
         DataPath_Registers_Inst2_n417, DataPath_Registers_Inst2_n416,
         DataPath_Registers_Inst2_n415, DataPath_Registers_Inst2_n414,
         DataPath_Registers_Inst2_n413, DataPath_Registers_Inst2_n412,
         DataPath_Registers_Inst2_n411, DataPath_Registers_Inst2_n410,
         DataPath_Registers_Inst2_n409, DataPath_Registers_Inst2_n408,
         DataPath_Registers_Inst2_n407, DataPath_Registers_Inst2_n406,
         DataPath_Registers_Inst2_n405, DataPath_Registers_Inst2_n404,
         DataPath_Registers_Inst2_n403, DataPath_Registers_Inst2_n402,
         DataPath_Registers_Inst2_n401, DataPath_Registers_Inst2_n400,
         DataPath_Registers_Inst2_n399, DataPath_Registers_Inst2_n398,
         DataPath_Registers_Inst2_n397, DataPath_Registers_Inst2_n396,
         DataPath_Registers_Inst2_n395, DataPath_Registers_Inst2_n394,
         DataPath_Registers_Inst2_n393, DataPath_Registers_Inst2_n392,
         DataPath_Registers_Inst2_n391, DataPath_Registers_Inst2_n390,
         DataPath_Registers_Inst2_n389, DataPath_Registers_Inst2_n388,
         DataPath_Registers_Inst2_n387, DataPath_Registers_Inst2_n386,
         DataPath_Registers_Inst2_n385, DataPath_Registers_Inst2_n384,
         DataPath_Registers_Inst2_n383, DataPath_Registers_Inst2_n382,
         DataPath_Registers_Inst2_n381, DataPath_Registers_Inst2_n380,
         DataPath_Registers_Inst2_n379, DataPath_Registers_Inst2_n378,
         DataPath_Registers_Inst2_n377, DataPath_Registers_Inst2_n376,
         DataPath_Registers_Inst2_n375, DataPath_Registers_Inst2_n374,
         DataPath_Registers_Inst2_n373, DataPath_Registers_Inst2_n372,
         DataPath_Registers_Inst2_n371, DataPath_Registers_Inst2_n370,
         DataPath_Registers_Inst2_n369, DataPath_Registers_Inst2_n368,
         DataPath_Registers_Inst2_n367, DataPath_Registers_Inst2_n366,
         DataPath_Registers_Inst2_n365, DataPath_Registers_Inst2_n364,
         DataPath_Registers_Inst2_n363, DataPath_Registers_Inst2_n362,
         DataPath_Registers_Inst2_n361, DataPath_Registers_Inst2_n360,
         DataPath_Registers_Inst2_n359, DataPath_Registers_Inst2_n358,
         DataPath_Registers_Inst2_n357, DataPath_Registers_Inst2_n356,
         DataPath_Registers_Inst2_n355, DataPath_Registers_Inst2_n354,
         DataPath_Registers_Inst2_n353, DataPath_Registers_Inst2_n352,
         DataPath_Registers_Inst2_n351, DataPath_Registers_Inst2_n350,
         DataPath_Registers_Inst2_n349, DataPath_Registers_Inst2_n348,
         DataPath_Registers_Inst2_n347, DataPath_Registers_Inst2_n346,
         DataPath_Registers_Inst2_n345, DataPath_Registers_Inst2_n344,
         DataPath_Registers_Inst2_n343, DataPath_Registers_Inst2_n342,
         DataPath_Registers_Inst2_n341, DataPath_Registers_Inst2_n340,
         DataPath_Registers_Inst2_n339, DataPath_Registers_Inst2_n338,
         DataPath_Registers_Inst2_n337, DataPath_Registers_Inst2_n212,
         DataPath_Registers_Inst2_n210, DataPath_Registers_Inst2_n208,
         DataPath_Registers_Inst2_n206, DataPath_Registers_Inst2_n204,
         DataPath_Registers_Inst2_n203, DataPath_Registers_Inst2_n202,
         DataPath_Registers_Inst2_n201, DataPath_Registers_Inst2_n6,
         DataPath_Registers_Inst2_n324, DataPath_Registers_Inst2_n323,
         DataPath_Registers_Inst2_n322, DataPath_Registers_Inst2_n321,
         DataPath_Registers_Inst2_n320, DataPath_Registers_Inst2_n319,
         DataPath_Registers_Inst2_n318, DataPath_Registers_Inst2_n317,
         DataPath_Registers_Inst2_n316, DataPath_Registers_Inst2_n315,
         DataPath_Registers_Inst2_n314, DataPath_Registers_Inst2_n313,
         DataPath_Registers_Inst2_n312, DataPath_Registers_Inst2_n311,
         DataPath_Registers_Inst2_n310, DataPath_Registers_Inst2_n309,
         DataPath_Registers_Inst2_n308, DataPath_Registers_Inst2_n307,
         DataPath_Registers_Inst2_n306, DataPath_Registers_Inst2_n305,
         DataPath_Registers_Inst2_n304, DataPath_Registers_Inst2_n303,
         DataPath_Registers_Inst2_n301, DataPath_Registers_Inst2_n300,
         DataPath_Registers_Inst2_n299, DataPath_Registers_Inst2_n298,
         DataPath_Registers_Inst2_n297, DataPath_Registers_Inst2_n296,
         DataPath_Registers_Inst2_n295, DataPath_Registers_Inst2_n294,
         DataPath_Registers_Inst2_n293, DataPath_Registers_Inst2_n292,
         DataPath_Registers_Inst2_n291, DataPath_Registers_Inst2_n290,
         DataPath_Registers_Inst2_n289, DataPath_Registers_Inst2_n288,
         DataPath_Registers_Inst2_n287, DataPath_Registers_Inst2_n286,
         DataPath_Registers_Inst2_n285, DataPath_Registers_Inst2_n284,
         DataPath_Registers_Inst2_n283, DataPath_Registers_Inst2_n282,
         DataPath_Registers_Inst2_n281, DataPath_Registers_Inst2_n280,
         DataPath_Registers_Inst2_n279, DataPath_Registers_Inst2_n278,
         DataPath_Registers_Inst2_n277, DataPath_Registers_Inst2_n276,
         DataPath_Registers_Inst2_n275, DataPath_Registers_Inst2_n274,
         DataPath_Registers_Inst2_n273, DataPath_Registers_Inst2_n272,
         DataPath_Registers_Inst2_n271, DataPath_Registers_Inst2_n270,
         DataPath_Registers_Inst2_n269, DataPath_Registers_Inst2_n268,
         DataPath_Registers_Inst2_n266, DataPath_Registers_Inst2_n264,
         DataPath_Registers_Inst2_n263, DataPath_Registers_Inst2_n262,
         DataPath_Registers_Inst2_n261, DataPath_Registers_Inst2_n260,
         DataPath_Registers_Inst2_n259, DataPath_Registers_Inst2_n258,
         DataPath_Registers_Inst2_n257, DataPath_Registers_Inst2_n256,
         DataPath_Registers_Inst2_n255, DataPath_Registers_Inst2_n254,
         DataPath_Registers_Inst2_n253, DataPath_Registers_Inst2_n252,
         DataPath_Registers_Inst2_n251, DataPath_Registers_Inst2_n250,
         DataPath_Registers_Inst2_n249, DataPath_Registers_Inst2_n248,
         DataPath_Registers_Inst2_n246, DataPath_Registers_Inst2_n245,
         DataPath_Registers_Inst2_n242, DataPath_Registers_Inst2_n241,
         DataPath_Registers_Inst2_n240, DataPath_Registers_Inst2_n236,
         DataPath_Registers_Inst2_n235, DataPath_Registers_Inst2_n232,
         DataPath_Registers_Inst2_n231, DataPath_Registers_Inst2_n230,
         DataPath_Registers_Inst2_n227, DataPath_Registers_Inst2_n225,
         DataPath_Registers_Inst2_n224, DataPath_Registers_Inst2_n220,
         DataPath_Registers_Inst2_n219, DataPath_Registers_Inst2_n215,
         DataPath_Registers_Inst2_in4_0_, DataPath_Registers_Inst2_in4_1_,
         DataPath_Registers_Inst2_in4_2_, DataPath_Registers_Inst2_in4_3_,
         DataPath_Registers_Inst2_in4_4_, DataPath_Registers_Inst2_in4_5_,
         DataPath_Registers_Inst2_in4_6_, DataPath_Registers_Inst2_in4_7_,
         DataPath_Registers_Inst2_in3_0_, DataPath_Registers_Inst2_in3_1_,
         DataPath_Registers_Inst2_in3_2_, DataPath_Registers_Inst2_in3_3_,
         DataPath_Registers_Inst2_in3_4_, DataPath_Registers_Inst2_in3_5_,
         DataPath_Registers_Inst2_in3_6_, DataPath_Registers_Inst2_in3_7_,
         DataPath_Registers_Inst2_in2_0_, DataPath_Registers_Inst2_in2_1_,
         DataPath_Registers_Inst2_in2_2_, DataPath_Registers_Inst2_in2_3_,
         DataPath_Registers_Inst2_in2_4_, DataPath_Registers_Inst2_in2_5_,
         DataPath_Registers_Inst2_in2_6_, DataPath_Registers_Inst2_in2_7_,
         DataPath_Registers_Inst2_in1_0_, DataPath_Registers_Inst2_in1_1_,
         DataPath_Registers_Inst2_in1_2_, DataPath_Registers_Inst2_in1_3_,
         DataPath_Registers_Inst2_in1_4_, DataPath_Registers_Inst2_in1_5_,
         DataPath_Registers_Inst2_in1_6_, DataPath_Registers_Inst2_in1_7_,
         DataPath_Registers_Inst2_S12_0_, DataPath_Registers_Inst2_S12_1_,
         DataPath_Registers_Inst2_S12_2_, DataPath_Registers_Inst2_S12_3_,
         DataPath_Registers_Inst2_S12_4_, DataPath_Registers_Inst2_S12_5_,
         DataPath_Registers_Inst2_S12_6_, DataPath_Registers_Inst2_S12_7_,
         DataPath_Registers_Inst2_S14_0_, DataPath_Registers_Inst2_S14_1_,
         DataPath_Registers_Inst2_S14_2_, DataPath_Registers_Inst2_S14_3_,
         DataPath_Registers_Inst2_S14_4_, DataPath_Registers_Inst2_S14_5_,
         DataPath_Registers_Inst2_S14_6_, DataPath_Registers_Inst2_S14_7_,
         DataPath_Registers_Inst2_S8_0_, DataPath_Registers_Inst2_S8_1_,
         DataPath_Registers_Inst2_S8_2_, DataPath_Registers_Inst2_S8_3_,
         DataPath_Registers_Inst2_S8_4_, DataPath_Registers_Inst2_S8_5_,
         DataPath_Registers_Inst2_S8_6_, DataPath_Registers_Inst2_S8_7_,
         DataPath_Registers_Inst2_S15_0_, DataPath_Registers_Inst2_S15_1_,
         DataPath_Registers_Inst2_S15_2_, DataPath_Registers_Inst2_S15_3_,
         DataPath_Registers_Inst2_S15_4_, DataPath_Registers_Inst2_S15_5_,
         DataPath_Registers_Inst2_S15_6_, DataPath_Registers_Inst2_S15_7_,
         DataPath_Registers_Inst2_S7_0_, DataPath_Registers_Inst2_S7_1_,
         DataPath_Registers_Inst2_S7_2_, DataPath_Registers_Inst2_S7_3_,
         DataPath_Registers_Inst2_S7_4_, DataPath_Registers_Inst2_S7_5_,
         DataPath_Registers_Inst2_S7_6_, DataPath_Registers_Inst2_S7_7_,
         DataPath_Registers_Inst2_S10_0_, DataPath_Registers_Inst2_S10_1_,
         DataPath_Registers_Inst2_S10_2_, DataPath_Registers_Inst2_S10_3_,
         DataPath_Registers_Inst2_S10_4_, DataPath_Registers_Inst2_S10_5_,
         DataPath_Registers_Inst2_S10_6_, DataPath_Registers_Inst2_S10_7_,
         DataPath_Registers_Inst2_S11_0_, DataPath_Registers_Inst2_S11_1_,
         DataPath_Registers_Inst2_S11_2_, DataPath_Registers_Inst2_S11_3_,
         DataPath_Registers_Inst2_S11_4_, DataPath_Registers_Inst2_S11_5_,
         DataPath_Registers_Inst2_S11_6_, DataPath_Registers_Inst2_S11_7_,
         DataPath_Registers_Inst2_S6_0_, DataPath_Registers_Inst2_S6_1_,
         DataPath_Registers_Inst2_S6_2_, DataPath_Registers_Inst2_S6_3_,
         DataPath_Registers_Inst2_S6_4_, DataPath_Registers_Inst2_S6_5_,
         DataPath_Registers_Inst2_S6_6_, DataPath_Registers_Inst2_S6_7_,
         DataPath_Registers_Inst2_S4_0_, DataPath_Registers_Inst2_S4_1_,
         DataPath_Registers_Inst2_S4_2_, DataPath_Registers_Inst2_S4_3_,
         DataPath_Registers_Inst2_S4_4_, DataPath_Registers_Inst2_S4_5_,
         DataPath_Registers_Inst2_S4_6_, DataPath_Registers_Inst2_S4_7_,
         DataPath_Registers_Inst2_S3_0_, DataPath_Registers_Inst2_S3_1_,
         DataPath_Registers_Inst2_S3_2_, DataPath_Registers_Inst2_S3_3_,
         DataPath_Registers_Inst2_S3_4_, DataPath_Registers_Inst2_S3_5_,
         DataPath_Registers_Inst2_S3_6_, DataPath_Registers_Inst2_S3_7_,
         DataPath_Registers_Inst2_S2_0_, DataPath_Registers_Inst2_S2_1_,
         DataPath_Registers_Inst2_S2_2_, DataPath_Registers_Inst2_S2_3_,
         DataPath_Registers_Inst2_S2_4_, DataPath_Registers_Inst2_S2_5_,
         DataPath_Registers_Inst2_S2_6_, DataPath_Registers_Inst2_S2_7_,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n12,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n11,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n10,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n8,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n7,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n12,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n11,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n10,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n8,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n7,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n12,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n11,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n10,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n8,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n7,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n12,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n11,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n10,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n8,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n7,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n12,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n11,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n10,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n8,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n7,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n12,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n11,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n10,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n8,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n7,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n12,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n11,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n10,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n8,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n7,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n12,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n11,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n10,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n8,
         DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n7,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n12,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n11,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n10,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n8,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n7,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n12,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n11,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n10,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n8,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n7,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n12,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n11,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n10,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n8,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n7,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n12,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n11,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n10,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n8,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n7,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n11,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n10,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n9,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n7,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n6,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n11,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n10,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n9,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n7,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n6,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n11,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n10,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n9,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n7,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n6,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n11,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n10,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n9,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n7,
         DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n6,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n12,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n11,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n10,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n8,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n7,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n12,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n11,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n10,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n8,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n7,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n12,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n11,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n10,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n8,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n7,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n12,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n11,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n10,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n8,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n7,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n12,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n11,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n10,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n8,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n7,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n11,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n10,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n8,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n7,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n11,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n10,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n8,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n7,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n11,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n10,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n8,
         DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n7,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n11,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n10,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n8,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n7,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n11,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n10,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n8,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n7,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n11,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n10,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n8,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n7,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n11,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n10,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n8,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n7,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n11,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n10,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n8,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n7,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n11,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n10,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n9,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n7,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n6,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n11,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n10,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n9,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n7,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n6,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n11,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n10,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n9,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n7,
         DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n6,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n11,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n10,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n8,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n7,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n11,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n10,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n8,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n7,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n10,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n9,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n7,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n6,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n11,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n10,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n8,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n7,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n11,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n10,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n8,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n7,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n11,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n10,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n8,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n7,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n11,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n10,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n8,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n7,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n10,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n9,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n7,
         DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n6,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n11,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n10,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n9,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n7,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n6,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n11,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n10,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n9,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n7,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n6,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n11,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n10,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n9,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n7,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n6,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n11,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n10,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n9,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n7,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n6,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n11,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n10,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n9,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n7,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n6,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n11,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n10,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n9,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n7,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n6,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n11,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n10,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n9,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n7,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n6,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n11,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n10,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n9,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n7,
         DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n6,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n11,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n10,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n8,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n7,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n11,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n10,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n8,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n7,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n11,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n10,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n8,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n7,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n11,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n10,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n8,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n7,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n11,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n10,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n8,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n7,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n11,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n10,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n8,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n7,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n11,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n10,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n8,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n7,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n11,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n10,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n8,
         DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n7,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n11,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n10,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n8,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n7,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n11,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n10,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n8,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n7,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n11,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n10,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n8,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n7,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n11,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n10,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n8,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n7,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n11,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n10,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n8,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n7,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n11,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n10,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n9,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n7,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n6,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n11,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n10,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n9,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n7,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n6,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n11,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n10,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n9,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n7,
         DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n6,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n11,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n10,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n8,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n7,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n11,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n10,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n9,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n7,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n6,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n11,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n10,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n9,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n7,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n6,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n11,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n10,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n9,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n7,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n6,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n11,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n10,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n9,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n7,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n6,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n11,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n10,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n9,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n7,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n6,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n11,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n10,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n9,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n7,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n6,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n11,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n10,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n9,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n7,
         DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n6,
         DataPath_Registers_Inst2_GEN_reg1_n230,
         DataPath_Registers_Inst2_GEN_reg1_n229,
         DataPath_Registers_Inst2_GEN_reg1_n228,
         DataPath_Registers_Inst2_GEN_reg1_n227,
         DataPath_Registers_Inst2_GEN_reg1_n226,
         DataPath_Registers_Inst2_GEN_reg1_n225,
         DataPath_Registers_Inst2_GEN_reg1_n224,
         DataPath_Registers_Inst2_GEN_reg1_n223,
         DataPath_Registers_Inst2_GEN_reg1_n222,
         DataPath_Registers_Inst2_GEN_reg1_n221,
         DataPath_Registers_Inst2_GEN_reg1_n220,
         DataPath_Registers_Inst2_GEN_reg1_n219,
         DataPath_Registers_Inst2_GEN_reg1_n218,
         DataPath_Registers_Inst2_GEN_reg1_n217,
         DataPath_Registers_Inst2_GEN_reg1_n216,
         DataPath_Registers_Inst2_GEN_reg1_n215,
         DataPath_Registers_Inst2_GEN_reg1_n214,
         DataPath_Registers_Inst2_GEN_reg1_n213,
         DataPath_Registers_Inst2_GEN_reg1_n212,
         DataPath_Registers_Inst2_GEN_reg1_n211,
         DataPath_Registers_Inst2_GEN_reg1_n210,
         DataPath_Registers_Inst2_GEN_reg1_n209,
         DataPath_Registers_Inst2_GEN_reg1_n208,
         DataPath_Registers_Inst2_GEN_reg1_n207,
         DataPath_Registers_Inst2_GEN_reg1_n206,
         DataPath_Registers_Inst2_GEN_reg1_n205,
         DataPath_Registers_Inst2_GEN_reg1_n204,
         DataPath_Registers_Inst2_GEN_reg1_n203,
         DataPath_Registers_Inst2_GEN_reg1_n202,
         DataPath_Registers_Inst2_GEN_reg1_n201,
         DataPath_Registers_Inst2_GEN_reg1_n200,
         DataPath_Registers_Inst2_GEN_reg1_n199,
         DataPath_Registers_Inst2_GEN_reg1_n198,
         DataPath_Registers_Inst2_GEN_reg1_n197,
         DataPath_Registers_Inst2_GEN_reg1_n196,
         DataPath_Registers_Inst2_GEN_reg1_n163,
         DataPath_Registers_Inst2_GEN_reg1_n162,
         DataPath_Registers_Inst2_GEN_reg1_n161,
         DataPath_Registers_Inst2_GEN_reg1_n160,
         DataPath_Registers_Inst2_GEN_reg1_n159,
         DataPath_Registers_Inst2_GEN_reg1_n158,
         DataPath_Registers_Inst2_GEN_reg1_n157,
         DataPath_Registers_Inst2_GEN_reg1_n156,
         DataPath_Registers_Inst2_GEN_reg1_n155,
         DataPath_Registers_Inst2_GEN_reg1_n154,
         DataPath_Registers_Inst2_GEN_reg1_n153,
         DataPath_Registers_Inst2_GEN_reg1_n152,
         DataPath_Registers_Inst2_GEN_reg1_n151,
         DataPath_Registers_Inst2_GEN_reg1_n150,
         DataPath_Registers_Inst2_GEN_reg1_n149,
         DataPath_Registers_Inst2_GEN_reg1_n148,
         DataPath_Registers_Inst2_GEN_reg1_n147,
         DataPath_Registers_Inst2_GEN_reg1_n146,
         DataPath_Registers_Inst2_GEN_reg1_n145,
         DataPath_Registers_Inst2_GEN_reg1_n144,
         DataPath_Registers_Inst2_GEN_reg1_n143,
         DataPath_Registers_Inst2_GEN_reg1_n142,
         DataPath_Registers_Inst2_GEN_reg1_n141,
         DataPath_Registers_Inst2_GEN_reg1_n140,
         DataPath_Registers_Inst2_GEN_reg1_n139,
         DataPath_Registers_Inst2_GEN_reg1_n138,
         DataPath_Registers_Inst2_GEN_reg1_n137,
         DataPath_Registers_Inst2_GEN_reg1_n136,
         DataPath_Registers_Inst2_GEN_reg1_n135,
         DataPath_Registers_Inst2_GEN_reg1_n134,
         DataPath_Registers_Inst2_GEN_reg1_n133,
         DataPath_Registers_Inst2_GEN_reg1_n132,
         DataPath_Registers_Inst2_GEN_reg1_n131,
         DataPath_Registers_Inst2_GEN_reg1_n130,
         DataPath_Registers_Inst2_GEN_reg1_n129,
         DataPath_Registers_Inst2_GEN_reg1_n128,
         DataPath_Registers_Inst2_GEN_reg1_n127,
         DataPath_Registers_Inst2_GEN_reg1_n126,
         DataPath_Registers_Inst2_GEN_reg1_n125,
         DataPath_Registers_Inst2_GEN_reg1_n124,
         DataPath_Registers_Inst2_GEN_reg1_n123,
         DataPath_Registers_Inst2_GEN_reg1_n122,
         DataPath_Registers_Inst2_GEN_reg1_n121,
         DataPath_Registers_Inst2_GEN_reg1_n120,
         DataPath_Registers_Inst2_GEN_reg1_n119,
         DataPath_Registers_Inst2_GEN_reg1_n118,
         DataPath_Registers_Inst2_GEN_reg1_n117,
         DataPath_Registers_Inst2_GEN_reg1_n116,
         DataPath_Registers_Inst2_GEN_reg1_n115,
         DataPath_Registers_Inst2_GEN_reg1_n114,
         DataPath_Registers_Inst2_GEN_reg1_n113,
         DataPath_Registers_Inst2_GEN_reg1_n112,
         DataPath_Registers_Inst2_GEN_reg1_n111,
         DataPath_Registers_Inst2_GEN_reg1_n110,
         DataPath_Registers_Inst2_GEN_reg1_n109,
         DataPath_Registers_Inst2_GEN_reg1_n108,
         DataPath_Registers_Inst2_GEN_reg1_n107,
         DataPath_Registers_Inst2_GEN_reg1_n106,
         DataPath_Registers_Inst2_GEN_reg1_n105,
         DataPath_Registers_Inst2_GEN_reg1_n104,
         DataPath_Registers_Inst2_GEN_reg1_n103,
         DataPath_Registers_Inst2_GEN_reg1_n102,
         DataPath_Registers_Inst2_GEN_reg1_n101,
         DataPath_Registers_Inst2_GEN_reg1_n100,
         DataPath_Registers_Inst2_A1_n12, DataPath_Registers_Inst2_A1_n11,
         DataPath_Registers_Inst2_A1_n10, DataPath_Registers_Inst2_A2_n12,
         DataPath_Registers_Inst2_A2_n11, DataPath_Registers_Inst2_A2_n10,
         DataPath_Registers_Inst2_A3_n12, DataPath_Registers_Inst2_A3_n11,
         DataPath_Registers_Inst2_A3_n10, DataPath_Registers_Inst2_A4_n12,
         DataPath_Registers_Inst2_A4_n11, DataPath_Registers_Inst2_A4_n10,
         Key_Registers_INST1_n317, Key_Registers_INST1_n316,
         Key_Registers_INST1_n315, Key_Registers_INST1_n314,
         Key_Registers_INST1_n313, Key_Registers_INST1_n312,
         Key_Registers_INST1_n311, Key_Registers_INST1_n310,
         Key_Registers_INST1_n309, Key_Registers_INST1_n308,
         Key_Registers_INST1_n307, Key_Registers_INST1_n306,
         Key_Registers_INST1_n305, Key_Registers_INST1_n304,
         Key_Registers_INST1_n303, Key_Registers_INST1_n302,
         Key_Registers_INST1_n301, Key_Registers_INST1_n300,
         Key_Registers_INST1_n299, Key_Registers_INST1_n298,
         Key_Registers_INST1_n297, Key_Registers_INST1_n296,
         Key_Registers_INST1_n295, Key_Registers_INST1_n294,
         Key_Registers_INST1_n293, Key_Registers_INST1_n292,
         Key_Registers_INST1_n291, Key_Registers_INST1_n290,
         Key_Registers_INST1_n289, Key_Registers_INST1_n288,
         Key_Registers_INST1_n287, Key_Registers_INST1_n286,
         Key_Registers_INST1_n285, Key_Registers_INST1_n284,
         Key_Registers_INST1_n283, Key_Registers_INST1_n282,
         Key_Registers_INST1_n281, Key_Registers_INST1_n280,
         Key_Registers_INST1_n279, Key_Registers_INST1_n278,
         Key_Registers_INST1_n277, Key_Registers_INST1_n276,
         Key_Registers_INST1_n275, Key_Registers_INST1_n274,
         Key_Registers_INST1_n273, Key_Registers_INST1_n272,
         Key_Registers_INST1_n271, Key_Registers_INST1_n270,
         Key_Registers_INST1_n269, Key_Registers_INST1_n268,
         Key_Registers_INST1_n267, Key_Registers_INST1_n266,
         Key_Registers_INST1_n265, Key_Registers_INST1_n264,
         Key_Registers_INST1_n263, Key_Registers_INST1_n262,
         Key_Registers_INST1_n261, Key_Registers_INST1_n260,
         Key_Registers_INST1_n259, Key_Registers_INST1_n258,
         Key_Registers_INST1_n257, Key_Registers_INST1_n256,
         Key_Registers_INST1_n255, Key_Registers_INST1_n254,
         Key_Registers_INST1_n253, Key_Registers_INST1_n252,
         Key_Registers_INST1_n251, Key_Registers_INST1_n250,
         Key_Registers_INST1_n249, Key_Registers_INST1_n248,
         Key_Registers_INST1_n247, Key_Registers_INST1_n246,
         Key_Registers_INST1_n245, Key_Registers_INST1_n244,
         Key_Registers_INST1_n243, Key_Registers_INST1_n242,
         Key_Registers_INST1_n241, Key_Registers_INST1_n240,
         Key_Registers_INST1_n239, Key_Registers_INST1_n238,
         Key_Registers_INST1_n237, Key_Registers_INST1_n236,
         Key_Registers_INST1_n235, Key_Registers_INST1_n234,
         Key_Registers_INST1_n233, Key_Registers_INST1_n232,
         Key_Registers_INST1_n231, Key_Registers_INST1_n230,
         Key_Registers_INST1_n229, Key_Registers_INST1_n228,
         Key_Registers_INST1_n227, Key_Registers_INST1_n129,
         Key_Registers_INST1_n127, Key_Registers_INST1_n124,
         Key_Registers_INST1_n121, Key_Registers_INST1_n118,
         Key_Registers_INST1_n115, Key_Registers_INST1_n112,
         Key_Registers_INST1_n109, Key_Registers_INST1_n106,
         Key_Registers_INST1_n105, Key_Registers_INST1_n103,
         Key_Registers_INST1_n102, Key_Registers_INST1_n100,
         Key_Registers_INST1_n99, Key_Registers_INST1_n97,
         Key_Registers_INST1_n96, Key_Registers_INST1_n94,
         Key_Registers_INST1_n93, Key_Registers_INST1_n91,
         Key_Registers_INST1_n90, Key_Registers_INST1_n88,
         Key_Registers_INST1_n87, Key_Registers_INST1_n85,
         Key_Registers_INST1_n84, Key_Registers_INST1_n82,
         Key_Registers_INST1_n81, Key_Registers_INST1_n79,
         Key_Registers_INST1_n78, Key_Registers_INST1_n76,
         Key_Registers_INST1_n75, Key_Registers_INST1_n73,
         Key_Registers_INST1_n72, Key_Registers_INST1_n226,
         Key_Registers_INST1_n225, Key_Registers_INST1_n224,
         Key_Registers_INST1_n223, Key_Registers_INST1_n222,
         Key_Registers_INST1_n221, Key_Registers_INST1_n220,
         Key_Registers_INST1_n219, Key_Registers_INST1_n218,
         Key_Registers_INST1_n217, Key_Registers_INST1_n216,
         Key_Registers_INST1_n215, Key_Registers_INST1_n214,
         Key_Registers_INST1_n213, Key_Registers_INST1_n212,
         Key_Registers_INST1_n211, Key_Registers_INST1_n210,
         Key_Registers_INST1_n209, Key_Registers_INST1_n208,
         Key_Registers_INST1_n207, Key_Registers_INST1_n206,
         Key_Registers_INST1_n205, Key_Registers_INST1_n204,
         Key_Registers_INST1_n203, Key_Registers_INST1_n202,
         Key_Registers_INST1_n201, Key_Registers_INST1_n200,
         Key_Registers_INST1_n199, Key_Registers_INST1_n198,
         Key_Registers_INST1_n197, Key_Registers_INST1_n196,
         Key_Registers_INST1_n195, Key_Registers_INST1_n194,
         Key_Registers_INST1_n193, Key_Registers_INST1_n192,
         Key_Registers_INST1_n191, Key_Registers_INST1_n190,
         Key_Registers_INST1_n189, Key_Registers_INST1_n188,
         Key_Registers_INST1_n187, Key_Registers_INST1_n186,
         Key_Registers_INST1_n185, Key_Registers_INST1_n184,
         Key_Registers_INST1_n183, Key_Registers_INST1_n182,
         Key_Registers_INST1_n181, Key_Registers_INST1_n180,
         Key_Registers_INST1_n179, Key_Registers_INST1_n178,
         Key_Registers_INST1_n177, Key_Registers_INST1_n176,
         Key_Registers_INST1_n175, Key_Registers_INST1_n174,
         Key_Registers_INST1_n173, Key_Registers_INST1_n172,
         Key_Registers_INST1_n171, Key_Registers_INST1_n170,
         Key_Registers_INST1_n169, Key_Registers_INST1_n168,
         Key_Registers_INST1_n167, Key_Registers_INST1_n166,
         Key_Registers_INST1_n165, Key_Registers_INST1_n164,
         Key_Registers_INST1_n163, Key_Registers_INST1_n162,
         Key_Registers_INST1_n161, Key_Registers_INST1_n160,
         Key_Registers_INST1_n159, Key_Registers_INST1_n158,
         Key_Registers_INST1_n157, Key_Registers_INST1_n156,
         Key_Registers_INST1_n155, Key_Registers_INST1_n154,
         Key_Registers_INST1_n152, Key_Registers_INST1_n151,
         Key_Registers_INST1_n149, Key_Registers_INST1_n148,
         Key_Registers_INST1_n146, Key_Registers_INST1_n145,
         Key_Registers_INST1_n143, Key_Registers_INST1_n142,
         Key_Registers_INST1_n140, Key_Registers_INST1_n139,
         Key_Registers_INST1_n137, Key_Registers_INST1_n136,
         Key_Registers_INST1_n134, Key_Registers_INST1_n133,
         Key_Registers_INST1_n131, Key_Registers_INST1_n130,
         Key_Registers_INST1_n128, Key_Registers_INST1_n126,
         Key_Registers_INST1_n125, Key_Registers_INST1_n123,
         Key_Registers_INST1_n122, Key_Registers_INST1_n120,
         Key_Registers_INST1_n119, Key_Registers_INST1_n117,
         Key_Registers_INST1_n116, Key_Registers_INST1_n114,
         Key_Registers_INST1_n113, Key_Registers_INST1_n111,
         Key_Registers_INST1_n110, Key_Registers_INST1_n108,
         Key_Registers_INST1_n107, Key_Registers_INST1_n104,
         Key_Registers_INST1_n101, Key_Registers_INST1_n98,
         Key_Registers_INST1_n95, Key_Registers_INST1_n92,
         Key_Registers_INST1_n89, Key_Registers_INST1_n86,
         Key_Registers_INST1_n83, Key_Registers_INST1_n80,
         Key_Registers_INST1_n77, Key_Registers_INST1_n74,
         Key_Registers_INST1_n71, Key_Registers_INST1_n68,
         Key_Registers_INST1_n65, Key_Registers_INST1_n62,
         Key_Registers_INST1_n59, Key_Registers_INST1_n56,
         Key_Registers_INST1_n53, Key_Registers_INST1_n50,
         Key_Registers_INST1_n47, Key_Registers_INST1_n44,
         Key_Registers_INST1_n41, Key_Registers_INST1_n38,
         Key_Registers_INST1_n35, Key_Registers_INST1_S8_0_,
         Key_Registers_INST1_S8_1_, Key_Registers_INST1_S8_2_,
         Key_Registers_INST1_S8_3_, Key_Registers_INST1_S8_4_,
         Key_Registers_INST1_S8_5_, Key_Registers_INST1_S8_6_,
         Key_Registers_INST1_S8_7_, Key_Registers_INST1_S4_0_,
         Key_Registers_INST1_S4_1_, Key_Registers_INST1_S4_2_,
         Key_Registers_INST1_S4_3_, Key_Registers_INST1_S4_4_,
         Key_Registers_INST1_S4_5_, Key_Registers_INST1_S4_6_,
         Key_Registers_INST1_S4_7_, Key_Registers_INST1_ScanFF_S3_SFF_0_n11,
         Key_Registers_INST1_ScanFF_S3_SFF_0_n10,
         Key_Registers_INST1_ScanFF_S3_SFF_0_n8,
         Key_Registers_INST1_ScanFF_S3_SFF_0_n7,
         Key_Registers_INST1_ScanFF_S3_SFF_1_n10,
         Key_Registers_INST1_ScanFF_S3_SFF_1_n9,
         Key_Registers_INST1_ScanFF_S3_SFF_1_n7,
         Key_Registers_INST1_ScanFF_S3_SFF_1_n6,
         Key_Registers_INST1_ScanFF_S3_SFF_2_n10,
         Key_Registers_INST1_ScanFF_S3_SFF_2_n9,
         Key_Registers_INST1_ScanFF_S3_SFF_2_n7,
         Key_Registers_INST1_ScanFF_S3_SFF_2_n6,
         Key_Registers_INST1_ScanFF_S3_SFF_3_n10,
         Key_Registers_INST1_ScanFF_S3_SFF_3_n9,
         Key_Registers_INST1_ScanFF_S3_SFF_3_n7,
         Key_Registers_INST1_ScanFF_S3_SFF_3_n6,
         Key_Registers_INST1_ScanFF_S3_SFF_4_n10,
         Key_Registers_INST1_ScanFF_S3_SFF_4_n9,
         Key_Registers_INST1_ScanFF_S3_SFF_4_n7,
         Key_Registers_INST1_ScanFF_S3_SFF_4_n6,
         Key_Registers_INST1_ScanFF_S3_SFF_5_n10,
         Key_Registers_INST1_ScanFF_S3_SFF_5_n9,
         Key_Registers_INST1_ScanFF_S3_SFF_5_n7,
         Key_Registers_INST1_ScanFF_S3_SFF_5_n6,
         Key_Registers_INST1_ScanFF_S3_SFF_6_n10,
         Key_Registers_INST1_ScanFF_S3_SFF_6_n9,
         Key_Registers_INST1_ScanFF_S3_SFF_6_n7,
         Key_Registers_INST1_ScanFF_S3_SFF_6_n6,
         Key_Registers_INST1_ScanFF_S3_SFF_7_n10,
         Key_Registers_INST1_ScanFF_S3_SFF_7_n9,
         Key_Registers_INST1_ScanFF_S3_SFF_7_n7,
         Key_Registers_INST1_ScanFF_S3_SFF_7_n6,
         Key_Registers_INST1_ScanFF_S7_SFF_0_n12,
         Key_Registers_INST1_ScanFF_S7_SFF_0_n11,
         Key_Registers_INST1_ScanFF_S7_SFF_0_n10,
         Key_Registers_INST1_ScanFF_S7_SFF_0_n8,
         Key_Registers_INST1_ScanFF_S7_SFF_0_n7,
         Key_Registers_INST1_ScanFF_S7_SFF_1_n13,
         Key_Registers_INST1_ScanFF_S7_SFF_1_n12,
         Key_Registers_INST1_ScanFF_S7_SFF_1_n11,
         Key_Registers_INST1_ScanFF_S7_SFF_1_n10,
         Key_Registers_INST1_ScanFF_S7_SFF_1_n8,
         Key_Registers_INST1_ScanFF_S7_SFF_1_n7,
         Key_Registers_INST1_ScanFF_S7_SFF_2_n13,
         Key_Registers_INST1_ScanFF_S7_SFF_2_n12,
         Key_Registers_INST1_ScanFF_S7_SFF_2_n11,
         Key_Registers_INST1_ScanFF_S7_SFF_2_n10,
         Key_Registers_INST1_ScanFF_S7_SFF_2_n8,
         Key_Registers_INST1_ScanFF_S7_SFF_2_n7,
         Key_Registers_INST1_ScanFF_S7_SFF_3_n13,
         Key_Registers_INST1_ScanFF_S7_SFF_3_n12,
         Key_Registers_INST1_ScanFF_S7_SFF_3_n11,
         Key_Registers_INST1_ScanFF_S7_SFF_3_n10,
         Key_Registers_INST1_ScanFF_S7_SFF_3_n8,
         Key_Registers_INST1_ScanFF_S7_SFF_3_n7,
         Key_Registers_INST1_ScanFF_S7_SFF_4_n13,
         Key_Registers_INST1_ScanFF_S7_SFF_4_n12,
         Key_Registers_INST1_ScanFF_S7_SFF_4_n11,
         Key_Registers_INST1_ScanFF_S7_SFF_4_n10,
         Key_Registers_INST1_ScanFF_S7_SFF_4_n8,
         Key_Registers_INST1_ScanFF_S7_SFF_4_n7,
         Key_Registers_INST1_ScanFF_S7_SFF_5_n13,
         Key_Registers_INST1_ScanFF_S7_SFF_5_n12,
         Key_Registers_INST1_ScanFF_S7_SFF_5_n11,
         Key_Registers_INST1_ScanFF_S7_SFF_5_n10,
         Key_Registers_INST1_ScanFF_S7_SFF_5_n8,
         Key_Registers_INST1_ScanFF_S7_SFF_5_n7,
         Key_Registers_INST1_ScanFF_S7_SFF_6_n13,
         Key_Registers_INST1_ScanFF_S7_SFF_6_n12,
         Key_Registers_INST1_ScanFF_S7_SFF_6_n11,
         Key_Registers_INST1_ScanFF_S7_SFF_6_n10,
         Key_Registers_INST1_ScanFF_S7_SFF_6_n8,
         Key_Registers_INST1_ScanFF_S7_SFF_6_n7,
         Key_Registers_INST1_ScanFF_S7_SFF_7_n13,
         Key_Registers_INST1_ScanFF_S7_SFF_7_n12,
         Key_Registers_INST1_ScanFF_S7_SFF_7_n11,
         Key_Registers_INST1_ScanFF_S7_SFF_7_n10,
         Key_Registers_INST1_ScanFF_S7_SFF_7_n8,
         Key_Registers_INST1_ScanFF_S7_SFF_7_n7,
         Key_Registers_INST1_ScanFF_S11_SFF_0_n14,
         Key_Registers_INST1_ScanFF_S11_SFF_0_n13,
         Key_Registers_INST1_ScanFF_S11_SFF_0_n12,
         Key_Registers_INST1_ScanFF_S11_SFF_0_n11,
         Key_Registers_INST1_ScanFF_S11_SFF_0_n10,
         Key_Registers_INST1_ScanFF_S11_SFF_0_n8,
         Key_Registers_INST1_ScanFF_S11_SFF_0_n7,
         Key_Registers_INST1_ScanFF_S11_SFF_1_n14,
         Key_Registers_INST1_ScanFF_S11_SFF_1_n13,
         Key_Registers_INST1_ScanFF_S11_SFF_1_n12,
         Key_Registers_INST1_ScanFF_S11_SFF_1_n11,
         Key_Registers_INST1_ScanFF_S11_SFF_1_n10,
         Key_Registers_INST1_ScanFF_S11_SFF_1_n8,
         Key_Registers_INST1_ScanFF_S11_SFF_1_n7,
         Key_Registers_INST1_ScanFF_S11_SFF_2_n14,
         Key_Registers_INST1_ScanFF_S11_SFF_2_n13,
         Key_Registers_INST1_ScanFF_S11_SFF_2_n12,
         Key_Registers_INST1_ScanFF_S11_SFF_2_n11,
         Key_Registers_INST1_ScanFF_S11_SFF_2_n10,
         Key_Registers_INST1_ScanFF_S11_SFF_2_n8,
         Key_Registers_INST1_ScanFF_S11_SFF_2_n7,
         Key_Registers_INST1_ScanFF_S11_SFF_3_n14,
         Key_Registers_INST1_ScanFF_S11_SFF_3_n13,
         Key_Registers_INST1_ScanFF_S11_SFF_3_n12,
         Key_Registers_INST1_ScanFF_S11_SFF_3_n11,
         Key_Registers_INST1_ScanFF_S11_SFF_3_n10,
         Key_Registers_INST1_ScanFF_S11_SFF_3_n8,
         Key_Registers_INST1_ScanFF_S11_SFF_3_n7,
         Key_Registers_INST1_ScanFF_S11_SFF_4_n14,
         Key_Registers_INST1_ScanFF_S11_SFF_4_n13,
         Key_Registers_INST1_ScanFF_S11_SFF_4_n12,
         Key_Registers_INST1_ScanFF_S11_SFF_4_n11,
         Key_Registers_INST1_ScanFF_S11_SFF_4_n10,
         Key_Registers_INST1_ScanFF_S11_SFF_4_n8,
         Key_Registers_INST1_ScanFF_S11_SFF_4_n7,
         Key_Registers_INST1_ScanFF_S11_SFF_5_n11,
         Key_Registers_INST1_ScanFF_S11_SFF_5_n10,
         Key_Registers_INST1_ScanFF_S11_SFF_5_n9,
         Key_Registers_INST1_ScanFF_S11_SFF_5_n7,
         Key_Registers_INST1_ScanFF_S11_SFF_5_n6,
         Key_Registers_INST1_ScanFF_S11_SFF_6_n13,
         Key_Registers_INST1_ScanFF_S11_SFF_6_n12,
         Key_Registers_INST1_ScanFF_S11_SFF_6_n11,
         Key_Registers_INST1_ScanFF_S11_SFF_6_n10,
         Key_Registers_INST1_ScanFF_S11_SFF_6_n9,
         Key_Registers_INST1_ScanFF_S11_SFF_6_n7,
         Key_Registers_INST1_ScanFF_S11_SFF_6_n6,
         Key_Registers_INST1_ScanFF_S11_SFF_7_n13,
         Key_Registers_INST1_ScanFF_S11_SFF_7_n12,
         Key_Registers_INST1_ScanFF_S11_SFF_7_n11,
         Key_Registers_INST1_ScanFF_S11_SFF_7_n10,
         Key_Registers_INST1_ScanFF_S11_SFF_7_n9,
         Key_Registers_INST1_ScanFF_S11_SFF_7_n7,
         Key_Registers_INST1_ScanFF_S11_SFF_7_n6,
         Key_Registers_INST1_ScanFF_S15_SFF_0_n12,
         Key_Registers_INST1_ScanFF_S15_SFF_0_n11,
         Key_Registers_INST1_ScanFF_S15_SFF_0_n10,
         Key_Registers_INST1_ScanFF_S15_SFF_0_n8,
         Key_Registers_INST1_ScanFF_S15_SFF_0_n7,
         Key_Registers_INST1_ScanFF_S15_SFF_1_n13,
         Key_Registers_INST1_ScanFF_S15_SFF_1_n12,
         Key_Registers_INST1_ScanFF_S15_SFF_1_n11,
         Key_Registers_INST1_ScanFF_S15_SFF_1_n10,
         Key_Registers_INST1_ScanFF_S15_SFF_1_n9,
         Key_Registers_INST1_ScanFF_S15_SFF_1_n7,
         Key_Registers_INST1_ScanFF_S15_SFF_1_n6,
         Key_Registers_INST1_ScanFF_S15_SFF_2_n13,
         Key_Registers_INST1_ScanFF_S15_SFF_2_n12,
         Key_Registers_INST1_ScanFF_S15_SFF_2_n11,
         Key_Registers_INST1_ScanFF_S15_SFF_2_n10,
         Key_Registers_INST1_ScanFF_S15_SFF_2_n9,
         Key_Registers_INST1_ScanFF_S15_SFF_2_n7,
         Key_Registers_INST1_ScanFF_S15_SFF_2_n6,
         Key_Registers_INST1_ScanFF_S15_SFF_3_n13,
         Key_Registers_INST1_ScanFF_S15_SFF_3_n12,
         Key_Registers_INST1_ScanFF_S15_SFF_3_n11,
         Key_Registers_INST1_ScanFF_S15_SFF_3_n10,
         Key_Registers_INST1_ScanFF_S15_SFF_3_n9,
         Key_Registers_INST1_ScanFF_S15_SFF_3_n7,
         Key_Registers_INST1_ScanFF_S15_SFF_3_n6,
         Key_Registers_INST1_ScanFF_S15_SFF_4_n13,
         Key_Registers_INST1_ScanFF_S15_SFF_4_n12,
         Key_Registers_INST1_ScanFF_S15_SFF_4_n11,
         Key_Registers_INST1_ScanFF_S15_SFF_4_n10,
         Key_Registers_INST1_ScanFF_S15_SFF_4_n9,
         Key_Registers_INST1_ScanFF_S15_SFF_4_n7,
         Key_Registers_INST1_ScanFF_S15_SFF_4_n6,
         Key_Registers_INST1_ScanFF_S15_SFF_5_n13,
         Key_Registers_INST1_ScanFF_S15_SFF_5_n12,
         Key_Registers_INST1_ScanFF_S15_SFF_5_n11,
         Key_Registers_INST1_ScanFF_S15_SFF_5_n10,
         Key_Registers_INST1_ScanFF_S15_SFF_5_n9,
         Key_Registers_INST1_ScanFF_S15_SFF_5_n7,
         Key_Registers_INST1_ScanFF_S15_SFF_5_n6,
         Key_Registers_INST1_ScanFF_S15_SFF_6_n13,
         Key_Registers_INST1_ScanFF_S15_SFF_6_n12,
         Key_Registers_INST1_ScanFF_S15_SFF_6_n11,
         Key_Registers_INST1_ScanFF_S15_SFF_6_n10,
         Key_Registers_INST1_ScanFF_S15_SFF_6_n9,
         Key_Registers_INST1_ScanFF_S15_SFF_6_n7,
         Key_Registers_INST1_ScanFF_S15_SFF_6_n6,
         Key_Registers_INST1_ScanFF_S15_SFF_7_n13,
         Key_Registers_INST1_ScanFF_S15_SFF_7_n12,
         Key_Registers_INST1_ScanFF_S15_SFF_7_n11,
         Key_Registers_INST1_ScanFF_S15_SFF_7_n10,
         Key_Registers_INST1_ScanFF_S15_SFF_7_n9,
         Key_Registers_INST1_ScanFF_S15_SFF_7_n7,
         Key_Registers_INST1_ScanFF_S15_SFF_7_n6,
         GF256Inv_o_InputAffine_Inst1_A1_n9,
         GF256Inv_o_InputAffine_Inst1_A1_n8,
         GF256Inv_o_InputAffine_Inst1_A1_n7,
         GF256Inv_o_InputAffine_Inst1_A1_n6,
         GF256Inv_o_InputAffine_Inst1_A1_n5,
         GF256Inv_o_InputAffine_Inst1_A1_n4,
         GF256Inv_o_InputAffine_Inst1_A1_n3,
         GF256Inv_o_InputAffine_Inst1_A2_n28,
         GF256Inv_o_InputAffine_Inst1_A2_n27,
         GF256Inv_o_InputAffine_Inst1_A2_n26,
         GF256Inv_o_InputAffine_Inst1_A2_n25,
         GF256Inv_o_InputAffine_Inst1_A2_n24,
         GF256Inv_o_InputAffine_Inst1_A2_n23,
         GF256Inv_o_InputAffine_Inst1_A2_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n81,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n80,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n79,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n78,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n77,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n76,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n75,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n74,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n73,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n72,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n71,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n70,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n69,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n68,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n67,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n66,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n65,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n64,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n63,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n62,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n61,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n60,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n59,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n58,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n57,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n56,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n55,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n54,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n53,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n52,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n51,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n50,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n49,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n48,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n47,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n46,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n45,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n44,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n43,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n42,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n41,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n40,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n39,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n38,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n59,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n58,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n57,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n56,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n55,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n54,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n53,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n52,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n51,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n50,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n49,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n48,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n47,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n46,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n45,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n44,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n43,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n42,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n41,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n40,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n39,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n38,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n37,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n36,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n35,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n34,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n33,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n32,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n31,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n30,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n29,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n28,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n27,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n26,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n25,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n24,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n23,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n21,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n20,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n19,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n18,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n17,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n16,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n15,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n11,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n10,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n9,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n8,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n61,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n60,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n59,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n58,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n57,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n56,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n55,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n54,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n53,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n52,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n51,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n50,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n49,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n48,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n47,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n46,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n45,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n44,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n43,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n42,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n41,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n40,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n39,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n38,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n37,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n36,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n35,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n34,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n33,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n32,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n31,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n30,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n29,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n28,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n27,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n26,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n17,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n16,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n15,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n14,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n13,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n12,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n11,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n10,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n98,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n97,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n96,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n95,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n94,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n93,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n92,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n91,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n90,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n89,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n88,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n87,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n86,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n85,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n84,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n83,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n82,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n81,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n80,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n79,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n78,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n77,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n76,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n75,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n74,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n73,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n72,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n71,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n70,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n69,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n68,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n67,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n66,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n65,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n61,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n59,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n56,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n54,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n53,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n52,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n51,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n50,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n49,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n48,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n47,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n7,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n61,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n59,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n56,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_n8,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n39,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n38,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n37,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n36,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n35,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n33,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n25,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n24,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n23,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n21,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n20,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n28,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n27,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n26,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n25,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n24,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n23,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n20,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n19,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n18,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n17,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n16,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n17,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n16,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n15,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n14,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n13,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n24,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n23,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n21,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n20,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n19,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n18,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n17,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n7,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n61,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n59,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n56,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_n8,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n39,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n38,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n37,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n36,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n35,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n33,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n25,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n24,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n23,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n21,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n20,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n28,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n27,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n26,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n25,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n24,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n23,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n20,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n19,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n18,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n17,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n16,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n17,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n16,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n15,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n14,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n13,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n24,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n23,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n22,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n21,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n20,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n19,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n18,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n17,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n6,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n5,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n133,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n132,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n131,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n130,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n129,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n128,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n100,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n110,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n109,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n108,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n107,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n106,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n105,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n104,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n103,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n102,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n101,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n98,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n133,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n132,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n131,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n130,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n129,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n128,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n100,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n110,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n109,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n108,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n107,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n106,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n105,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n104,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n103,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n102,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n101,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99,
         GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n98,
         Inst_Controller_n178, Inst_Controller_n177, Inst_Controller_n176,
         Inst_Controller_n175, Inst_Controller_n174, Inst_Controller_n173,
         Inst_Controller_n172, Inst_Controller_n171, Inst_Controller_n170,
         Inst_Controller_n169, Inst_Controller_n168, Inst_Controller_n167,
         Inst_Controller_n166, Inst_Controller_n165, Inst_Controller_n164,
         Inst_Controller_n163, Inst_Controller_n162, Inst_Controller_n161,
         Inst_Controller_n160, Inst_Controller_n159, Inst_Controller_n158,
         Inst_Controller_n157, Inst_Controller_n156, Inst_Controller_n155,
         Inst_Controller_n154, Inst_Controller_n153, Inst_Controller_n152,
         Inst_Controller_n151, Inst_Controller_n150, Inst_Controller_n149,
         Inst_Controller_n148, Inst_Controller_n147, Inst_Controller_n146,
         Inst_Controller_n145, Inst_Controller_n144, Inst_Controller_n143,
         Inst_Controller_n142, Inst_Controller_n141, Inst_Controller_n140,
         Inst_Controller_n139, Inst_Controller_n138, Inst_Controller_n137,
         Inst_Controller_n136, Inst_Controller_n135, Inst_Controller_n134,
         Inst_Controller_n133, Inst_Controller_n132, Inst_Controller_n131,
         Inst_Controller_n130, Inst_Controller_n129, Inst_Controller_n128,
         Inst_Controller_n127, Inst_Controller_n126, Inst_Controller_n125,
         Inst_Controller_n124, Inst_Controller_n123, Inst_Controller_n122,
         Inst_Controller_n121, Inst_Controller_n120, Inst_Controller_n119,
         Inst_Controller_n118, Inst_Controller_n117, Inst_Controller_n116,
         Inst_Controller_n115, Inst_Controller_n100, Inst_Controller_n99,
         Inst_Controller_n98, Inst_Controller_n97, Inst_Controller_n94,
         Inst_Controller_n91, Inst_Controller_n90, Inst_Controller_n6,
         Inst_Controller_n114, Inst_Controller_n113, Inst_Controller_n112,
         Inst_Controller_n111, Inst_Controller_n110, Inst_Controller_n109,
         Inst_Controller_n108, Inst_Controller_n107, Inst_Controller_n106,
         Inst_Controller_n105, Inst_Controller_n104, Inst_Controller_n103,
         Inst_Controller_n44, Inst_Controller_n39, Inst_Controller_n37,
         Inst_Controller_n35, Inst_Controller_n33, Inst_Controller_n26,
         Inst_Controller_n25, Inst_Controller_n24, Inst_Controller_n23,
         Inst_Controller_n22, Inst_Controller_n21, Inst_Controller_n20,
         Inst_Controller_n19, Inst_Controller_N86, Inst_Controller_N84,
         Inst_Controller_N83, Inst_Controller_N82, Inst_Controller_N81,
         Inst_Controller_PerRoundCounter_0_, Inst_Controller_n179;
  wire   [7:0] KeyOut1;
  wire   [7:0] KeyForSchedule1;
  wire   [7:0] S0_output1;
  wire   [7:0] KeySchedule_out1;
  wire   [7:0] MCout_xor_SKey_2;
  wire   [7:0] K_ciphertext1;
  wire   [7:0] Affined_Inv_K0_xor_K12_1;
  wire   [7:0] OutputReg_in1;
  wire   [7:0] OutputReg1;
  wire   [7:0] OutputReg2;
  wire   [7:0] Rcon_1;
  wire   [7:0] Rcon_internal;
  wire   [7:0] StateIn1;
  wire   [7:0] StateIn2;
  wire   [1:0] SboxIn_sel;
  wire   [7:1] SboxIn1;
  wire   [7:0] KeyToSbox1;
  wire   [1:0] KeyIn_sel;
  wire   [7:0] KeyIn1;
  wire   [7:0] KeySchedule_Inst1_Reg_in;
  wire   [7:0] KeySchedule_Inst1_S_key2_reg;
  wire   [7:0] KeySchedule_Inst1_Reg_out;
  wire   [7:0] KeySchedule_Inst1_Key_out_tmp;
  wire   [7:0] KeySchedule_Inst1_Affined_Inv_K0;
  wire   [7:0] DataPath_Registers_Inst1_reg_A_output4_1;
  wire   [7:0] DataPath_Registers_Inst1_reg_A_output3_1;
  wire   [7:0] DataPath_Registers_Inst1_reg_A_output2_1;
  wire   [7:0] DataPath_Registers_Inst1_reg_A_output1_1;
  wire   [7:0] DataPath_Registers_Inst1_out4;
  wire   [7:0] DataPath_Registers_Inst1_out3;
  wire   [7:0] DataPath_Registers_Inst1_out2;
  wire   [7:0] DataPath_Registers_Inst1_out1;
  wire   [7:0] DataPath_Registers_Inst1_S12_in;
  wire   [7:0] DataPath_Registers_Inst1_S8_in;
  wire   [7:0] DataPath_Registers_Inst1_S4_in;
  wire   [7:0] DataPath_Registers_Inst2_reg_A_output4_1;
  wire   [7:0] DataPath_Registers_Inst2_reg_A_output3_1;
  wire   [7:0] DataPath_Registers_Inst2_reg_A_output2_1;
  wire   [7:0] DataPath_Registers_Inst2_reg_A_output1_1;
  wire   [7:0] DataPath_Registers_Inst2_out4;
  wire   [7:0] DataPath_Registers_Inst2_out3;
  wire   [7:0] DataPath_Registers_Inst2_out2;
  wire   [7:0] DataPath_Registers_Inst2_out1;
  wire   [7:0] DataPath_Registers_Inst2_S12_in;
  wire   [7:0] DataPath_Registers_Inst2_S8_in;
  wire   [7:0] DataPath_Registers_Inst2_S4_in;
  wire   [7:0] Key_Registers_INST1_S14_in;
  wire   [7:0] Key_Registers_INST1_S10_in;
  wire   [7:0] Key_Registers_INST1_S6_in;
  wire   [7:0] Key_Registers_INST1_S2_in;
  wire   [7:0] GF256Inv_o_InputAffine_Inst1_inv_input2_reg;
  wire   [7:0] GF256Inv_o_InputAffine_Inst1_inv_input1_reg;
  wire   [7:0] GF256Inv_o_InputAffine_Inst1_inv_input2;
  wire   [7:0] GF256Inv_o_InputAffine_Inst1_inv_input1;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg
;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg
;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg
;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg
;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg3;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg3;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg3;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg3;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg2;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg2;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg
;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg2;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg2;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg1;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg1;
  wire   [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2;
  wire   [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1;
  wire   [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2;
  wire   [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg1;
  wire   [3:0] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg1;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu_reg
;
  wire  
         [3:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd
;
  wire  
         [3:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd
;
  wire  
         [4:2] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y
;
  wire  
         [8:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x_reg
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y
;
  wire  
         [4:1] GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x
;

  DFF_X1 Done_reg ( .D(done_internal), .CK(clk), .Q(Done), .QN() );
  INV_X1 U288 ( .A(n331), .ZN(n164) );
  INV_X1 U289 ( .A(n316), .ZN(n314) );
  INV_X1 U290 ( .A(n317), .ZN(n315) );
  NOR2_X2 U291 ( .A1(SboxIn_sel[0]), .A2(SboxIn_sel[1]), .ZN(n332) );
  INV_X1 U293 ( .A(key[0]), .ZN(n274) );
  OR2_X1 U294 ( .A1(KeyIn_sel[1]), .A2(KeyIn_sel[0]), .ZN(n261) );
  INV_X1 U295 ( .A(KeyIn_sel[0]), .ZN(n251) );
  NOR2_X1 U296 ( .A1(KeyIn_sel[1]), .A2(n251), .ZN(n259) );
  XOR2_X1 U297 ( .A(KeyForSchedule1[0]), .B(KeyOut1[0]), .Z(n171) );
  AOI22_X1 U298 ( .A1(KeySchedule_out1[0]), .A2(n259), .B1(n171), .B2(
        KeyIn_sel[1]), .ZN(n252) );
  OAI21_X1 U299 ( .B1(n274), .B2(n261), .A(n252), .ZN(KeyIn1[0]) );
  INV_X1 U300 ( .A(key[1]), .ZN(n280) );
  XOR2_X1 U301 ( .A(KeyForSchedule1[1]), .B(KeyOut1[1]), .Z(n172) );
  AOI22_X1 U302 ( .A1(KeySchedule_out1[1]), .A2(n259), .B1(n172), .B2(
        KeyIn_sel[1]), .ZN(n253) );
  OAI21_X1 U303 ( .B1(n280), .B2(n261), .A(n253), .ZN(KeyIn1[1]) );
  INV_X1 U304 ( .A(key[2]), .ZN(n286) );
  XOR2_X1 U305 ( .A(KeyForSchedule1[2]), .B(KeyOut1[2]), .Z(n173) );
  AOI22_X1 U306 ( .A1(KeySchedule_out1[2]), .A2(n259), .B1(n173), .B2(
        KeyIn_sel[1]), .ZN(n254) );
  OAI21_X1 U307 ( .B1(n286), .B2(n261), .A(n254), .ZN(KeyIn1[2]) );
  INV_X1 U308 ( .A(key[3]), .ZN(n292) );
  XOR2_X1 U309 ( .A(KeyForSchedule1[3]), .B(KeyOut1[3]), .Z(n174) );
  AOI22_X1 U310 ( .A1(KeySchedule_out1[3]), .A2(n259), .B1(n174), .B2(
        KeyIn_sel[1]), .ZN(n255) );
  OAI21_X1 U311 ( .B1(n292), .B2(n261), .A(n255), .ZN(KeyIn1[3]) );
  INV_X1 U312 ( .A(key[4]), .ZN(n298) );
  XOR2_X1 U313 ( .A(KeyForSchedule1[4]), .B(KeyOut1[4]), .Z(n175) );
  AOI22_X1 U314 ( .A1(KeySchedule_out1[4]), .A2(n259), .B1(n175), .B2(
        KeyIn_sel[1]), .ZN(n256) );
  OAI21_X1 U315 ( .B1(n298), .B2(n261), .A(n256), .ZN(KeyIn1[4]) );
  INV_X1 U316 ( .A(key[5]), .ZN(n304) );
  XOR2_X1 U317 ( .A(KeyForSchedule1[5]), .B(KeyOut1[5]), .Z(n176) );
  AOI22_X1 U318 ( .A1(KeySchedule_out1[5]), .A2(n259), .B1(n176), .B2(
        KeyIn_sel[1]), .ZN(n257) );
  OAI21_X1 U319 ( .B1(n304), .B2(n261), .A(n257), .ZN(KeyIn1[5]) );
  INV_X1 U320 ( .A(key[6]), .ZN(n310) );
  XOR2_X1 U321 ( .A(KeyForSchedule1[6]), .B(KeyOut1[6]), .Z(n177) );
  AOI22_X1 U322 ( .A1(KeySchedule_out1[6]), .A2(n259), .B1(n177), .B2(
        KeyIn_sel[1]), .ZN(n258) );
  OAI21_X1 U323 ( .B1(n310), .B2(n261), .A(n258), .ZN(KeyIn1[6]) );
  INV_X1 U324 ( .A(key[7]), .ZN(n321) );
  XOR2_X1 U325 ( .A(KeyForSchedule1[7]), .B(KeyOut1[7]), .Z(n178) );
  AOI22_X1 U326 ( .A1(KeySchedule_out1[7]), .A2(n259), .B1(n178), .B2(
        KeyIn_sel[1]), .ZN(n260) );
  OAI21_X1 U327 ( .B1(n321), .B2(n261), .A(n260), .ZN(KeyIn1[7]) );
  INV_X1 U328 ( .A(Output_Sel), .ZN(n269) );
  AOI22_X1 U329 ( .A1(Output_Sel), .A2(Affined_Inv_K0_xor_K12_1[0]), .B1(
        K_ciphertext1[0]), .B2(n269), .ZN(n262) );
  XNOR2_X1 U330 ( .A(S0_output1[0]), .B(n262), .ZN(OutputReg_in1[0]) );
  AOI22_X1 U331 ( .A1(Output_Sel), .A2(Affined_Inv_K0_xor_K12_1[1]), .B1(
        K_ciphertext1[1]), .B2(n269), .ZN(n263) );
  XNOR2_X1 U332 ( .A(S0_output1[1]), .B(n263), .ZN(OutputReg_in1[1]) );
  AOI22_X1 U333 ( .A1(Output_Sel), .A2(Affined_Inv_K0_xor_K12_1[2]), .B1(
        K_ciphertext1[2]), .B2(n269), .ZN(n264) );
  XNOR2_X1 U334 ( .A(S0_output1[2]), .B(n264), .ZN(OutputReg_in1[2]) );
  AOI22_X1 U335 ( .A1(Output_Sel), .A2(Affined_Inv_K0_xor_K12_1[3]), .B1(
        K_ciphertext1[3]), .B2(n269), .ZN(n265) );
  XNOR2_X1 U336 ( .A(S0_output1[3]), .B(n265), .ZN(OutputReg_in1[3]) );
  AOI22_X1 U337 ( .A1(Output_Sel), .A2(Affined_Inv_K0_xor_K12_1[4]), .B1(
        K_ciphertext1[4]), .B2(n269), .ZN(n266) );
  XNOR2_X1 U338 ( .A(S0_output1[4]), .B(n266), .ZN(OutputReg_in1[4]) );
  AOI22_X1 U339 ( .A1(Output_Sel), .A2(Affined_Inv_K0_xor_K12_1[5]), .B1(
        K_ciphertext1[5]), .B2(n269), .ZN(n267) );
  XNOR2_X1 U340 ( .A(S0_output1[5]), .B(n267), .ZN(OutputReg_in1[5]) );
  AOI22_X1 U341 ( .A1(Output_Sel), .A2(Affined_Inv_K0_xor_K12_1[6]), .B1(
        K_ciphertext1[6]), .B2(n269), .ZN(n268) );
  XNOR2_X1 U342 ( .A(S0_output1[6]), .B(n268), .ZN(OutputReg_in1[6]) );
  AOI22_X1 U343 ( .A1(Output_Sel), .A2(Affined_Inv_K0_xor_K12_1[7]), .B1(
        K_ciphertext1[7]), .B2(n269), .ZN(n270) );
  XNOR2_X1 U344 ( .A(S0_output1[7]), .B(n270), .ZN(OutputReg_in1[7]) );
  AND2_X1 U345 ( .A1(ShowRcon), .A2(Rcon_internal[0]), .ZN(Rcon_1[0]) );
  AND2_X1 U346 ( .A1(ShowRcon), .A2(Rcon_internal[1]), .ZN(Rcon_1[1]) );
  AND2_X1 U347 ( .A1(ShowRcon), .A2(Rcon_internal[2]), .ZN(Rcon_1[2]) );
  AND2_X1 U348 ( .A1(ShowRcon), .A2(Rcon_internal[3]), .ZN(Rcon_1[3]) );
  AND2_X1 U349 ( .A1(ShowRcon), .A2(Rcon_internal[4]), .ZN(Rcon_1[4]) );
  AND2_X1 U350 ( .A1(ShowRcon), .A2(Rcon_internal[5]), .ZN(Rcon_1[5]) );
  AND2_X1 U351 ( .A1(ShowRcon), .A2(Rcon_internal[6]), .ZN(Rcon_1[6]) );
  AND2_X1 U352 ( .A1(ShowRcon), .A2(Rcon_internal[7]), .ZN(Rcon_1[7]) );
  INV_X1 U353 ( .A(SboxIn_sel[0]), .ZN(n271) );
  NAND2_X1 U354 ( .A1(n271), .A2(SboxIn_sel[1]), .ZN(n317) );
  NAND2_X1 U355 ( .A1(SboxIn_sel[0]), .A2(SboxIn_sel[1]), .ZN(n316) );
  AOI22_X1 U356 ( .A1(n315), .A2(KeySchedule_out1[0]), .B1(n314), .B2(n171), 
        .ZN(n277) );
  NOR2_X1 U357 ( .A1(SboxIn_sel[1]), .A2(n271), .ZN(n319) );
  OAI22_X1 U358 ( .A1(KeySchedule_out1[0]), .A2(n317), .B1(n171), .B2(n316), 
        .ZN(n272) );
  AOI22_X1 U359 ( .A1(KeyToSbox1[0]), .A2(n319), .B1(S0_output1[0]), .B2(n272), 
        .ZN(n276) );
  INV_X1 U360 ( .A(input1[0]), .ZN(n273) );
  OAI221_X1 U361 ( .B1(key[0]), .B2(input1[0]), .C1(n274), .C2(n273), .A(n332), 
        .ZN(n275) );
  OAI211_X1 U362 ( .C1(S0_output1[0]), .C2(n277), .A(n276), .B(n275), .ZN(
        GF256Inv_o_InputAffine_Inst1_inv_input1[2]) );
  AOI22_X1 U363 ( .A1(n315), .A2(KeySchedule_out1[1]), .B1(n314), .B2(n172), 
        .ZN(n283) );
  OAI22_X1 U364 ( .A1(KeySchedule_out1[1]), .A2(n317), .B1(n172), .B2(n316), 
        .ZN(n278) );
  AOI22_X1 U365 ( .A1(n319), .A2(KeyToSbox1[1]), .B1(S0_output1[1]), .B2(n278), 
        .ZN(n282) );
  INV_X1 U366 ( .A(input1[1]), .ZN(n279) );
  OAI221_X1 U367 ( .B1(key[1]), .B2(input1[1]), .C1(n280), .C2(n279), .A(n332), 
        .ZN(n281) );
  OAI211_X1 U368 ( .C1(S0_output1[1]), .C2(n283), .A(n282), .B(n281), .ZN(
        SboxIn1[1]) );
  AOI22_X1 U369 ( .A1(n315), .A2(KeySchedule_out1[2]), .B1(n314), .B2(n173), 
        .ZN(n289) );
  OAI22_X1 U370 ( .A1(KeySchedule_out1[2]), .A2(n317), .B1(n173), .B2(n316), 
        .ZN(n284) );
  AOI22_X1 U371 ( .A1(n319), .A2(KeyToSbox1[2]), .B1(S0_output1[2]), .B2(n284), 
        .ZN(n288) );
  INV_X1 U372 ( .A(input1[2]), .ZN(n285) );
  OAI221_X1 U373 ( .B1(key[2]), .B2(input1[2]), .C1(n286), .C2(n285), .A(n332), 
        .ZN(n287) );
  OAI211_X1 U374 ( .C1(S0_output1[2]), .C2(n289), .A(n288), .B(n287), .ZN(
        SboxIn1[2]) );
  AOI22_X1 U375 ( .A1(n315), .A2(KeySchedule_out1[3]), .B1(n314), .B2(n174), 
        .ZN(n295) );
  OAI22_X1 U376 ( .A1(KeySchedule_out1[3]), .A2(n317), .B1(n174), .B2(n316), 
        .ZN(n290) );
  AOI22_X1 U377 ( .A1(n319), .A2(KeyToSbox1[3]), .B1(S0_output1[3]), .B2(n290), 
        .ZN(n294) );
  INV_X1 U378 ( .A(input1[3]), .ZN(n291) );
  OAI221_X1 U379 ( .B1(key[3]), .B2(input1[3]), .C1(n292), .C2(n291), .A(n332), 
        .ZN(n293) );
  OAI211_X1 U380 ( .C1(S0_output1[3]), .C2(n295), .A(n294), .B(n293), .ZN(
        SboxIn1[3]) );
  AOI22_X1 U381 ( .A1(n315), .A2(KeySchedule_out1[4]), .B1(n314), .B2(n175), 
        .ZN(n301) );
  OAI22_X1 U382 ( .A1(KeySchedule_out1[4]), .A2(n317), .B1(n175), .B2(n316), 
        .ZN(n296) );
  AOI22_X1 U383 ( .A1(n319), .A2(KeyToSbox1[4]), .B1(S0_output1[4]), .B2(n296), 
        .ZN(n300) );
  INV_X1 U384 ( .A(input1[4]), .ZN(n297) );
  OAI221_X1 U385 ( .B1(key[4]), .B2(input1[4]), .C1(n298), .C2(n297), .A(n332), 
        .ZN(n299) );
  OAI211_X1 U386 ( .C1(S0_output1[4]), .C2(n301), .A(n300), .B(n299), .ZN(
        SboxIn1[4]) );
  AOI22_X1 U387 ( .A1(n315), .A2(KeySchedule_out1[5]), .B1(n314), .B2(n176), 
        .ZN(n307) );
  OAI22_X1 U388 ( .A1(KeySchedule_out1[5]), .A2(n317), .B1(n176), .B2(n316), 
        .ZN(n302) );
  AOI22_X1 U389 ( .A1(n319), .A2(KeyToSbox1[5]), .B1(S0_output1[5]), .B2(n302), 
        .ZN(n306) );
  INV_X1 U390 ( .A(input1[5]), .ZN(n303) );
  OAI221_X1 U391 ( .B1(key[5]), .B2(input1[5]), .C1(n304), .C2(n303), .A(n332), 
        .ZN(n305) );
  OAI211_X1 U392 ( .C1(S0_output1[5]), .C2(n307), .A(n306), .B(n305), .ZN(
        SboxIn1[5]) );
  AOI22_X1 U393 ( .A1(n315), .A2(KeySchedule_out1[6]), .B1(n314), .B2(n177), 
        .ZN(n313) );
  OAI22_X1 U394 ( .A1(KeySchedule_out1[6]), .A2(n317), .B1(n177), .B2(n316), 
        .ZN(n308) );
  AOI22_X1 U395 ( .A1(n319), .A2(KeyToSbox1[6]), .B1(S0_output1[6]), .B2(n308), 
        .ZN(n312) );
  INV_X1 U396 ( .A(input1[6]), .ZN(n309) );
  OAI221_X1 U397 ( .B1(key[6]), .B2(input1[6]), .C1(n310), .C2(n309), .A(n332), 
        .ZN(n311) );
  OAI211_X1 U398 ( .C1(S0_output1[6]), .C2(n313), .A(n312), .B(n311), .ZN(
        SboxIn1[6]) );
  AOI22_X1 U399 ( .A1(n315), .A2(KeySchedule_out1[7]), .B1(n314), .B2(n178), 
        .ZN(n324) );
  OAI22_X1 U400 ( .A1(KeySchedule_out1[7]), .A2(n317), .B1(n178), .B2(n316), 
        .ZN(n318) );
  AOI22_X1 U401 ( .A1(n319), .A2(KeyToSbox1[7]), .B1(S0_output1[7]), .B2(n318), 
        .ZN(n323) );
  INV_X1 U402 ( .A(input1[7]), .ZN(n320) );
  OAI221_X1 U403 ( .B1(key[7]), .B2(input1[7]), .C1(n321), .C2(n320), .A(n332), 
        .ZN(n322) );
  OAI211_X1 U404 ( .C1(S0_output1[7]), .C2(n324), .A(n323), .B(n322), .ZN(
        SboxIn1[7]) );
  XOR2_X1 U405 ( .A(Corr_63_5_), .B(output1_A_1_), .Z(output1[1]) );
  XOR2_X1 U406 ( .A(Corr_63_5_), .B(output1_A_2_), .Z(output1[2]) );
  XOR2_X1 U407 ( .A(Corr_63_5_), .B(output1_A_4_), .Z(output1[4]) );
  XOR2_X1 U408 ( .A(Corr_63_5_), .B(output1_A_5_), .Z(output1[5]) );
  AOI22_X1 U409 ( .A1(SboxIn_sel[1]), .A2(MCout_xor_SKey_2[7]), .B1(n332), 
        .B2(input2[7]), .ZN(n325) );
  INV_X1 U410 ( .A(n325), .ZN(n170) );
  AOI22_X1 U411 ( .A1(SboxIn_sel[1]), .A2(MCout_xor_SKey_2[6]), .B1(n332), 
        .B2(input2[6]), .ZN(n326) );
  INV_X1 U412 ( .A(n326), .ZN(n169) );
  AOI22_X1 U413 ( .A1(SboxIn_sel[1]), .A2(MCout_xor_SKey_2[5]), .B1(n332), 
        .B2(input2[5]), .ZN(n327) );
  INV_X1 U414 ( .A(n327), .ZN(n168) );
  AOI22_X1 U415 ( .A1(SboxIn_sel[1]), .A2(MCout_xor_SKey_2[4]), .B1(n332), 
        .B2(input2[4]), .ZN(n328) );
  INV_X1 U416 ( .A(n328), .ZN(n167) );
  AOI22_X1 U417 ( .A1(SboxIn_sel[1]), .A2(MCout_xor_SKey_2[3]), .B1(n332), 
        .B2(input2[3]), .ZN(n329) );
  INV_X1 U418 ( .A(n329), .ZN(n166) );
  AOI22_X1 U419 ( .A1(SboxIn_sel[1]), .A2(MCout_xor_SKey_2[2]), .B1(n332), 
        .B2(input2[2]), .ZN(n330) );
  INV_X1 U420 ( .A(n330), .ZN(n165) );
  AOI22_X1 U421 ( .A1(SboxIn_sel[1]), .A2(MCout_xor_SKey_2[1]), .B1(n332), 
        .B2(input2[1]), .ZN(n331) );
  AOI22_X1 U422 ( .A1(SboxIn_sel[1]), .A2(MCout_xor_SKey_2[0]), .B1(n332), 
        .B2(input2[0]), .ZN(n333) );
  INV_X1 U423 ( .A(n333), .ZN(GF256Inv_o_InputAffine_Inst1_inv_input2[2]) );
  XOR2_X1 Affine_OutInv1_U12 ( .A(n175), .B(n178), .Z(
        Affined_Inv_K0_xor_K12_1[7]) );
  XNOR2_X1 Affine_OutInv1_U11 ( .A(Affine_OutInv1_n4), .B(Affine_OutInv1_n3), 
        .ZN(Affined_Inv_K0_xor_K12_1[4]) );
  XNOR2_X1 Affine_OutInv1_U10 ( .A(n177), .B(n174), .ZN(Affine_OutInv1_n4) );
  XOR2_X1 Affine_OutInv1_U9 ( .A(n178), .B(Affined_Inv_K0_xor_K12_1[5]), .Z(
        Affined_Inv_K0_xor_K12_1[3]) );
  XNOR2_X1 Affine_OutInv1_U8 ( .A(n173), .B(Affine_OutInv1_n2), .ZN(
        Affined_Inv_K0_xor_K12_1[2]) );
  XOR2_X1 Affine_OutInv1_U7 ( .A(n176), .B(n178), .Z(Affine_OutInv1_n2) );
  XNOR2_X1 Affine_OutInv1_U6 ( .A(n174), .B(Affine_OutInv1_n1), .ZN(
        Affined_Inv_K0_xor_K12_1[1]) );
  XOR2_X1 Affine_OutInv1_U5 ( .A(n171), .B(n175), .Z(Affine_OutInv1_n1) );
  XNOR2_X1 Affine_OutInv1_U4 ( .A(n176), .B(Affined_Inv_K0_xor_K12_1[6]), .ZN(
        Affined_Inv_K0_xor_K12_1[0]) );
  XNOR2_X1 Affine_OutInv1_U3 ( .A(Affine_OutInv1_n3), .B(
        Affined_Inv_K0_xor_K12_1[5]), .ZN(Affined_Inv_K0_xor_K12_1[6]) );
  XNOR2_X1 Affine_OutInv1_U2 ( .A(n171), .B(n172), .ZN(Affine_OutInv1_n3) );
  XNOR2_X1 Affine_OutInv1_U1 ( .A(n175), .B(n177), .ZN(
        Affined_Inv_K0_xor_K12_1[5]) );
  OAI21_X1 OutputReg_U37 ( .B1(OutputReg_n67), .B2(OutputReg_n27), .A(
        OutputReg_n66), .ZN(OutputReg_n36) );
  NAND2_X1 OutputReg_U36 ( .A1(OutputReg_n65), .A2(MCout_xor_SKey_2[7]), .ZN(
        OutputReg_n66) );
  OAI21_X1 OutputReg_U35 ( .B1(OutputReg_n67), .B2(OutputReg_n26), .A(
        OutputReg_n64), .ZN(OutputReg_n37) );
  NAND2_X1 OutputReg_U34 ( .A1(OutputReg_n65), .A2(MCout_xor_SKey_2[6]), .ZN(
        OutputReg_n64) );
  OAI21_X1 OutputReg_U33 ( .B1(OutputReg_n67), .B2(OutputReg_n25), .A(
        OutputReg_n63), .ZN(OutputReg_n38) );
  NAND2_X1 OutputReg_U32 ( .A1(OutputReg_n65), .A2(MCout_xor_SKey_2[5]), .ZN(
        OutputReg_n63) );
  OAI21_X1 OutputReg_U31 ( .B1(OutputReg_n67), .B2(OutputReg_n24), .A(
        OutputReg_n62), .ZN(OutputReg_n39) );
  NAND2_X1 OutputReg_U30 ( .A1(OutputReg_n65), .A2(MCout_xor_SKey_2[4]), .ZN(
        OutputReg_n62) );
  OAI21_X1 OutputReg_U29 ( .B1(OutputReg_n67), .B2(OutputReg_n23), .A(
        OutputReg_n61), .ZN(OutputReg_n40) );
  NAND2_X1 OutputReg_U28 ( .A1(OutputReg_n65), .A2(MCout_xor_SKey_2[3]), .ZN(
        OutputReg_n61) );
  OAI21_X1 OutputReg_U27 ( .B1(OutputReg_n67), .B2(OutputReg_n22), .A(
        OutputReg_n60), .ZN(OutputReg_n41) );
  NAND2_X1 OutputReg_U26 ( .A1(OutputReg_n65), .A2(MCout_xor_SKey_2[2]), .ZN(
        OutputReg_n60) );
  OAI21_X1 OutputReg_U25 ( .B1(OutputReg_n67), .B2(OutputReg_n21), .A(
        OutputReg_n59), .ZN(OutputReg_n42) );
  NAND2_X1 OutputReg_U24 ( .A1(OutputReg_n65), .A2(MCout_xor_SKey_2[1]), .ZN(
        OutputReg_n59) );
  OAI21_X1 OutputReg_U23 ( .B1(OutputReg_n67), .B2(OutputReg_n20), .A(
        OutputReg_n58), .ZN(OutputReg_n43) );
  NAND2_X1 OutputReg_U22 ( .A1(OutputReg_n65), .A2(MCout_xor_SKey_2[0]), .ZN(
        OutputReg_n58) );
  OAI21_X1 OutputReg_U21 ( .B1(OutputReg_n67), .B2(OutputReg_n35), .A(
        OutputReg_n57), .ZN(OutputReg_n44) );
  NAND2_X1 OutputReg_U20 ( .A1(OutputReg_n65), .A2(OutputReg_in1[7]), .ZN(
        OutputReg_n57) );
  OAI21_X1 OutputReg_U19 ( .B1(OutputReg_n67), .B2(OutputReg_n34), .A(
        OutputReg_n56), .ZN(OutputReg_n45) );
  NAND2_X1 OutputReg_U18 ( .A1(OutputReg_n65), .A2(OutputReg_in1[6]), .ZN(
        OutputReg_n56) );
  OAI21_X1 OutputReg_U17 ( .B1(OutputReg_n67), .B2(OutputReg_n33), .A(
        OutputReg_n55), .ZN(OutputReg_n46) );
  NAND2_X1 OutputReg_U16 ( .A1(OutputReg_n65), .A2(OutputReg_in1[5]), .ZN(
        OutputReg_n55) );
  OAI21_X1 OutputReg_U15 ( .B1(OutputReg_n67), .B2(OutputReg_n32), .A(
        OutputReg_n54), .ZN(OutputReg_n47) );
  NAND2_X1 OutputReg_U14 ( .A1(OutputReg_n65), .A2(OutputReg_in1[4]), .ZN(
        OutputReg_n54) );
  OAI21_X1 OutputReg_U13 ( .B1(OutputReg_n67), .B2(OutputReg_n31), .A(
        OutputReg_n53), .ZN(OutputReg_n48) );
  NAND2_X1 OutputReg_U12 ( .A1(OutputReg_n65), .A2(OutputReg_in1[3]), .ZN(
        OutputReg_n53) );
  OAI21_X1 OutputReg_U11 ( .B1(OutputReg_n67), .B2(OutputReg_n30), .A(
        OutputReg_n52), .ZN(OutputReg_n49) );
  NAND2_X1 OutputReg_U10 ( .A1(OutputReg_n65), .A2(OutputReg_in1[2]), .ZN(
        OutputReg_n52) );
  OAI21_X1 OutputReg_U9 ( .B1(OutputReg_n67), .B2(OutputReg_n29), .A(
        OutputReg_n19), .ZN(OutputReg_n50) );
  NAND2_X1 OutputReg_U8 ( .A1(OutputReg_n65), .A2(OutputReg_in1[1]), .ZN(
        OutputReg_n19) );
  OAI21_X1 OutputReg_U7 ( .B1(OutputReg_n67), .B2(OutputReg_n28), .A(
        OutputReg_n18), .ZN(OutputReg_n51) );
  NAND2_X1 OutputReg_U6 ( .A1(OutputReg_n65), .A2(OutputReg_in1[0]), .ZN(
        OutputReg_n18) );
  NOR2_X1 OutputReg_U5 ( .A1(rst), .A2(done_internal), .ZN(OutputReg_n17) );
  NOR2_X2 OutputReg_U4 ( .A1(rst), .A2(OutputReg_n17), .ZN(OutputReg_n65) );
  INV_X1 OutputReg_U3 ( .A(OutputReg_n17), .ZN(OutputReg_n67) );
  DFF_X1 OutputReg_Q_reg_0_ ( .D(OutputReg_n51), .CK(clk), .Q(OutputReg1[0]), 
        .QN(OutputReg_n28) );
  DFF_X1 OutputReg_Q_reg_1_ ( .D(OutputReg_n50), .CK(clk), .Q(OutputReg1[1]), 
        .QN(OutputReg_n29) );
  DFF_X1 OutputReg_Q_reg_2_ ( .D(OutputReg_n49), .CK(clk), .Q(OutputReg1[2]), 
        .QN(OutputReg_n30) );
  DFF_X1 OutputReg_Q_reg_3_ ( .D(OutputReg_n48), .CK(clk), .Q(OutputReg1[3]), 
        .QN(OutputReg_n31) );
  DFF_X1 OutputReg_Q_reg_4_ ( .D(OutputReg_n47), .CK(clk), .Q(OutputReg1[4]), 
        .QN(OutputReg_n32) );
  DFF_X1 OutputReg_Q_reg_5_ ( .D(OutputReg_n46), .CK(clk), .Q(OutputReg1[5]), 
        .QN(OutputReg_n33) );
  DFF_X1 OutputReg_Q_reg_6_ ( .D(OutputReg_n45), .CK(clk), .Q(OutputReg1[6]), 
        .QN(OutputReg_n34) );
  DFF_X1 OutputReg_Q_reg_7_ ( .D(OutputReg_n44), .CK(clk), .Q(OutputReg1[7]), 
        .QN(OutputReg_n35) );
  DFF_X1 OutputReg_Q_reg_8_ ( .D(OutputReg_n43), .CK(clk), .Q(OutputReg2[0]), 
        .QN(OutputReg_n20) );
  DFF_X1 OutputReg_Q_reg_9_ ( .D(OutputReg_n42), .CK(clk), .Q(OutputReg2[1]), 
        .QN(OutputReg_n21) );
  DFF_X1 OutputReg_Q_reg_10_ ( .D(OutputReg_n41), .CK(clk), .Q(OutputReg2[2]), 
        .QN(OutputReg_n22) );
  DFF_X1 OutputReg_Q_reg_11_ ( .D(OutputReg_n40), .CK(clk), .Q(OutputReg2[3]), 
        .QN(OutputReg_n23) );
  DFF_X1 OutputReg_Q_reg_12_ ( .D(OutputReg_n39), .CK(clk), .Q(OutputReg2[4]), 
        .QN(OutputReg_n24) );
  DFF_X1 OutputReg_Q_reg_13_ ( .D(OutputReg_n38), .CK(clk), .Q(OutputReg2[5]), 
        .QN(OutputReg_n25) );
  DFF_X1 OutputReg_Q_reg_14_ ( .D(OutputReg_n37), .CK(clk), .Q(OutputReg2[6]), 
        .QN(OutputReg_n26) );
  DFF_X1 OutputReg_Q_reg_15_ ( .D(OutputReg_n36), .CK(clk), .Q(OutputReg2[7]), 
        .QN(OutputReg_n27) );
  XNOR2_X1 Affine_output_Inst_U11 ( .A(output1_A_4_), .B(
        Affine_output_Inst_n12), .ZN(output1[3]) );
  XNOR2_X1 Affine_output_Inst_U10 ( .A(Affine_output_Inst_n11), .B(
        output1_A_5_), .ZN(output1_A_2_) );
  XNOR2_X1 Affine_output_Inst_U9 ( .A(output1[7]), .B(OutputReg1[2]), .ZN(
        Affine_output_Inst_n11) );
  XOR2_X1 Affine_output_Inst_U8 ( .A(OutputReg1[6]), .B(OutputReg1[0]), .Z(
        output1_A_5_) );
  XNOR2_X1 Affine_output_Inst_U7 ( .A(Affine_output_Inst_n10), .B(
        OutputReg1[1]), .ZN(output1_A_1_) );
  XNOR2_X1 Affine_output_Inst_U6 ( .A(OutputReg1[5]), .B(OutputReg1[4]), .ZN(
        Affine_output_Inst_n10) );
  XNOR2_X1 Affine_output_Inst_U5 ( .A(OutputReg1[1]), .B(
        Affine_output_Inst_n12), .ZN(output1[0]) );
  XNOR2_X1 Affine_output_Inst_U4 ( .A(OutputReg1[6]), .B(OutputReg1[4]), .ZN(
        Affine_output_Inst_n12) );
  XOR2_X1 Affine_output_Inst_U3 ( .A(OutputReg1[5]), .B(output1[6]), .Z(
        output1_A_4_) );
  XOR2_X1 Affine_output_Inst_U2 ( .A(OutputReg1[3]), .B(OutputReg1[7]), .Z(
        output1[6]) );
  XOR2_X1 Affine_output_Inst_U1 ( .A(OutputReg1[5]), .B(OutputReg1[3]), .Z(
        output1[7]) );
  XNOR2_X1 Affine_outputC_Inst_U11 ( .A(output2[4]), .B(
        Affine_outputC_Inst_n12), .ZN(output2[3]) );
  XNOR2_X1 Affine_outputC_Inst_U10 ( .A(Affine_outputC_Inst_n11), .B(
        output2[5]), .ZN(output2[2]) );
  XNOR2_X1 Affine_outputC_Inst_U9 ( .A(output2[7]), .B(OutputReg2[2]), .ZN(
        Affine_outputC_Inst_n11) );
  XOR2_X1 Affine_outputC_Inst_U8 ( .A(OutputReg2[6]), .B(OutputReg2[0]), .Z(
        output2[5]) );
  XNOR2_X1 Affine_outputC_Inst_U7 ( .A(Affine_outputC_Inst_n10), .B(
        OutputReg2[1]), .ZN(output2[1]) );
  XNOR2_X1 Affine_outputC_Inst_U6 ( .A(OutputReg2[5]), .B(OutputReg2[4]), .ZN(
        Affine_outputC_Inst_n10) );
  XNOR2_X1 Affine_outputC_Inst_U5 ( .A(OutputReg2[1]), .B(
        Affine_outputC_Inst_n12), .ZN(output2[0]) );
  XNOR2_X1 Affine_outputC_Inst_U4 ( .A(OutputReg2[6]), .B(OutputReg2[4]), .ZN(
        Affine_outputC_Inst_n12) );
  XOR2_X1 Affine_outputC_Inst_U3 ( .A(OutputReg2[5]), .B(output2[6]), .Z(
        output2[4]) );
  XOR2_X1 Affine_outputC_Inst_U2 ( .A(OutputReg2[3]), .B(OutputReg2[7]), .Z(
        output2[6]) );
  XOR2_X1 Affine_outputC_Inst_U1 ( .A(OutputReg2[5]), .B(OutputReg2[3]), .Z(
        output2[7]) );
  XOR2_X1 KeySchedule_Inst1_U24 ( .A(KeySchedule_Inst1_Affined_Inv_K0[7]), .B(
        StateIn1[7]), .Z(KeySchedule_Inst1_Reg_in[7]) );
  XOR2_X1 KeySchedule_Inst1_U23 ( .A(KeySchedule_Inst1_Affined_Inv_K0[6]), .B(
        StateIn1[6]), .Z(KeySchedule_Inst1_Reg_in[6]) );
  XOR2_X1 KeySchedule_Inst1_U22 ( .A(KeySchedule_Inst1_Affined_Inv_K0[5]), .B(
        StateIn1[5]), .Z(KeySchedule_Inst1_Reg_in[5]) );
  XOR2_X1 KeySchedule_Inst1_U21 ( .A(KeySchedule_Inst1_Affined_Inv_K0[4]), .B(
        StateIn1[4]), .Z(KeySchedule_Inst1_Reg_in[4]) );
  XOR2_X1 KeySchedule_Inst1_U20 ( .A(KeySchedule_Inst1_Affined_Inv_K0[3]), .B(
        StateIn1[3]), .Z(KeySchedule_Inst1_Reg_in[3]) );
  XOR2_X1 KeySchedule_Inst1_U19 ( .A(KeySchedule_Inst1_Affined_Inv_K0[2]), .B(
        StateIn1[2]), .Z(KeySchedule_Inst1_Reg_in[2]) );
  XOR2_X1 KeySchedule_Inst1_U18 ( .A(KeySchedule_Inst1_Affined_Inv_K0[1]), .B(
        StateIn1[1]), .Z(KeySchedule_Inst1_Reg_in[1]) );
  XOR2_X1 KeySchedule_Inst1_U17 ( .A(KeySchedule_Inst1_Affined_Inv_K0[0]), .B(
        StateIn1[0]), .Z(KeySchedule_Inst1_Reg_in[0]) );
  XOR2_X1 KeySchedule_Inst1_U16 ( .A(KeySchedule_Inst1_Key_out_tmp[7]), .B(
        Rcon_1[7]), .Z(KeySchedule_out1[7]) );
  XOR2_X1 KeySchedule_Inst1_U15 ( .A(KeySchedule_Inst1_Key_out_tmp[6]), .B(
        Rcon_1[6]), .Z(KeySchedule_out1[6]) );
  XOR2_X1 KeySchedule_Inst1_U14 ( .A(KeySchedule_Inst1_Key_out_tmp[5]), .B(
        Rcon_1[5]), .Z(KeySchedule_out1[5]) );
  XOR2_X1 KeySchedule_Inst1_U13 ( .A(KeySchedule_Inst1_Key_out_tmp[4]), .B(
        Rcon_1[4]), .Z(KeySchedule_out1[4]) );
  XOR2_X1 KeySchedule_Inst1_U12 ( .A(KeySchedule_Inst1_Key_out_tmp[3]), .B(
        Rcon_1[3]), .Z(KeySchedule_out1[3]) );
  XOR2_X1 KeySchedule_Inst1_U11 ( .A(KeySchedule_Inst1_Key_out_tmp[2]), .B(
        Rcon_1[2]), .Z(KeySchedule_out1[2]) );
  XOR2_X1 KeySchedule_Inst1_U10 ( .A(KeySchedule_Inst1_Key_out_tmp[1]), .B(
        Rcon_1[1]), .Z(KeySchedule_out1[1]) );
  XOR2_X1 KeySchedule_Inst1_U9 ( .A(KeySchedule_Inst1_Key_out_tmp[0]), .B(
        Rcon_1[0]), .Z(KeySchedule_out1[0]) );
  XOR2_X1 KeySchedule_Inst1_U8 ( .A(KeySchedule_Inst1_Reg_out[7]), .B(
        KeySchedule_Inst1_S_key2_reg[7]), .Z(K_ciphertext1[7]) );
  XOR2_X1 KeySchedule_Inst1_U7 ( .A(KeySchedule_Inst1_Reg_out[6]), .B(
        KeySchedule_Inst1_S_key2_reg[6]), .Z(K_ciphertext1[6]) );
  XOR2_X1 KeySchedule_Inst1_U6 ( .A(KeySchedule_Inst1_Reg_out[5]), .B(
        KeySchedule_Inst1_S_key2_reg[5]), .Z(K_ciphertext1[5]) );
  XOR2_X1 KeySchedule_Inst1_U5 ( .A(KeySchedule_Inst1_Reg_out[4]), .B(
        KeySchedule_Inst1_S_key2_reg[4]), .Z(K_ciphertext1[4]) );
  XOR2_X1 KeySchedule_Inst1_U4 ( .A(KeySchedule_Inst1_Reg_out[3]), .B(
        KeySchedule_Inst1_S_key2_reg[3]), .Z(K_ciphertext1[3]) );
  XOR2_X1 KeySchedule_Inst1_U3 ( .A(KeySchedule_Inst1_Reg_out[2]), .B(
        KeySchedule_Inst1_S_key2_reg[2]), .Z(K_ciphertext1[2]) );
  XOR2_X1 KeySchedule_Inst1_U2 ( .A(KeySchedule_Inst1_Reg_out[1]), .B(
        KeySchedule_Inst1_S_key2_reg[1]), .Z(K_ciphertext1[1]) );
  XOR2_X1 KeySchedule_Inst1_U1 ( .A(KeySchedule_Inst1_Reg_out[0]), .B(
        KeySchedule_Inst1_S_key2_reg[0]), .Z(K_ciphertext1[0]) );
  XOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U12 ( .A(KeyOut1[4]), .B(KeyOut1[7]), .Z(KeySchedule_Inst1_Affined_Inv_K0[7]) );
  XNOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U11 ( .A(
        KeySchedule_Inst1_Affine_OutInv1_n4), .B(
        KeySchedule_Inst1_Affine_OutInv1_n3), .ZN(
        KeySchedule_Inst1_Affined_Inv_K0[4]) );
  XOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U10 ( .A(KeyOut1[6]), .B(KeyOut1[3]), .Z(KeySchedule_Inst1_Affine_OutInv1_n3) );
  XOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U9 ( .A(
        KeySchedule_Inst1_Affined_Inv_K0[5]), .B(KeyOut1[7]), .Z(
        KeySchedule_Inst1_Affined_Inv_K0[3]) );
  XNOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U8 ( .A(
        KeySchedule_Inst1_Affine_OutInv1_n2), .B(KeyOut1[2]), .ZN(
        KeySchedule_Inst1_Affined_Inv_K0[2]) );
  XNOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U7 ( .A(KeyOut1[5]), .B(KeyOut1[7]), .ZN(KeySchedule_Inst1_Affine_OutInv1_n2) );
  XNOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U6 ( .A(
        KeySchedule_Inst1_Affine_OutInv1_n1), .B(KeyOut1[3]), .ZN(
        KeySchedule_Inst1_Affined_Inv_K0[1]) );
  XNOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U5 ( .A(KeyOut1[0]), .B(KeyOut1[4]), .ZN(KeySchedule_Inst1_Affine_OutInv1_n1) );
  XOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U4 ( .A(KeyOut1[5]), .B(
        KeySchedule_Inst1_Affined_Inv_K0[6]), .Z(
        KeySchedule_Inst1_Affined_Inv_K0[0]) );
  XNOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U3 ( .A(
        KeySchedule_Inst1_Affined_Inv_K0[5]), .B(
        KeySchedule_Inst1_Affine_OutInv1_n4), .ZN(
        KeySchedule_Inst1_Affined_Inv_K0[6]) );
  XNOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U2 ( .A(KeyOut1[0]), .B(KeyOut1[1]), .ZN(KeySchedule_Inst1_Affine_OutInv1_n4) );
  XOR2_X1 KeySchedule_Inst1_Affine_OutInv1_U1 ( .A(KeyOut1[4]), .B(KeyOut1[6]), 
        .Z(KeySchedule_Inst1_Affined_Inv_K0[5]) );
  XNOR2_X1 KeySchedule_Inst1_A1_U11 ( .A(KeySchedule_Inst1_Key_out_tmp[4]), 
        .B(KeySchedule_Inst1_A1_n14), .ZN(KeySchedule_Inst1_Key_out_tmp[3]) );
  XNOR2_X1 KeySchedule_Inst1_A1_U10 ( .A(KeySchedule_Inst1_Key_out_tmp[5]), 
        .B(KeySchedule_Inst1_A1_n13), .ZN(KeySchedule_Inst1_Key_out_tmp[2]) );
  XOR2_X1 KeySchedule_Inst1_A1_U9 ( .A(KeySchedule_Inst1_Key_out_tmp[7]), .B(
        K_ciphertext1[2]), .Z(KeySchedule_Inst1_A1_n13) );
  XNOR2_X1 KeySchedule_Inst1_A1_U8 ( .A(K_ciphertext1[6]), .B(K_ciphertext1[0]), .ZN(KeySchedule_Inst1_Key_out_tmp[5]) );
  XOR2_X1 KeySchedule_Inst1_A1_U7 ( .A(K_ciphertext1[1]), .B(
        KeySchedule_Inst1_A1_n14), .Z(KeySchedule_Inst1_Key_out_tmp[0]) );
  XNOR2_X1 KeySchedule_Inst1_A1_U6 ( .A(K_ciphertext1[6]), .B(K_ciphertext1[4]), .ZN(KeySchedule_Inst1_A1_n14) );
  XNOR2_X1 KeySchedule_Inst1_A1_U5 ( .A(K_ciphertext1[1]), .B(
        KeySchedule_Inst1_A1_n12), .ZN(KeySchedule_Inst1_Key_out_tmp[1]) );
  XOR2_X1 KeySchedule_Inst1_A1_U4 ( .A(K_ciphertext1[5]), .B(K_ciphertext1[4]), 
        .Z(KeySchedule_Inst1_A1_n12) );
  XNOR2_X1 KeySchedule_Inst1_A1_U3 ( .A(K_ciphertext1[5]), .B(
        KeySchedule_Inst1_Key_out_tmp[6]), .ZN(
        KeySchedule_Inst1_Key_out_tmp[4]) );
  XNOR2_X1 KeySchedule_Inst1_A1_U2 ( .A(K_ciphertext1[3]), .B(K_ciphertext1[7]), .ZN(KeySchedule_Inst1_Key_out_tmp[6]) );
  XOR2_X1 KeySchedule_Inst1_A1_U1 ( .A(K_ciphertext1[5]), .B(K_ciphertext1[3]), 
        .Z(KeySchedule_Inst1_Key_out_tmp[7]) );
  OAI21_X1 KeySchedule_Inst1_GEN_reg_U18 ( .B1(KeySchedule_Inst1_GEN_reg_n26), 
        .B2(KeySchedule_Inst1_GEN_reg_n16), .A(KeySchedule_Inst1_GEN_reg_n34), 
        .ZN(KeySchedule_Inst1_GEN_reg_n24) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg_U17 ( .A1(KeySchedule_Inst1_GEN_reg_n26), 
        .A2(KeySchedule_Inst1_Reg_in[7]), .ZN(KeySchedule_Inst1_GEN_reg_n34)
         );
  OAI21_X1 KeySchedule_Inst1_GEN_reg_U16 ( .B1(KeySchedule_Inst1_GEN_reg_n26), 
        .B2(KeySchedule_Inst1_GEN_reg_n15), .A(KeySchedule_Inst1_GEN_reg_n33), 
        .ZN(KeySchedule_Inst1_GEN_reg_n23) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg_U15 ( .A1(KeySchedule_Inst1_GEN_reg_n26), 
        .A2(KeySchedule_Inst1_Reg_in[6]), .ZN(KeySchedule_Inst1_GEN_reg_n33)
         );
  OAI21_X1 KeySchedule_Inst1_GEN_reg_U14 ( .B1(KeySchedule_Inst1_GEN_reg_n26), 
        .B2(KeySchedule_Inst1_GEN_reg_n14), .A(KeySchedule_Inst1_GEN_reg_n32), 
        .ZN(KeySchedule_Inst1_GEN_reg_n22) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg_U13 ( .A1(KeySchedule_Inst1_GEN_reg_n26), 
        .A2(KeySchedule_Inst1_Reg_in[5]), .ZN(KeySchedule_Inst1_GEN_reg_n32)
         );
  OAI21_X1 KeySchedule_Inst1_GEN_reg_U12 ( .B1(KeySchedule_Inst1_GEN_reg_n26), 
        .B2(KeySchedule_Inst1_GEN_reg_n13), .A(KeySchedule_Inst1_GEN_reg_n31), 
        .ZN(KeySchedule_Inst1_GEN_reg_n21) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg_U11 ( .A1(KeySchedule_Inst1_GEN_reg_n26), 
        .A2(KeySchedule_Inst1_Reg_in[4]), .ZN(KeySchedule_Inst1_GEN_reg_n31)
         );
  OAI21_X1 KeySchedule_Inst1_GEN_reg_U10 ( .B1(KeySchedule_Inst1_GEN_reg_n26), 
        .B2(KeySchedule_Inst1_GEN_reg_n12), .A(KeySchedule_Inst1_GEN_reg_n30), 
        .ZN(KeySchedule_Inst1_GEN_reg_n20) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg_U9 ( .A1(KeySchedule_Inst1_GEN_reg_n26), 
        .A2(KeySchedule_Inst1_Reg_in[3]), .ZN(KeySchedule_Inst1_GEN_reg_n30)
         );
  OAI21_X1 KeySchedule_Inst1_GEN_reg_U8 ( .B1(KeySchedule_Inst1_GEN_reg_n26), 
        .B2(KeySchedule_Inst1_GEN_reg_n11), .A(KeySchedule_Inst1_GEN_reg_n29), 
        .ZN(KeySchedule_Inst1_GEN_reg_n19) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg_U7 ( .A1(KeySchedule_Inst1_GEN_reg_n26), 
        .A2(KeySchedule_Inst1_Reg_in[2]), .ZN(KeySchedule_Inst1_GEN_reg_n29)
         );
  OAI21_X1 KeySchedule_Inst1_GEN_reg_U6 ( .B1(KeySchedule_Inst1_GEN_reg_n26), 
        .B2(KeySchedule_Inst1_GEN_reg_n10), .A(KeySchedule_Inst1_GEN_reg_n28), 
        .ZN(KeySchedule_Inst1_GEN_reg_n18) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg_U5 ( .A1(KeySchedule_Inst1_GEN_reg_n26), 
        .A2(KeySchedule_Inst1_Reg_in[1]), .ZN(KeySchedule_Inst1_GEN_reg_n28)
         );
  OAI21_X1 KeySchedule_Inst1_GEN_reg_U4 ( .B1(KeySchedule_Inst1_GEN_reg_n26), 
        .B2(KeySchedule_Inst1_GEN_reg_n9), .A(KeySchedule_Inst1_GEN_reg_n27), 
        .ZN(KeySchedule_Inst1_GEN_reg_n17) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg_U3 ( .A1(KeySchedule_Inst1_GEN_reg_n26), 
        .A2(KeySchedule_Inst1_Reg_in[0]), .ZN(KeySchedule_Inst1_GEN_reg_n27)
         );
  BUF_X1 KeySchedule_Inst1_GEN_reg_U2 ( .A(KeyScheduleRegisterEN), .Z(
        KeySchedule_Inst1_GEN_reg_n26) );
  DFF_X1 KeySchedule_Inst1_GEN_reg_Q_reg_0_ ( .D(KeySchedule_Inst1_GEN_reg_n17), .CK(clk), .Q(KeySchedule_Inst1_Reg_out[0]), .QN(KeySchedule_Inst1_GEN_reg_n9) );
  DFF_X1 KeySchedule_Inst1_GEN_reg_Q_reg_1_ ( .D(KeySchedule_Inst1_GEN_reg_n18), .CK(clk), .Q(KeySchedule_Inst1_Reg_out[1]), .QN(
        KeySchedule_Inst1_GEN_reg_n10) );
  DFF_X1 KeySchedule_Inst1_GEN_reg_Q_reg_2_ ( .D(KeySchedule_Inst1_GEN_reg_n19), .CK(clk), .Q(KeySchedule_Inst1_Reg_out[2]), .QN(
        KeySchedule_Inst1_GEN_reg_n11) );
  DFF_X1 KeySchedule_Inst1_GEN_reg_Q_reg_3_ ( .D(KeySchedule_Inst1_GEN_reg_n20), .CK(clk), .Q(KeySchedule_Inst1_Reg_out[3]), .QN(
        KeySchedule_Inst1_GEN_reg_n12) );
  DFF_X1 KeySchedule_Inst1_GEN_reg_Q_reg_4_ ( .D(KeySchedule_Inst1_GEN_reg_n21), .CK(clk), .Q(KeySchedule_Inst1_Reg_out[4]), .QN(
        KeySchedule_Inst1_GEN_reg_n13) );
  DFF_X1 KeySchedule_Inst1_GEN_reg_Q_reg_5_ ( .D(KeySchedule_Inst1_GEN_reg_n22), .CK(clk), .Q(KeySchedule_Inst1_Reg_out[5]), .QN(
        KeySchedule_Inst1_GEN_reg_n14) );
  DFF_X1 KeySchedule_Inst1_GEN_reg_Q_reg_6_ ( .D(KeySchedule_Inst1_GEN_reg_n23), .CK(clk), .Q(KeySchedule_Inst1_Reg_out[6]), .QN(
        KeySchedule_Inst1_GEN_reg_n15) );
  DFF_X1 KeySchedule_Inst1_GEN_reg_Q_reg_7_ ( .D(KeySchedule_Inst1_GEN_reg_n24), .CK(clk), .Q(KeySchedule_Inst1_Reg_out[7]), .QN(
        KeySchedule_Inst1_GEN_reg_n16) );
  OAI21_X1 KeySchedule_Inst1_GEN_reg2_U18 ( .B1(KeySchedule_Inst1_GEN_reg2_n49), .B2(KeySchedule_Inst1_GEN_reg2_n40), .A(KeySchedule_Inst1_GEN_reg2_n57), 
        .ZN(KeySchedule_Inst1_GEN_reg2_n32) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg2_U17 ( .A1(KeySchedule_Inst1_GEN_reg2_n49), .A2(StateIn2[0]), .ZN(KeySchedule_Inst1_GEN_reg2_n57) );
  OAI21_X1 KeySchedule_Inst1_GEN_reg2_U16 ( .B1(KeySchedule_Inst1_GEN_reg2_n49), .B2(KeySchedule_Inst1_GEN_reg2_n39), .A(KeySchedule_Inst1_GEN_reg2_n56), 
        .ZN(KeySchedule_Inst1_GEN_reg2_n31) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg2_U15 ( .A1(KeySchedule_Inst1_GEN_reg2_n49), .A2(StateIn2[1]), .ZN(KeySchedule_Inst1_GEN_reg2_n56) );
  OAI21_X1 KeySchedule_Inst1_GEN_reg2_U14 ( .B1(KeySchedule_Inst1_GEN_reg2_n49), .B2(KeySchedule_Inst1_GEN_reg2_n38), .A(KeySchedule_Inst1_GEN_reg2_n55), 
        .ZN(KeySchedule_Inst1_GEN_reg2_n30) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg2_U13 ( .A1(KeySchedule_Inst1_GEN_reg2_n49), .A2(StateIn2[2]), .ZN(KeySchedule_Inst1_GEN_reg2_n55) );
  OAI21_X1 KeySchedule_Inst1_GEN_reg2_U12 ( .B1(KeySchedule_Inst1_GEN_reg2_n49), .B2(KeySchedule_Inst1_GEN_reg2_n37), .A(KeySchedule_Inst1_GEN_reg2_n54), 
        .ZN(KeySchedule_Inst1_GEN_reg2_n29) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg2_U11 ( .A1(KeySchedule_Inst1_GEN_reg2_n49), .A2(StateIn2[3]), .ZN(KeySchedule_Inst1_GEN_reg2_n54) );
  OAI21_X1 KeySchedule_Inst1_GEN_reg2_U10 ( .B1(KeySchedule_Inst1_GEN_reg2_n49), .B2(KeySchedule_Inst1_GEN_reg2_n36), .A(KeySchedule_Inst1_GEN_reg2_n53), 
        .ZN(KeySchedule_Inst1_GEN_reg2_n28) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg2_U9 ( .A1(KeySchedule_Inst1_GEN_reg2_n49), 
        .A2(StateIn2[4]), .ZN(KeySchedule_Inst1_GEN_reg2_n53) );
  OAI21_X1 KeySchedule_Inst1_GEN_reg2_U8 ( .B1(KeySchedule_Inst1_GEN_reg2_n49), 
        .B2(KeySchedule_Inst1_GEN_reg2_n35), .A(KeySchedule_Inst1_GEN_reg2_n52), .ZN(KeySchedule_Inst1_GEN_reg2_n27) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg2_U7 ( .A1(KeySchedule_Inst1_GEN_reg2_n49), 
        .A2(StateIn2[5]), .ZN(KeySchedule_Inst1_GEN_reg2_n52) );
  OAI21_X1 KeySchedule_Inst1_GEN_reg2_U6 ( .B1(KeySchedule_Inst1_GEN_reg2_n49), 
        .B2(KeySchedule_Inst1_GEN_reg2_n34), .A(KeySchedule_Inst1_GEN_reg2_n51), .ZN(KeySchedule_Inst1_GEN_reg2_n26) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg2_U5 ( .A1(KeySchedule_Inst1_GEN_reg2_n49), 
        .A2(StateIn2[6]), .ZN(KeySchedule_Inst1_GEN_reg2_n51) );
  OAI21_X1 KeySchedule_Inst1_GEN_reg2_U4 ( .B1(KeySchedule_Inst1_GEN_reg2_n49), 
        .B2(KeySchedule_Inst1_GEN_reg2_n33), .A(KeySchedule_Inst1_GEN_reg2_n50), .ZN(KeySchedule_Inst1_GEN_reg2_n25) );
  NAND2_X1 KeySchedule_Inst1_GEN_reg2_U3 ( .A1(KeySchedule_Inst1_GEN_reg2_n49), 
        .A2(StateIn2[7]), .ZN(KeySchedule_Inst1_GEN_reg2_n50) );
  BUF_X1 KeySchedule_Inst1_GEN_reg2_U2 ( .A(KeyScheduleRegisterEN), .Z(
        KeySchedule_Inst1_GEN_reg2_n49) );
  DFF_X1 KeySchedule_Inst1_GEN_reg2_Q_reg_0_ ( .D(
        KeySchedule_Inst1_GEN_reg2_n32), .CK(clk), .Q(
        KeySchedule_Inst1_S_key2_reg[0]), .QN(KeySchedule_Inst1_GEN_reg2_n40)
         );
  DFF_X1 KeySchedule_Inst1_GEN_reg2_Q_reg_1_ ( .D(
        KeySchedule_Inst1_GEN_reg2_n31), .CK(clk), .Q(
        KeySchedule_Inst1_S_key2_reg[1]), .QN(KeySchedule_Inst1_GEN_reg2_n39)
         );
  DFF_X1 KeySchedule_Inst1_GEN_reg2_Q_reg_2_ ( .D(
        KeySchedule_Inst1_GEN_reg2_n30), .CK(clk), .Q(
        KeySchedule_Inst1_S_key2_reg[2]), .QN(KeySchedule_Inst1_GEN_reg2_n38)
         );
  DFF_X1 KeySchedule_Inst1_GEN_reg2_Q_reg_3_ ( .D(
        KeySchedule_Inst1_GEN_reg2_n29), .CK(clk), .Q(
        KeySchedule_Inst1_S_key2_reg[3]), .QN(KeySchedule_Inst1_GEN_reg2_n37)
         );
  DFF_X1 KeySchedule_Inst1_GEN_reg2_Q_reg_4_ ( .D(
        KeySchedule_Inst1_GEN_reg2_n28), .CK(clk), .Q(
        KeySchedule_Inst1_S_key2_reg[4]), .QN(KeySchedule_Inst1_GEN_reg2_n36)
         );
  DFF_X1 KeySchedule_Inst1_GEN_reg2_Q_reg_5_ ( .D(
        KeySchedule_Inst1_GEN_reg2_n27), .CK(clk), .Q(
        KeySchedule_Inst1_S_key2_reg[5]), .QN(KeySchedule_Inst1_GEN_reg2_n35)
         );
  DFF_X1 KeySchedule_Inst1_GEN_reg2_Q_reg_6_ ( .D(
        KeySchedule_Inst1_GEN_reg2_n26), .CK(clk), .Q(
        KeySchedule_Inst1_S_key2_reg[6]), .QN(KeySchedule_Inst1_GEN_reg2_n34)
         );
  DFF_X1 KeySchedule_Inst1_GEN_reg2_Q_reg_7_ ( .D(
        KeySchedule_Inst1_GEN_reg2_n25), .CK(clk), .Q(
        KeySchedule_Inst1_S_key2_reg[7]), .QN(KeySchedule_Inst1_GEN_reg2_n33)
         );
  INV_X1 DataPath_Registers_Inst1_U279 ( .A(DataPath_Registers_Inst1_n529), 
        .ZN(DataPath_Registers_Inst1_n6) );
  OAI22_X1 DataPath_Registers_Inst1_U278 ( .A1(DataPath_Registers_Inst1_n365), 
        .A2(DataPath_Registers_Inst1_n528), .B1(DataPath_Registers_Inst1_n201), 
        .B2(DataPath_Registers_Inst1_n361), .ZN(DataPath_Registers_Inst1_n529)
         );
  XOR2_X1 DataPath_Registers_Inst1_U277 ( .A(DataPath_Registers_Inst1_n527), 
        .B(DataPath_Registers_Inst1_n526), .Z(DataPath_Registers_Inst1_out4[7]) );
  XOR2_X1 DataPath_Registers_Inst1_U276 ( .A(DataPath_Registers_Inst1_n525), 
        .B(DataPath_Registers_Inst1_n524), .Z(DataPath_Registers_Inst1_out4[6]) );
  XOR2_X1 DataPath_Registers_Inst1_U275 ( .A(DataPath_Registers_Inst1_n523), 
        .B(DataPath_Registers_Inst1_n522), .Z(DataPath_Registers_Inst1_out4[5]) );
  XNOR2_X1 DataPath_Registers_Inst1_U274 ( .A(DataPath_Registers_Inst1_n521), 
        .B(DataPath_Registers_Inst1_n520), .ZN(
        DataPath_Registers_Inst1_out4[4]) );
  XNOR2_X1 DataPath_Registers_Inst1_U273 ( .A(DataPath_Registers_Inst1_n519), 
        .B(DataPath_Registers_Inst1_n518), .ZN(
        DataPath_Registers_Inst1_out4[3]) );
  XOR2_X1 DataPath_Registers_Inst1_U272 ( .A(DataPath_Registers_Inst1_n517), 
        .B(DataPath_Registers_Inst1_n516), .Z(DataPath_Registers_Inst1_out4[2]) );
  XNOR2_X1 DataPath_Registers_Inst1_U271 ( .A(DataPath_Registers_Inst1_n515), 
        .B(DataPath_Registers_Inst1_n514), .ZN(
        DataPath_Registers_Inst1_out4[1]) );
  XOR2_X1 DataPath_Registers_Inst1_U270 ( .A(DataPath_Registers_Inst1_n513), 
        .B(DataPath_Registers_Inst1_n528), .Z(DataPath_Registers_Inst1_out4[0]) );
  XNOR2_X1 DataPath_Registers_Inst1_U269 ( .A(DataPath_Registers_Inst1_n512), 
        .B(DataPath_Registers_Inst1_n511), .ZN(
        DataPath_Registers_Inst1_out3[7]) );
  XNOR2_X1 DataPath_Registers_Inst1_U268 ( .A(DataPath_Registers_Inst1_n510), 
        .B(DataPath_Registers_Inst1_n509), .ZN(
        DataPath_Registers_Inst1_out3[6]) );
  XNOR2_X1 DataPath_Registers_Inst1_U267 ( .A(DataPath_Registers_Inst1_n508), 
        .B(DataPath_Registers_Inst1_n507), .ZN(
        DataPath_Registers_Inst1_out3[5]) );
  XOR2_X1 DataPath_Registers_Inst1_U266 ( .A(DataPath_Registers_Inst1_n506), 
        .B(DataPath_Registers_Inst1_n505), .Z(DataPath_Registers_Inst1_out3[4]) );
  XOR2_X1 DataPath_Registers_Inst1_U265 ( .A(DataPath_Registers_Inst1_n504), 
        .B(DataPath_Registers_Inst1_n503), .Z(DataPath_Registers_Inst1_out3[3]) );
  XNOR2_X1 DataPath_Registers_Inst1_U264 ( .A(DataPath_Registers_Inst1_n502), 
        .B(DataPath_Registers_Inst1_n501), .ZN(
        DataPath_Registers_Inst1_out3[2]) );
  XOR2_X1 DataPath_Registers_Inst1_U263 ( .A(DataPath_Registers_Inst1_n500), 
        .B(DataPath_Registers_Inst1_n499), .Z(DataPath_Registers_Inst1_out3[1]) );
  XNOR2_X1 DataPath_Registers_Inst1_U262 ( .A(DataPath_Registers_Inst1_n498), 
        .B(DataPath_Registers_Inst1_n497), .ZN(
        DataPath_Registers_Inst1_out3[0]) );
  XNOR2_X1 DataPath_Registers_Inst1_U261 ( .A(DataPath_Registers_Inst1_n496), 
        .B(DataPath_Registers_Inst1_n512), .ZN(
        DataPath_Registers_Inst1_out2[7]) );
  XNOR2_X1 DataPath_Registers_Inst1_U260 ( .A(DataPath_Registers_Inst1_n495), 
        .B(DataPath_Registers_Inst1_n526), .ZN(DataPath_Registers_Inst1_n512)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U259 ( .A(DataPath_Registers_Inst1_n494), 
        .B(DataPath_Registers_Inst1_n510), .ZN(
        DataPath_Registers_Inst1_out2[6]) );
  XNOR2_X1 DataPath_Registers_Inst1_U258 ( .A(DataPath_Registers_Inst1_n493), 
        .B(DataPath_Registers_Inst1_n524), .ZN(DataPath_Registers_Inst1_n510)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U257 ( .A(DataPath_Registers_Inst1_n492), 
        .B(DataPath_Registers_Inst1_n508), .ZN(
        DataPath_Registers_Inst1_out2[5]) );
  XNOR2_X1 DataPath_Registers_Inst1_U256 ( .A(DataPath_Registers_Inst1_n491), 
        .B(DataPath_Registers_Inst1_n522), .ZN(DataPath_Registers_Inst1_n508)
         );
  XOR2_X1 DataPath_Registers_Inst1_U255 ( .A(DataPath_Registers_Inst1_n490), 
        .B(DataPath_Registers_Inst1_n505), .Z(DataPath_Registers_Inst1_out2[4]) );
  XNOR2_X1 DataPath_Registers_Inst1_U254 ( .A(DataPath_Registers_Inst1_n489), 
        .B(DataPath_Registers_Inst1_n520), .ZN(DataPath_Registers_Inst1_n505)
         );
  XOR2_X1 DataPath_Registers_Inst1_U253 ( .A(DataPath_Registers_Inst1_n488), 
        .B(DataPath_Registers_Inst1_n503), .Z(DataPath_Registers_Inst1_out2[3]) );
  XNOR2_X1 DataPath_Registers_Inst1_U252 ( .A(DataPath_Registers_Inst1_n487), 
        .B(DataPath_Registers_Inst1_n518), .ZN(DataPath_Registers_Inst1_n503)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U251 ( .A(DataPath_Registers_Inst1_n486), 
        .B(DataPath_Registers_Inst1_n502), .ZN(
        DataPath_Registers_Inst1_out2[2]) );
  XNOR2_X1 DataPath_Registers_Inst1_U250 ( .A(DataPath_Registers_Inst1_n485), 
        .B(DataPath_Registers_Inst1_n516), .ZN(DataPath_Registers_Inst1_n502)
         );
  XOR2_X1 DataPath_Registers_Inst1_U249 ( .A(DataPath_Registers_Inst1_n484), 
        .B(DataPath_Registers_Inst1_n499), .Z(DataPath_Registers_Inst1_out2[1]) );
  XNOR2_X1 DataPath_Registers_Inst1_U248 ( .A(DataPath_Registers_Inst1_n483), 
        .B(DataPath_Registers_Inst1_n514), .ZN(DataPath_Registers_Inst1_n499)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U247 ( .A(DataPath_Registers_Inst1_n482), 
        .B(DataPath_Registers_Inst1_n498), .ZN(
        DataPath_Registers_Inst1_out2[0]) );
  XNOR2_X1 DataPath_Registers_Inst1_U246 ( .A(DataPath_Registers_Inst1_n481), 
        .B(DataPath_Registers_Inst1_n528), .ZN(DataPath_Registers_Inst1_n498)
         );
  OAI21_X1 DataPath_Registers_Inst1_U245 ( .B1(DataPath_Registers_Inst1_n245), 
        .B2(DataPath_Registers_Inst1_n480), .A(DataPath_Registers_Inst1_n479), 
        .ZN(DataPath_Registers_Inst1_n528) );
  AOI21_X1 DataPath_Registers_Inst1_U244 ( .B1(DataPath_Registers_Inst1_n353), 
        .B2(DataPath_Registers_Inst1_S6_0_), .A(DataPath_Registers_Inst1_n478), 
        .ZN(DataPath_Registers_Inst1_n479) );
  AOI221_X1 DataPath_Registers_Inst1_U243 ( .B1(
        DataPath_Registers_Inst1_in3_7_), .B2(DataPath_Registers_Inst1_n477), 
        .C1(DataPath_Registers_Inst1_n476), .C2(DataPath_Registers_Inst1_n475), 
        .A(DataPath_Registers_Inst1_n474), .ZN(DataPath_Registers_Inst1_n478)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U242 ( .A(DataPath_Registers_Inst1_n527), 
        .B(DataPath_Registers_Inst1_n495), .ZN(
        DataPath_Registers_Inst1_out1[7]) );
  XOR2_X1 DataPath_Registers_Inst1_U241 ( .A(DataPath_Registers_Inst1_n496), 
        .B(DataPath_Registers_Inst1_n511), .Z(DataPath_Registers_Inst1_n527)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U240 ( .A(DataPath_Registers_Inst1_n525), 
        .B(DataPath_Registers_Inst1_n493), .ZN(
        DataPath_Registers_Inst1_out1[6]) );
  XOR2_X1 DataPath_Registers_Inst1_U239 ( .A(DataPath_Registers_Inst1_n494), 
        .B(DataPath_Registers_Inst1_n509), .Z(DataPath_Registers_Inst1_n525)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U238 ( .A(DataPath_Registers_Inst1_n523), 
        .B(DataPath_Registers_Inst1_n491), .ZN(
        DataPath_Registers_Inst1_out1[5]) );
  XOR2_X1 DataPath_Registers_Inst1_U237 ( .A(DataPath_Registers_Inst1_n492), 
        .B(DataPath_Registers_Inst1_n507), .Z(DataPath_Registers_Inst1_n523)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U236 ( .A(DataPath_Registers_Inst1_n521), 
        .B(DataPath_Registers_Inst1_n489), .ZN(
        DataPath_Registers_Inst1_out1[4]) );
  XOR2_X1 DataPath_Registers_Inst1_U235 ( .A(DataPath_Registers_Inst1_n506), 
        .B(DataPath_Registers_Inst1_n490), .Z(DataPath_Registers_Inst1_n521)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U234 ( .A(DataPath_Registers_Inst1_n519), 
        .B(DataPath_Registers_Inst1_n487), .ZN(
        DataPath_Registers_Inst1_out1[3]) );
  XOR2_X1 DataPath_Registers_Inst1_U233 ( .A(DataPath_Registers_Inst1_n504), 
        .B(DataPath_Registers_Inst1_n488), .Z(DataPath_Registers_Inst1_n519)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U232 ( .A(DataPath_Registers_Inst1_n517), 
        .B(DataPath_Registers_Inst1_n485), .ZN(
        DataPath_Registers_Inst1_out1[2]) );
  XOR2_X1 DataPath_Registers_Inst1_U231 ( .A(DataPath_Registers_Inst1_n486), 
        .B(DataPath_Registers_Inst1_n501), .Z(DataPath_Registers_Inst1_n517)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U230 ( .A(DataPath_Registers_Inst1_n515), 
        .B(DataPath_Registers_Inst1_n483), .ZN(
        DataPath_Registers_Inst1_out1[1]) );
  XOR2_X1 DataPath_Registers_Inst1_U229 ( .A(DataPath_Registers_Inst1_n500), 
        .B(DataPath_Registers_Inst1_n484), .Z(DataPath_Registers_Inst1_n515)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U228 ( .A(DataPath_Registers_Inst1_n513), 
        .B(DataPath_Registers_Inst1_n481), .ZN(
        DataPath_Registers_Inst1_out1[0]) );
  XOR2_X1 DataPath_Registers_Inst1_U227 ( .A(DataPath_Registers_Inst1_n482), 
        .B(DataPath_Registers_Inst1_n497), .Z(DataPath_Registers_Inst1_n513)
         );
  OAI21_X1 DataPath_Registers_Inst1_U226 ( .B1(DataPath_Registers_Inst1_n359), 
        .B2(DataPath_Registers_Inst1_n268), .A(DataPath_Registers_Inst1_n473), 
        .ZN(DataPath_Registers_Inst1_n324) );
  NAND2_X1 DataPath_Registers_Inst1_U225 ( .A1(DataPath_Registers_Inst1_n361), 
        .A2(DataPath_Registers_Inst1_S8_in[0]), .ZN(
        DataPath_Registers_Inst1_n473) );
  INV_X1 DataPath_Registers_Inst1_U224 ( .A(DataPath_Registers_Inst1_n472), 
        .ZN(DataPath_Registers_Inst1_n323) );
  OAI22_X1 DataPath_Registers_Inst1_U223 ( .A1(DataPath_Registers_Inst1_n365), 
        .A2(DataPath_Registers_Inst1_n526), .B1(DataPath_Registers_Inst1_n203), 
        .B2(DataPath_Registers_Inst1_n360), .ZN(DataPath_Registers_Inst1_n472)
         );
  OAI222_X1 DataPath_Registers_Inst1_U222 ( .A1(DataPath_Registers_Inst1_n471), 
        .A2(DataPath_Registers_Inst1_n474), .B1(DataPath_Registers_Inst1_n480), 
        .B2(DataPath_Registers_Inst1_n266), .C1(DataPath_Registers_Inst1_n354), 
        .C2(DataPath_Registers_Inst1_n470), .ZN(DataPath_Registers_Inst1_n526)
         );
  INV_X1 DataPath_Registers_Inst1_U221 ( .A(DataPath_Registers_Inst1_S6_7_), 
        .ZN(DataPath_Registers_Inst1_n470) );
  XNOR2_X1 DataPath_Registers_Inst1_U220 ( .A(DataPath_Registers_Inst1_in3_6_), 
        .B(DataPath_Registers_Inst1_n469), .ZN(DataPath_Registers_Inst1_n471)
         );
  AOI22_X1 DataPath_Registers_Inst1_U219 ( .A1(DataPath_Registers_Inst1_in2_7_), .A2(DataPath_Registers_Inst1_in2_6_), .B1(DataPath_Registers_Inst1_n468), 
        .B2(DataPath_Registers_Inst1_n467), .ZN(DataPath_Registers_Inst1_n469)
         );
  AOI22_X1 DataPath_Registers_Inst1_U218 ( .A1(DataPath_Registers_Inst1_n359), 
        .A2(DataPath_Registers_Inst1_n495), .B1(DataPath_Registers_Inst1_n347), 
        .B2(DataPath_Registers_Inst1_n364), .ZN(DataPath_Registers_Inst1_n322)
         );
  AOI22_X1 DataPath_Registers_Inst1_U217 ( .A1(DataPath_Registers_Inst1_n466), 
        .A2(DataPath_Registers_Inst1_n465), .B1(DataPath_Registers_Inst1_n203), 
        .B2(DataPath_Registers_Inst1_n474), .ZN(DataPath_Registers_Inst1_n495)
         );
  XOR2_X1 DataPath_Registers_Inst1_U216 ( .A(DataPath_Registers_Inst1_n464), 
        .B(DataPath_Registers_Inst1_n468), .Z(DataPath_Registers_Inst1_n465)
         );
  XOR2_X1 DataPath_Registers_Inst1_U215 ( .A(DataPath_Registers_Inst1_n463), 
        .B(DataPath_Registers_Inst1_in1_6_), .Z(DataPath_Registers_Inst1_n464)
         );
  AOI22_X1 DataPath_Registers_Inst1_U214 ( .A1(DataPath_Registers_Inst1_n359), 
        .A2(DataPath_Registers_Inst1_n506), .B1(DataPath_Registers_Inst1_n264), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n321)
         );
  AOI222_X1 DataPath_Registers_Inst1_U213 ( .A1(DataPath_Registers_Inst1_S3_4_), .A2(DataPath_Registers_Inst1_n462), .B1(DataPath_Registers_Inst1_n466), .B2(
        DataPath_Registers_Inst1_n461), .C1(DataPath_Registers_Inst1_n353), 
        .C2(DataPath_Registers_Inst1_S11_4_), .ZN(
        DataPath_Registers_Inst1_n506) );
  XNOR2_X1 DataPath_Registers_Inst1_U212 ( .A(DataPath_Registers_Inst1_n460), 
        .B(DataPath_Registers_Inst1_n459), .ZN(DataPath_Registers_Inst1_n461)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U211 ( .A(DataPath_Registers_Inst1_n458), 
        .B(DataPath_Registers_Inst1_in3_4_), .ZN(DataPath_Registers_Inst1_n460) );
  OAI21_X1 DataPath_Registers_Inst1_U210 ( .B1(DataPath_Registers_Inst1_n359), 
        .B2(DataPath_Registers_Inst1_n262), .A(DataPath_Registers_Inst1_n457), 
        .ZN(DataPath_Registers_Inst1_n320) );
  NAND2_X1 DataPath_Registers_Inst1_U209 ( .A1(DataPath_Registers_Inst1_n361), 
        .A2(DataPath_Registers_Inst1_S12_in[0]), .ZN(
        DataPath_Registers_Inst1_n457) );
  OAI21_X1 DataPath_Registers_Inst1_U208 ( .B1(DataPath_Registers_Inst1_n360), 
        .B2(DataPath_Registers_Inst1_n261), .A(DataPath_Registers_Inst1_n456), 
        .ZN(DataPath_Registers_Inst1_n319) );
  NAND2_X1 DataPath_Registers_Inst1_U207 ( .A1(DataPath_Registers_Inst1_n361), 
        .A2(DataPath_Registers_Inst1_S12_in[1]), .ZN(
        DataPath_Registers_Inst1_n456) );
  OAI21_X1 DataPath_Registers_Inst1_U206 ( .B1(DataPath_Registers_Inst1_n358), 
        .B2(DataPath_Registers_Inst1_n260), .A(DataPath_Registers_Inst1_n455), 
        .ZN(DataPath_Registers_Inst1_n318) );
  NAND2_X1 DataPath_Registers_Inst1_U205 ( .A1(DataPath_Registers_Inst1_n362), 
        .A2(DataPath_Registers_Inst1_S12_in[2]), .ZN(
        DataPath_Registers_Inst1_n455) );
  OAI21_X1 DataPath_Registers_Inst1_U204 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n259), .A(DataPath_Registers_Inst1_n454), 
        .ZN(DataPath_Registers_Inst1_n317) );
  NAND2_X1 DataPath_Registers_Inst1_U203 ( .A1(DataPath_Registers_Inst1_n362), 
        .A2(DataPath_Registers_Inst1_S12_in[3]), .ZN(
        DataPath_Registers_Inst1_n454) );
  OAI21_X1 DataPath_Registers_Inst1_U202 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n258), .A(DataPath_Registers_Inst1_n453), 
        .ZN(DataPath_Registers_Inst1_n316) );
  NAND2_X1 DataPath_Registers_Inst1_U201 ( .A1(DataPath_Registers_Inst1_n362), 
        .A2(DataPath_Registers_Inst1_S12_in[4]), .ZN(
        DataPath_Registers_Inst1_n453) );
  OAI21_X1 DataPath_Registers_Inst1_U200 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n257), .A(DataPath_Registers_Inst1_n452), 
        .ZN(DataPath_Registers_Inst1_n315) );
  NAND2_X1 DataPath_Registers_Inst1_U199 ( .A1(DataPath_Registers_Inst1_n362), 
        .A2(DataPath_Registers_Inst1_S12_in[5]), .ZN(
        DataPath_Registers_Inst1_n452) );
  OAI21_X1 DataPath_Registers_Inst1_U198 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n256), .A(DataPath_Registers_Inst1_n451), 
        .ZN(DataPath_Registers_Inst1_n314) );
  NAND2_X1 DataPath_Registers_Inst1_U197 ( .A1(DataPath_Registers_Inst1_n362), 
        .A2(DataPath_Registers_Inst1_S12_in[6]), .ZN(
        DataPath_Registers_Inst1_n451) );
  OAI21_X1 DataPath_Registers_Inst1_U196 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n255), .A(DataPath_Registers_Inst1_n450), 
        .ZN(DataPath_Registers_Inst1_n313) );
  NAND2_X1 DataPath_Registers_Inst1_U195 ( .A1(DataPath_Registers_Inst1_n363), 
        .A2(DataPath_Registers_Inst1_S12_in[7]), .ZN(
        DataPath_Registers_Inst1_n450) );
  OAI21_X1 DataPath_Registers_Inst1_U194 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n254), .A(DataPath_Registers_Inst1_n449), 
        .ZN(DataPath_Registers_Inst1_n312) );
  NAND2_X1 DataPath_Registers_Inst1_U193 ( .A1(DataPath_Registers_Inst1_n363), 
        .A2(DataPath_Registers_Inst1_S8_in[1]), .ZN(
        DataPath_Registers_Inst1_n449) );
  OAI21_X1 DataPath_Registers_Inst1_U192 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n253), .A(DataPath_Registers_Inst1_n448), 
        .ZN(DataPath_Registers_Inst1_n311) );
  NAND2_X1 DataPath_Registers_Inst1_U191 ( .A1(DataPath_Registers_Inst1_n363), 
        .A2(DataPath_Registers_Inst1_S8_in[2]), .ZN(
        DataPath_Registers_Inst1_n448) );
  OAI21_X1 DataPath_Registers_Inst1_U190 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n252), .A(DataPath_Registers_Inst1_n447), 
        .ZN(DataPath_Registers_Inst1_n310) );
  NAND2_X1 DataPath_Registers_Inst1_U189 ( .A1(DataPath_Registers_Inst1_n363), 
        .A2(DataPath_Registers_Inst1_S8_in[3]), .ZN(
        DataPath_Registers_Inst1_n447) );
  OAI21_X1 DataPath_Registers_Inst1_U188 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n251), .A(DataPath_Registers_Inst1_n446), 
        .ZN(DataPath_Registers_Inst1_n309) );
  NAND2_X1 DataPath_Registers_Inst1_U187 ( .A1(DataPath_Registers_Inst1_n363), 
        .A2(DataPath_Registers_Inst1_S8_in[4]), .ZN(
        DataPath_Registers_Inst1_n446) );
  OAI21_X1 DataPath_Registers_Inst1_U186 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n250), .A(DataPath_Registers_Inst1_n445), 
        .ZN(DataPath_Registers_Inst1_n308) );
  NAND2_X1 DataPath_Registers_Inst1_U185 ( .A1(DataPath_Registers_Inst1_n363), 
        .A2(DataPath_Registers_Inst1_S8_in[5]), .ZN(
        DataPath_Registers_Inst1_n445) );
  OAI21_X1 DataPath_Registers_Inst1_U184 ( .B1(DataPath_Registers_Inst1_n363), 
        .B2(DataPath_Registers_Inst1_n249), .A(DataPath_Registers_Inst1_n444), 
        .ZN(DataPath_Registers_Inst1_n307) );
  NAND2_X1 DataPath_Registers_Inst1_U183 ( .A1(DataPath_Registers_Inst1_n363), 
        .A2(DataPath_Registers_Inst1_S8_in[6]), .ZN(
        DataPath_Registers_Inst1_n444) );
  OAI21_X1 DataPath_Registers_Inst1_U182 ( .B1(DataPath_Registers_Inst1_n356), 
        .B2(DataPath_Registers_Inst1_n248), .A(DataPath_Registers_Inst1_n443), 
        .ZN(DataPath_Registers_Inst1_n306) );
  NAND2_X1 DataPath_Registers_Inst1_U181 ( .A1(DataPath_Registers_Inst1_n363), 
        .A2(DataPath_Registers_Inst1_S8_in[7]), .ZN(
        DataPath_Registers_Inst1_n443) );
  MUX2_X1 DataPath_Registers_Inst1_U180 ( .A(DataPath_Registers_Inst1_S4_in[0]), .B(DataPath_Registers_Inst1_S4_0_), .S(DataPath_Registers_Inst1_n366), .Z(
        DataPath_Registers_Inst1_n305) );
  AOI22_X1 DataPath_Registers_Inst1_U179 ( .A1(DataPath_Registers_Inst1_n358), 
        .A2(DataPath_Registers_Inst1_n482), .B1(DataPath_Registers_Inst1_n246), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n304)
         );
  AOI22_X1 DataPath_Registers_Inst1_U178 ( .A1(DataPath_Registers_Inst1_n352), 
        .A2(StateIn1[0]), .B1(DataPath_Registers_Inst1_S4_0_), .B2(
        DataPath_Registers_Inst1_n354), .ZN(DataPath_Registers_Inst1_n482) );
  AOI22_X1 DataPath_Registers_Inst1_U177 ( .A1(DataPath_Registers_Inst1_n360), 
        .A2(DataPath_Registers_Inst1_n497), .B1(DataPath_Registers_Inst1_n245), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n303)
         );
  AOI22_X1 DataPath_Registers_Inst1_U176 ( .A1(DataPath_Registers_Inst1_n359), 
        .A2(DataPath_Registers_Inst1_n481), .B1(DataPath_Registers_Inst1_n346), 
        .B2(DataPath_Registers_Inst1_n364), .ZN(DataPath_Registers_Inst1_n301)
         );
  AOI22_X1 DataPath_Registers_Inst1_U175 ( .A1(DataPath_Registers_Inst1_n466), 
        .A2(DataPath_Registers_Inst1_n440), .B1(DataPath_Registers_Inst1_n201), 
        .B2(DataPath_Registers_Inst1_n474), .ZN(DataPath_Registers_Inst1_n481)
         );
  AOI22_X1 DataPath_Registers_Inst1_U174 ( .A1(DataPath_Registers_Inst1_in2_7_), .A2(DataPath_Registers_Inst1_n439), .B1(DataPath_Registers_Inst1_n438), .B2(
        DataPath_Registers_Inst1_n467), .ZN(DataPath_Registers_Inst1_n440) );
  OAI21_X1 DataPath_Registers_Inst1_U173 ( .B1(DataPath_Registers_Inst1_n361), 
        .B2(DataPath_Registers_Inst1_n242), .A(DataPath_Registers_Inst1_n437), 
        .ZN(DataPath_Registers_Inst1_n300) );
  NAND2_X1 DataPath_Registers_Inst1_U172 ( .A1(DataPath_Registers_Inst1_n363), 
        .A2(DataPath_Registers_Inst1_S4_in[1]), .ZN(
        DataPath_Registers_Inst1_n437) );
  AOI22_X1 DataPath_Registers_Inst1_U171 ( .A1(DataPath_Registers_Inst1_n359), 
        .A2(DataPath_Registers_Inst1_n484), .B1(DataPath_Registers_Inst1_n241), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n299)
         );
  OAI22_X1 DataPath_Registers_Inst1_U170 ( .A1(DataPath_Registers_Inst1_n354), 
        .A2(StateIn1[1]), .B1(DataPath_Registers_Inst1_S4_1_), .B2(
        DataPath_Registers_Inst1_n353), .ZN(DataPath_Registers_Inst1_n484) );
  AOI22_X1 DataPath_Registers_Inst1_U169 ( .A1(DataPath_Registers_Inst1_n358), 
        .A2(DataPath_Registers_Inst1_n500), .B1(DataPath_Registers_Inst1_n240), 
        .B2(DataPath_Registers_Inst1_n364), .ZN(DataPath_Registers_Inst1_n298)
         );
  AOI222_X1 DataPath_Registers_Inst1_U168 ( .A1(DataPath_Registers_Inst1_S3_1_), .A2(DataPath_Registers_Inst1_n462), .B1(DataPath_Registers_Inst1_n466), .B2(
        DataPath_Registers_Inst1_n436), .C1(DataPath_Registers_Inst1_n353), 
        .C2(DataPath_Registers_Inst1_S11_1_), .ZN(
        DataPath_Registers_Inst1_n500) );
  XOR2_X1 DataPath_Registers_Inst1_U167 ( .A(DataPath_Registers_Inst1_n435), 
        .B(DataPath_Registers_Inst1_n434), .Z(DataPath_Registers_Inst1_n436)
         );
  XOR2_X1 DataPath_Registers_Inst1_U166 ( .A(DataPath_Registers_Inst1_in3_1_), 
        .B(DataPath_Registers_Inst1_n442), .Z(DataPath_Registers_Inst1_n435)
         );
  AOI22_X1 DataPath_Registers_Inst1_U165 ( .A1(DataPath_Registers_Inst1_n359), 
        .A2(DataPath_Registers_Inst1_n514), .B1(DataPath_Registers_Inst1_n350), 
        .B2(DataPath_Registers_Inst1_n364), .ZN(DataPath_Registers_Inst1_n297)
         );
  AOI222_X1 DataPath_Registers_Inst1_U164 ( .A1(DataPath_Registers_Inst1_S2_1_), .A2(DataPath_Registers_Inst1_n462), .B1(DataPath_Registers_Inst1_n466), .B2(
        DataPath_Registers_Inst1_n433), .C1(DataPath_Registers_Inst1_n353), 
        .C2(DataPath_Registers_Inst1_S6_1_), .ZN(DataPath_Registers_Inst1_n514) );
  XNOR2_X1 DataPath_Registers_Inst1_U163 ( .A(DataPath_Registers_Inst1_n432), 
        .B(DataPath_Registers_Inst1_in2_1_), .ZN(DataPath_Registers_Inst1_n433) );
  XOR2_X1 DataPath_Registers_Inst1_U162 ( .A(DataPath_Registers_Inst1_n442), 
        .B(DataPath_Registers_Inst1_n477), .Z(DataPath_Registers_Inst1_n432)
         );
  INV_X1 DataPath_Registers_Inst1_U161 ( .A(DataPath_Registers_Inst1_n475), 
        .ZN(DataPath_Registers_Inst1_n477) );
  XOR2_X1 DataPath_Registers_Inst1_U160 ( .A(DataPath_Registers_Inst1_n476), 
        .B(DataPath_Registers_Inst1_in3_0_), .Z(DataPath_Registers_Inst1_n442)
         );
  AOI22_X1 DataPath_Registers_Inst1_U159 ( .A1(DataPath_Registers_Inst1_n358), 
        .A2(DataPath_Registers_Inst1_n483), .B1(DataPath_Registers_Inst1_n345), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n296)
         );
  AOI22_X1 DataPath_Registers_Inst1_U158 ( .A1(DataPath_Registers_Inst1_n466), 
        .A2(DataPath_Registers_Inst1_n431), .B1(DataPath_Registers_Inst1_n202), 
        .B2(DataPath_Registers_Inst1_n474), .ZN(DataPath_Registers_Inst1_n483)
         );
  XOR2_X1 DataPath_Registers_Inst1_U157 ( .A(DataPath_Registers_Inst1_n430), 
        .B(DataPath_Registers_Inst1_n438), .Z(DataPath_Registers_Inst1_n431)
         );
  XOR2_X1 DataPath_Registers_Inst1_U156 ( .A(DataPath_Registers_Inst1_n475), 
        .B(DataPath_Registers_Inst1_in1_1_), .Z(DataPath_Registers_Inst1_n430)
         );
  XOR2_X1 DataPath_Registers_Inst1_U155 ( .A(DataPath_Registers_Inst1_n467), 
        .B(DataPath_Registers_Inst1_in2_0_), .Z(DataPath_Registers_Inst1_n475)
         );
  MUX2_X1 DataPath_Registers_Inst1_U154 ( .A(DataPath_Registers_Inst1_S4_in[2]), .B(DataPath_Registers_Inst1_S4_2_), .S(DataPath_Registers_Inst1_n366), .Z(
        DataPath_Registers_Inst1_n295) );
  AOI22_X1 DataPath_Registers_Inst1_U153 ( .A1(DataPath_Registers_Inst1_n358), 
        .A2(DataPath_Registers_Inst1_n486), .B1(DataPath_Registers_Inst1_n236), 
        .B2(DataPath_Registers_Inst1_n364), .ZN(DataPath_Registers_Inst1_n294)
         );
  AOI22_X1 DataPath_Registers_Inst1_U152 ( .A1(DataPath_Registers_Inst1_n353), 
        .A2(StateIn1[2]), .B1(DataPath_Registers_Inst1_S4_2_), .B2(
        DataPath_Registers_Inst1_n354), .ZN(DataPath_Registers_Inst1_n486) );
  AOI22_X1 DataPath_Registers_Inst1_U151 ( .A1(DataPath_Registers_Inst1_n357), 
        .A2(DataPath_Registers_Inst1_n501), .B1(DataPath_Registers_Inst1_n235), 
        .B2(DataPath_Registers_Inst1_n364), .ZN(DataPath_Registers_Inst1_n293)
         );
  AOI222_X1 DataPath_Registers_Inst1_U150 ( .A1(DataPath_Registers_Inst1_n429), 
        .A2(DataPath_Registers_Inst1_n466), .B1(DataPath_Registers_Inst1_n462), 
        .B2(DataPath_Registers_Inst1_S3_2_), .C1(DataPath_Registers_Inst1_n353), .C2(DataPath_Registers_Inst1_S11_2_), .ZN(DataPath_Registers_Inst1_n501) );
  XOR2_X1 DataPath_Registers_Inst1_U149 ( .A(DataPath_Registers_Inst1_in4_1_), 
        .B(DataPath_Registers_Inst1_n428), .Z(DataPath_Registers_Inst1_n429)
         );
  XOR2_X1 DataPath_Registers_Inst1_U148 ( .A(DataPath_Registers_Inst1_in3_1_), 
        .B(DataPath_Registers_Inst1_in3_2_), .Z(DataPath_Registers_Inst1_n428)
         );
  INV_X1 DataPath_Registers_Inst1_U147 ( .A(DataPath_Registers_Inst1_n427), 
        .ZN(DataPath_Registers_Inst1_n292) );
  OAI22_X1 DataPath_Registers_Inst1_U146 ( .A1(DataPath_Registers_Inst1_n365), 
        .A2(DataPath_Registers_Inst1_n516), .B1(DataPath_Registers_Inst1_n212), 
        .B2(DataPath_Registers_Inst1_n360), .ZN(DataPath_Registers_Inst1_n427)
         );
  OAI222_X1 DataPath_Registers_Inst1_U145 ( .A1(DataPath_Registers_Inst1_n426), 
        .A2(DataPath_Registers_Inst1_n474), .B1(DataPath_Registers_Inst1_n480), 
        .B2(DataPath_Registers_Inst1_n235), .C1(DataPath_Registers_Inst1_n354), 
        .C2(DataPath_Registers_Inst1_n425), .ZN(DataPath_Registers_Inst1_n516)
         );
  INV_X1 DataPath_Registers_Inst1_U144 ( .A(DataPath_Registers_Inst1_S6_2_), 
        .ZN(DataPath_Registers_Inst1_n425) );
  XNOR2_X1 DataPath_Registers_Inst1_U143 ( .A(DataPath_Registers_Inst1_in2_1_), 
        .B(DataPath_Registers_Inst1_n424), .ZN(DataPath_Registers_Inst1_n426)
         );
  XOR2_X1 DataPath_Registers_Inst1_U142 ( .A(DataPath_Registers_Inst1_in3_1_), 
        .B(DataPath_Registers_Inst1_in2_2_), .Z(DataPath_Registers_Inst1_n424)
         );
  AOI22_X1 DataPath_Registers_Inst1_U141 ( .A1(DataPath_Registers_Inst1_n358), 
        .A2(DataPath_Registers_Inst1_n485), .B1(DataPath_Registers_Inst1_n344), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n291)
         );
  AOI22_X1 DataPath_Registers_Inst1_U140 ( .A1(DataPath_Registers_Inst1_n466), 
        .A2(DataPath_Registers_Inst1_n423), .B1(DataPath_Registers_Inst1_n212), 
        .B2(DataPath_Registers_Inst1_n474), .ZN(DataPath_Registers_Inst1_n485)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U139 ( .A(DataPath_Registers_Inst1_n422), 
        .B(DataPath_Registers_Inst1_in2_1_), .ZN(DataPath_Registers_Inst1_n423) );
  XNOR2_X1 DataPath_Registers_Inst1_U138 ( .A(DataPath_Registers_Inst1_in1_1_), 
        .B(DataPath_Registers_Inst1_in1_2_), .ZN(DataPath_Registers_Inst1_n422) );
  OAI21_X1 DataPath_Registers_Inst1_U137 ( .B1(DataPath_Registers_Inst1_n356), 
        .B2(DataPath_Registers_Inst1_n232), .A(DataPath_Registers_Inst1_n421), 
        .ZN(DataPath_Registers_Inst1_n290) );
  NAND2_X1 DataPath_Registers_Inst1_U136 ( .A1(DataPath_Registers_Inst1_n363), 
        .A2(DataPath_Registers_Inst1_S4_in[3]), .ZN(
        DataPath_Registers_Inst1_n421) );
  AOI22_X1 DataPath_Registers_Inst1_U135 ( .A1(DataPath_Registers_Inst1_n362), 
        .A2(DataPath_Registers_Inst1_n488), .B1(DataPath_Registers_Inst1_n231), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n289)
         );
  OAI22_X1 DataPath_Registers_Inst1_U134 ( .A1(DataPath_Registers_Inst1_n354), 
        .A2(StateIn1[3]), .B1(DataPath_Registers_Inst1_S4_3_), .B2(
        DataPath_Registers_Inst1_n353), .ZN(DataPath_Registers_Inst1_n488) );
  AOI22_X1 DataPath_Registers_Inst1_U133 ( .A1(DataPath_Registers_Inst1_n362), 
        .A2(DataPath_Registers_Inst1_n504), .B1(DataPath_Registers_Inst1_n230), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n288)
         );
  AOI222_X1 DataPath_Registers_Inst1_U132 ( .A1(DataPath_Registers_Inst1_S3_3_), .A2(DataPath_Registers_Inst1_n462), .B1(DataPath_Registers_Inst1_n466), .B2(
        DataPath_Registers_Inst1_n420), .C1(DataPath_Registers_Inst1_n353), 
        .C2(DataPath_Registers_Inst1_S11_3_), .ZN(
        DataPath_Registers_Inst1_n504) );
  XNOR2_X1 DataPath_Registers_Inst1_U131 ( .A(DataPath_Registers_Inst1_n419), 
        .B(DataPath_Registers_Inst1_n418), .ZN(DataPath_Registers_Inst1_n420)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U130 ( .A(DataPath_Registers_Inst1_n458), 
        .B(DataPath_Registers_Inst1_in3_2_), .ZN(DataPath_Registers_Inst1_n419) );
  AOI22_X1 DataPath_Registers_Inst1_U129 ( .A1(DataPath_Registers_Inst1_n361), 
        .A2(DataPath_Registers_Inst1_n518), .B1(DataPath_Registers_Inst1_n349), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n287)
         );
  AOI222_X1 DataPath_Registers_Inst1_U128 ( .A1(DataPath_Registers_Inst1_S2_3_), .A2(DataPath_Registers_Inst1_n462), .B1(DataPath_Registers_Inst1_n466), .B2(
        DataPath_Registers_Inst1_n417), .C1(DataPath_Registers_Inst1_n353), 
        .C2(DataPath_Registers_Inst1_S6_3_), .ZN(DataPath_Registers_Inst1_n518) );
  XNOR2_X1 DataPath_Registers_Inst1_U127 ( .A(DataPath_Registers_Inst1_n416), 
        .B(DataPath_Registers_Inst1_n415), .ZN(DataPath_Registers_Inst1_n417)
         );
  XOR2_X1 DataPath_Registers_Inst1_U126 ( .A(DataPath_Registers_Inst1_n476), 
        .B(DataPath_Registers_Inst1_in3_2_), .Z(DataPath_Registers_Inst1_n415)
         );
  XOR2_X1 DataPath_Registers_Inst1_U125 ( .A(DataPath_Registers_Inst1_in2_3_), 
        .B(DataPath_Registers_Inst1_n414), .Z(DataPath_Registers_Inst1_n416)
         );
  AOI22_X1 DataPath_Registers_Inst1_U124 ( .A1(DataPath_Registers_Inst1_n360), 
        .A2(DataPath_Registers_Inst1_n487), .B1(DataPath_Registers_Inst1_n343), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n286)
         );
  AOI22_X1 DataPath_Registers_Inst1_U123 ( .A1(DataPath_Registers_Inst1_n466), 
        .A2(DataPath_Registers_Inst1_n413), .B1(DataPath_Registers_Inst1_n210), 
        .B2(DataPath_Registers_Inst1_n474), .ZN(DataPath_Registers_Inst1_n487)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U122 ( .A(DataPath_Registers_Inst1_n412), 
        .B(DataPath_Registers_Inst1_in1_2_), .ZN(DataPath_Registers_Inst1_n413) );
  XNOR2_X1 DataPath_Registers_Inst1_U121 ( .A(DataPath_Registers_Inst1_n414), 
        .B(DataPath_Registers_Inst1_n411), .ZN(DataPath_Registers_Inst1_n412)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U120 ( .A(DataPath_Registers_Inst1_n467), 
        .B(DataPath_Registers_Inst1_in2_2_), .ZN(DataPath_Registers_Inst1_n414) );
  OAI21_X1 DataPath_Registers_Inst1_U119 ( .B1(DataPath_Registers_Inst1_n358), 
        .B2(DataPath_Registers_Inst1_n227), .A(DataPath_Registers_Inst1_n410), 
        .ZN(DataPath_Registers_Inst1_n285) );
  NAND2_X1 DataPath_Registers_Inst1_U118 ( .A1(DataPath_Registers_Inst1_n361), 
        .A2(DataPath_Registers_Inst1_S4_in[4]), .ZN(
        DataPath_Registers_Inst1_n410) );
  AOI22_X1 DataPath_Registers_Inst1_U117 ( .A1(DataPath_Registers_Inst1_n357), 
        .A2(DataPath_Registers_Inst1_n490), .B1(DataPath_Registers_Inst1_n263), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n284)
         );
  OAI22_X1 DataPath_Registers_Inst1_U116 ( .A1(DataPath_Registers_Inst1_n354), 
        .A2(StateIn1[4]), .B1(DataPath_Registers_Inst1_S4_4_), .B2(
        DataPath_Registers_Inst1_n353), .ZN(DataPath_Registers_Inst1_n490) );
  MUX2_X1 DataPath_Registers_Inst1_U115 ( .A(DataPath_Registers_Inst1_S4_in[5]), .B(DataPath_Registers_Inst1_S4_5_), .S(DataPath_Registers_Inst1_n366), .Z(
        DataPath_Registers_Inst1_n283) );
  AOI22_X1 DataPath_Registers_Inst1_U114 ( .A1(DataPath_Registers_Inst1_n357), 
        .A2(DataPath_Registers_Inst1_n492), .B1(DataPath_Registers_Inst1_n225), 
        .B2(DataPath_Registers_Inst1_n364), .ZN(DataPath_Registers_Inst1_n282)
         );
  AOI22_X1 DataPath_Registers_Inst1_U113 ( .A1(DataPath_Registers_Inst1_n353), 
        .A2(StateIn1[5]), .B1(DataPath_Registers_Inst1_S4_5_), .B2(
        DataPath_Registers_Inst1_n354), .ZN(DataPath_Registers_Inst1_n492) );
  AOI22_X1 DataPath_Registers_Inst1_U112 ( .A1(DataPath_Registers_Inst1_n357), 
        .A2(DataPath_Registers_Inst1_n507), .B1(DataPath_Registers_Inst1_n224), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n281)
         );
  AOI222_X1 DataPath_Registers_Inst1_U111 ( .A1(DataPath_Registers_Inst1_n409), 
        .A2(DataPath_Registers_Inst1_n466), .B1(DataPath_Registers_Inst1_n462), 
        .B2(DataPath_Registers_Inst1_S3_5_), .C1(DataPath_Registers_Inst1_n353), .C2(DataPath_Registers_Inst1_S11_5_), .ZN(DataPath_Registers_Inst1_n507) );
  XOR2_X1 DataPath_Registers_Inst1_U110 ( .A(DataPath_Registers_Inst1_in4_4_), 
        .B(DataPath_Registers_Inst1_n408), .Z(DataPath_Registers_Inst1_n409)
         );
  XOR2_X1 DataPath_Registers_Inst1_U109 ( .A(DataPath_Registers_Inst1_in3_4_), 
        .B(DataPath_Registers_Inst1_in3_5_), .Z(DataPath_Registers_Inst1_n408)
         );
  INV_X1 DataPath_Registers_Inst1_U108 ( .A(DataPath_Registers_Inst1_n407), 
        .ZN(DataPath_Registers_Inst1_n280) );
  OAI22_X1 DataPath_Registers_Inst1_U107 ( .A1(DataPath_Registers_Inst1_n365), 
        .A2(DataPath_Registers_Inst1_n522), .B1(DataPath_Registers_Inst1_n208), 
        .B2(DataPath_Registers_Inst1_n360), .ZN(DataPath_Registers_Inst1_n407)
         );
  OAI222_X1 DataPath_Registers_Inst1_U106 ( .A1(DataPath_Registers_Inst1_n406), 
        .A2(DataPath_Registers_Inst1_n474), .B1(DataPath_Registers_Inst1_n480), 
        .B2(DataPath_Registers_Inst1_n224), .C1(DataPath_Registers_Inst1_n354), 
        .C2(DataPath_Registers_Inst1_n405), .ZN(DataPath_Registers_Inst1_n522)
         );
  INV_X1 DataPath_Registers_Inst1_U105 ( .A(DataPath_Registers_Inst1_S6_5_), 
        .ZN(DataPath_Registers_Inst1_n405) );
  XNOR2_X1 DataPath_Registers_Inst1_U104 ( .A(DataPath_Registers_Inst1_in2_5_), 
        .B(DataPath_Registers_Inst1_n404), .ZN(DataPath_Registers_Inst1_n406)
         );
  XOR2_X1 DataPath_Registers_Inst1_U103 ( .A(DataPath_Registers_Inst1_in3_4_), 
        .B(DataPath_Registers_Inst1_in2_4_), .Z(DataPath_Registers_Inst1_n404)
         );
  AOI22_X1 DataPath_Registers_Inst1_U102 ( .A1(DataPath_Registers_Inst1_n357), 
        .A2(DataPath_Registers_Inst1_n491), .B1(DataPath_Registers_Inst1_n342), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n279)
         );
  AOI22_X1 DataPath_Registers_Inst1_U101 ( .A1(DataPath_Registers_Inst1_n466), 
        .A2(DataPath_Registers_Inst1_n403), .B1(DataPath_Registers_Inst1_n208), 
        .B2(DataPath_Registers_Inst1_n474), .ZN(DataPath_Registers_Inst1_n491)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U100 ( .A(DataPath_Registers_Inst1_n402), 
        .B(DataPath_Registers_Inst1_in1_5_), .ZN(DataPath_Registers_Inst1_n403) );
  XNOR2_X1 DataPath_Registers_Inst1_U99 ( .A(DataPath_Registers_Inst1_in1_4_), 
        .B(DataPath_Registers_Inst1_in2_4_), .ZN(DataPath_Registers_Inst1_n402) );
  MUX2_X1 DataPath_Registers_Inst1_U98 ( .A(DataPath_Registers_Inst1_S4_in[6]), 
        .B(DataPath_Registers_Inst1_S4_6_), .S(DataPath_Registers_Inst1_n366), 
        .Z(DataPath_Registers_Inst1_n278) );
  AOI22_X1 DataPath_Registers_Inst1_U97 ( .A1(DataPath_Registers_Inst1_n357), 
        .A2(DataPath_Registers_Inst1_n494), .B1(DataPath_Registers_Inst1_n220), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n277)
         );
  AOI22_X1 DataPath_Registers_Inst1_U96 ( .A1(DataPath_Registers_Inst1_n353), 
        .A2(StateIn1[6]), .B1(DataPath_Registers_Inst1_S4_6_), .B2(
        DataPath_Registers_Inst1_n354), .ZN(DataPath_Registers_Inst1_n494) );
  AOI22_X1 DataPath_Registers_Inst1_U95 ( .A1(DataPath_Registers_Inst1_n356), 
        .A2(DataPath_Registers_Inst1_n509), .B1(DataPath_Registers_Inst1_n219), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n276)
         );
  AOI222_X1 DataPath_Registers_Inst1_U94 ( .A1(DataPath_Registers_Inst1_n401), 
        .A2(DataPath_Registers_Inst1_n466), .B1(DataPath_Registers_Inst1_n462), 
        .B2(DataPath_Registers_Inst1_S3_6_), .C1(DataPath_Registers_Inst1_n353), .C2(DataPath_Registers_Inst1_S11_6_), .ZN(DataPath_Registers_Inst1_n509) );
  XOR2_X1 DataPath_Registers_Inst1_U93 ( .A(DataPath_Registers_Inst1_in4_5_), 
        .B(DataPath_Registers_Inst1_n400), .Z(DataPath_Registers_Inst1_n401)
         );
  XOR2_X1 DataPath_Registers_Inst1_U92 ( .A(DataPath_Registers_Inst1_in3_5_), 
        .B(DataPath_Registers_Inst1_in3_6_), .Z(DataPath_Registers_Inst1_n400)
         );
  INV_X1 DataPath_Registers_Inst1_U91 ( .A(DataPath_Registers_Inst1_n399), 
        .ZN(DataPath_Registers_Inst1_n275) );
  OAI22_X1 DataPath_Registers_Inst1_U90 ( .A1(DataPath_Registers_Inst1_n364), 
        .A2(DataPath_Registers_Inst1_n524), .B1(DataPath_Registers_Inst1_n206), 
        .B2(DataPath_Registers_Inst1_n360), .ZN(DataPath_Registers_Inst1_n399)
         );
  OAI222_X1 DataPath_Registers_Inst1_U89 ( .A1(DataPath_Registers_Inst1_n398), 
        .A2(DataPath_Registers_Inst1_n474), .B1(DataPath_Registers_Inst1_n480), 
        .B2(DataPath_Registers_Inst1_n219), .C1(DataPath_Registers_Inst1_n354), 
        .C2(DataPath_Registers_Inst1_n397), .ZN(DataPath_Registers_Inst1_n524)
         );
  INV_X1 DataPath_Registers_Inst1_U88 ( .A(DataPath_Registers_Inst1_S6_6_), 
        .ZN(DataPath_Registers_Inst1_n397) );
  XOR2_X1 DataPath_Registers_Inst1_U87 ( .A(DataPath_Registers_Inst1_n468), 
        .B(DataPath_Registers_Inst1_n396), .Z(DataPath_Registers_Inst1_n398)
         );
  XOR2_X1 DataPath_Registers_Inst1_U86 ( .A(DataPath_Registers_Inst1_in3_5_), 
        .B(DataPath_Registers_Inst1_in2_5_), .Z(DataPath_Registers_Inst1_n396)
         );
  INV_X1 DataPath_Registers_Inst1_U85 ( .A(DataPath_Registers_Inst1_in2_6_), 
        .ZN(DataPath_Registers_Inst1_n468) );
  AOI22_X1 DataPath_Registers_Inst1_U84 ( .A1(DataPath_Registers_Inst1_n356), 
        .A2(DataPath_Registers_Inst1_n493), .B1(DataPath_Registers_Inst1_n341), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n274)
         );
  AOI22_X1 DataPath_Registers_Inst1_U83 ( .A1(DataPath_Registers_Inst1_n466), 
        .A2(DataPath_Registers_Inst1_n395), .B1(DataPath_Registers_Inst1_n206), 
        .B2(DataPath_Registers_Inst1_n474), .ZN(DataPath_Registers_Inst1_n493)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U82 ( .A(DataPath_Registers_Inst1_n394), 
        .B(DataPath_Registers_Inst1_in1_6_), .ZN(DataPath_Registers_Inst1_n395) );
  XNOR2_X1 DataPath_Registers_Inst1_U81 ( .A(DataPath_Registers_Inst1_in1_5_), 
        .B(DataPath_Registers_Inst1_in2_5_), .ZN(DataPath_Registers_Inst1_n394) );
  MUX2_X1 DataPath_Registers_Inst1_U80 ( .A(DataPath_Registers_Inst1_S4_in[7]), 
        .B(DataPath_Registers_Inst1_S4_7_), .S(DataPath_Registers_Inst1_n366), 
        .Z(DataPath_Registers_Inst1_n273) );
  AOI22_X1 DataPath_Registers_Inst1_U79 ( .A1(DataPath_Registers_Inst1_n356), 
        .A2(DataPath_Registers_Inst1_n496), .B1(DataPath_Registers_Inst1_n215), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n272)
         );
  AOI22_X1 DataPath_Registers_Inst1_U78 ( .A1(DataPath_Registers_Inst1_n351), 
        .A2(StateIn1[7]), .B1(DataPath_Registers_Inst1_S4_7_), .B2(
        DataPath_Registers_Inst1_n354), .ZN(DataPath_Registers_Inst1_n496) );
  AOI22_X1 DataPath_Registers_Inst1_U77 ( .A1(DataPath_Registers_Inst1_n356), 
        .A2(DataPath_Registers_Inst1_n511), .B1(DataPath_Registers_Inst1_n266), 
        .B2(DataPath_Registers_Inst1_n364), .ZN(DataPath_Registers_Inst1_n271)
         );
  AOI222_X1 DataPath_Registers_Inst1_U76 ( .A1(DataPath_Registers_Inst1_n393), 
        .A2(DataPath_Registers_Inst1_n466), .B1(DataPath_Registers_Inst1_n462), 
        .B2(DataPath_Registers_Inst1_S3_7_), .C1(DataPath_Registers_Inst1_n353), .C2(DataPath_Registers_Inst1_S11_7_), .ZN(DataPath_Registers_Inst1_n511) );
  XOR2_X1 DataPath_Registers_Inst1_U75 ( .A(DataPath_Registers_Inst1_in3_6_), 
        .B(DataPath_Registers_Inst1_n392), .Z(DataPath_Registers_Inst1_n393)
         );
  AOI22_X1 DataPath_Registers_Inst1_U74 ( .A1(DataPath_Registers_Inst1_in3_7_), 
        .A2(DataPath_Registers_Inst1_in4_6_), .B1(
        DataPath_Registers_Inst1_n391), .B2(DataPath_Registers_Inst1_n476), 
        .ZN(DataPath_Registers_Inst1_n392) );
  AOI22_X1 DataPath_Registers_Inst1_U73 ( .A1(DataPath_Registers_Inst1_n356), 
        .A2(DataPath_Registers_Inst1_n520), .B1(DataPath_Registers_Inst1_n348), 
        .B2(DataPath_Registers_Inst1_n365), .ZN(DataPath_Registers_Inst1_n270)
         );
  AOI222_X1 DataPath_Registers_Inst1_U72 ( .A1(DataPath_Registers_Inst1_S2_4_), 
        .A2(DataPath_Registers_Inst1_n462), .B1(DataPath_Registers_Inst1_n466), 
        .B2(DataPath_Registers_Inst1_n390), .C1(DataPath_Registers_Inst1_n353), 
        .C2(DataPath_Registers_Inst1_S6_4_), .ZN(DataPath_Registers_Inst1_n520) );
  XNOR2_X1 DataPath_Registers_Inst1_U71 ( .A(DataPath_Registers_Inst1_n389), 
        .B(DataPath_Registers_Inst1_in2_4_), .ZN(DataPath_Registers_Inst1_n390) );
  XNOR2_X1 DataPath_Registers_Inst1_U70 ( .A(DataPath_Registers_Inst1_n458), 
        .B(DataPath_Registers_Inst1_n388), .ZN(DataPath_Registers_Inst1_n389)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U69 ( .A(DataPath_Registers_Inst1_n476), 
        .B(DataPath_Registers_Inst1_in3_3_), .ZN(DataPath_Registers_Inst1_n458) );
  INV_X1 DataPath_Registers_Inst1_U68 ( .A(DataPath_Registers_Inst1_in3_7_), 
        .ZN(DataPath_Registers_Inst1_n476) );
  NAND2_X1 DataPath_Registers_Inst1_U67 ( .A1(DataPath_Registers_Inst1_n354), 
        .A2(DataPath_Registers_Inst1_n387), .ZN(DataPath_Registers_Inst1_n480)
         );
  AOI22_X1 DataPath_Registers_Inst1_U66 ( .A1(DataPath_Registers_Inst1_n355), 
        .A2(DataPath_Registers_Inst1_n489), .B1(DataPath_Registers_Inst1_n340), 
        .B2(DataPath_Registers_Inst1_n364), .ZN(DataPath_Registers_Inst1_n269)
         );
  AOI22_X1 DataPath_Registers_Inst1_U65 ( .A1(DataPath_Registers_Inst1_n466), 
        .A2(DataPath_Registers_Inst1_n386), .B1(DataPath_Registers_Inst1_n204), 
        .B2(DataPath_Registers_Inst1_n474), .ZN(DataPath_Registers_Inst1_n489)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U64 ( .A(DataPath_Registers_Inst1_n385), 
        .B(DataPath_Registers_Inst1_in1_4_), .ZN(DataPath_Registers_Inst1_n386) );
  XNOR2_X1 DataPath_Registers_Inst1_U63 ( .A(DataPath_Registers_Inst1_n411), 
        .B(DataPath_Registers_Inst1_n388), .ZN(DataPath_Registers_Inst1_n385)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U62 ( .A(DataPath_Registers_Inst1_n467), 
        .B(DataPath_Registers_Inst1_in2_3_), .ZN(DataPath_Registers_Inst1_n388) );
  INV_X1 DataPath_Registers_Inst1_U61 ( .A(DataPath_Registers_Inst1_in2_7_), 
        .ZN(DataPath_Registers_Inst1_n467) );
  AOI22_X1 DataPath_Registers_Inst1_U60 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst1_n384), .B1(DataPath_Registers_Inst1_n347), 
        .B2(DataPath_Registers_Inst1_n387), .ZN(S0_output1[7]) );
  XNOR2_X1 DataPath_Registers_Inst1_U59 ( .A(DataPath_Registers_Inst1_in1_6_), 
        .B(DataPath_Registers_Inst1_n383), .ZN(DataPath_Registers_Inst1_n384)
         );
  AOI22_X1 DataPath_Registers_Inst1_U58 ( .A1(DataPath_Registers_Inst1_in4_7_), 
        .A2(DataPath_Registers_Inst1_in4_6_), .B1(
        DataPath_Registers_Inst1_n391), .B2(DataPath_Registers_Inst1_n441), 
        .ZN(DataPath_Registers_Inst1_n383) );
  AOI22_X1 DataPath_Registers_Inst1_U57 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst1_n382), .B1(DataPath_Registers_Inst1_n341), 
        .B2(DataPath_Registers_Inst1_n387), .ZN(S0_output1[6]) );
  XNOR2_X1 DataPath_Registers_Inst1_U56 ( .A(DataPath_Registers_Inst1_in1_5_), 
        .B(DataPath_Registers_Inst1_n381), .ZN(DataPath_Registers_Inst1_n382)
         );
  AOI22_X1 DataPath_Registers_Inst1_U55 ( .A1(DataPath_Registers_Inst1_in4_5_), 
        .A2(DataPath_Registers_Inst1_in4_6_), .B1(
        DataPath_Registers_Inst1_n391), .B2(DataPath_Registers_Inst1_n380), 
        .ZN(DataPath_Registers_Inst1_n381) );
  INV_X1 DataPath_Registers_Inst1_U54 ( .A(DataPath_Registers_Inst1_in4_6_), 
        .ZN(DataPath_Registers_Inst1_n391) );
  AOI22_X1 DataPath_Registers_Inst1_U53 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst1_n379), .B1(DataPath_Registers_Inst1_n342), 
        .B2(DataPath_Registers_Inst1_n387), .ZN(S0_output1[5]) );
  XOR2_X1 DataPath_Registers_Inst1_U52 ( .A(DataPath_Registers_Inst1_n380), 
        .B(DataPath_Registers_Inst1_n378), .Z(DataPath_Registers_Inst1_n379)
         );
  XOR2_X1 DataPath_Registers_Inst1_U51 ( .A(DataPath_Registers_Inst1_in1_4_), 
        .B(DataPath_Registers_Inst1_in4_4_), .Z(DataPath_Registers_Inst1_n378)
         );
  INV_X1 DataPath_Registers_Inst1_U50 ( .A(DataPath_Registers_Inst1_in4_5_), 
        .ZN(DataPath_Registers_Inst1_n380) );
  AOI22_X1 DataPath_Registers_Inst1_U49 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst1_n377), .B1(DataPath_Registers_Inst1_n340), 
        .B2(DataPath_Registers_Inst1_n387), .ZN(S0_output1[4]) );
  XNOR2_X1 DataPath_Registers_Inst1_U48 ( .A(DataPath_Registers_Inst1_in4_4_), 
        .B(DataPath_Registers_Inst1_n376), .ZN(DataPath_Registers_Inst1_n377)
         );
  XOR2_X1 DataPath_Registers_Inst1_U47 ( .A(DataPath_Registers_Inst1_n411), 
        .B(DataPath_Registers_Inst1_n459), .Z(DataPath_Registers_Inst1_n376)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U46 ( .A(DataPath_Registers_Inst1_n441), 
        .B(DataPath_Registers_Inst1_in4_3_), .ZN(DataPath_Registers_Inst1_n459) );
  XNOR2_X1 DataPath_Registers_Inst1_U45 ( .A(DataPath_Registers_Inst1_n463), 
        .B(DataPath_Registers_Inst1_in1_3_), .ZN(DataPath_Registers_Inst1_n411) );
  AOI22_X1 DataPath_Registers_Inst1_U44 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst1_n375), .B1(DataPath_Registers_Inst1_n343), 
        .B2(DataPath_Registers_Inst1_n387), .ZN(S0_output1[3]) );
  XOR2_X1 DataPath_Registers_Inst1_U43 ( .A(DataPath_Registers_Inst1_n463), 
        .B(DataPath_Registers_Inst1_n374), .Z(DataPath_Registers_Inst1_n375)
         );
  XNOR2_X1 DataPath_Registers_Inst1_U42 ( .A(DataPath_Registers_Inst1_n373), 
        .B(DataPath_Registers_Inst1_in4_3_), .ZN(DataPath_Registers_Inst1_n374) );
  XNOR2_X1 DataPath_Registers_Inst1_U41 ( .A(DataPath_Registers_Inst1_n418), 
        .B(DataPath_Registers_Inst1_in1_2_), .ZN(DataPath_Registers_Inst1_n373) );
  XNOR2_X1 DataPath_Registers_Inst1_U40 ( .A(DataPath_Registers_Inst1_n441), 
        .B(DataPath_Registers_Inst1_in4_2_), .ZN(DataPath_Registers_Inst1_n418) );
  AOI22_X1 DataPath_Registers_Inst1_U39 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst1_n372), .B1(DataPath_Registers_Inst1_n344), 
        .B2(DataPath_Registers_Inst1_n387), .ZN(S0_output1[2]) );
  XNOR2_X1 DataPath_Registers_Inst1_U38 ( .A(DataPath_Registers_Inst1_in4_1_), 
        .B(DataPath_Registers_Inst1_n371), .ZN(DataPath_Registers_Inst1_n372)
         );
  XOR2_X1 DataPath_Registers_Inst1_U37 ( .A(DataPath_Registers_Inst1_in1_1_), 
        .B(DataPath_Registers_Inst1_in4_2_), .Z(DataPath_Registers_Inst1_n371)
         );
  AOI22_X1 DataPath_Registers_Inst1_U36 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst1_n370), .B1(DataPath_Registers_Inst1_n345), 
        .B2(DataPath_Registers_Inst1_n387), .ZN(S0_output1[1]) );
  XNOR2_X1 DataPath_Registers_Inst1_U35 ( .A(DataPath_Registers_Inst1_in4_1_), 
        .B(DataPath_Registers_Inst1_n369), .ZN(DataPath_Registers_Inst1_n370)
         );
  AOI22_X1 DataPath_Registers_Inst1_U34 ( .A1(DataPath_Registers_Inst1_n368), 
        .A2(DataPath_Registers_Inst1_n439), .B1(DataPath_Registers_Inst1_n438), 
        .B2(DataPath_Registers_Inst1_n434), .ZN(DataPath_Registers_Inst1_n369)
         );
  INV_X1 DataPath_Registers_Inst1_U33 ( .A(DataPath_Registers_Inst1_n438), 
        .ZN(DataPath_Registers_Inst1_n439) );
  XOR2_X1 DataPath_Registers_Inst1_U32 ( .A(DataPath_Registers_Inst1_n463), 
        .B(DataPath_Registers_Inst1_in1_0_), .Z(DataPath_Registers_Inst1_n438)
         );
  AOI22_X1 DataPath_Registers_Inst1_U31 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst1_n367), .B1(DataPath_Registers_Inst1_n346), 
        .B2(DataPath_Registers_Inst1_n387), .ZN(S0_output1[0]) );
  INV_X1 DataPath_Registers_Inst1_U30 ( .A(DoMC), .ZN(
        DataPath_Registers_Inst1_n387) );
  AOI22_X1 DataPath_Registers_Inst1_U29 ( .A1(DataPath_Registers_Inst1_n368), 
        .A2(DataPath_Registers_Inst1_n463), .B1(
        DataPath_Registers_Inst1_in1_7_), .B2(DataPath_Registers_Inst1_n434), 
        .ZN(DataPath_Registers_Inst1_n367) );
  INV_X1 DataPath_Registers_Inst1_U28 ( .A(DataPath_Registers_Inst1_in1_7_), 
        .ZN(DataPath_Registers_Inst1_n463) );
  INV_X1 DataPath_Registers_Inst1_U27 ( .A(DataPath_Registers_Inst1_n434), 
        .ZN(DataPath_Registers_Inst1_n368) );
  XOR2_X1 DataPath_Registers_Inst1_U26 ( .A(DataPath_Registers_Inst1_n441), 
        .B(DataPath_Registers_Inst1_in4_0_), .Z(DataPath_Registers_Inst1_n434)
         );
  INV_X1 DataPath_Registers_Inst1_U25 ( .A(DataPath_Registers_Inst1_in4_7_), 
        .ZN(DataPath_Registers_Inst1_n441) );
  INV_X2 DataPath_Registers_Inst1_U24 ( .A(DataPath_Registers_Inst1_n354), 
        .ZN(DataPath_Registers_Inst1_n353) );
  INV_X1 DataPath_Registers_Inst1_U23 ( .A(DataPath_Registers_Inst1_n480), 
        .ZN(DataPath_Registers_Inst1_n462) );
  NAND2_X1 DataPath_Registers_Inst1_U22 ( .A1(DataPath_Registers_Inst1_n354), 
        .A2(DoMC), .ZN(DataPath_Registers_Inst1_n474) );
  INV_X1 DataPath_Registers_Inst1_U21 ( .A(DataPath_Registers_Inst1_n474), 
        .ZN(DataPath_Registers_Inst1_n466) );
  INV_X2 DataPath_Registers_Inst1_U20 ( .A(DataPath_Registers_Inst1_n354), 
        .ZN(DataPath_Registers_Inst1_n351) );
  INV_X2 DataPath_Registers_Inst1_U19 ( .A(DataPath_Registers_Inst1_n354), 
        .ZN(DataPath_Registers_Inst1_n352) );
  INV_X1 DataPath_Registers_Inst1_U18 ( .A(DataPath_Registers_Inst1_n366), 
        .ZN(DataPath_Registers_Inst1_n358) );
  INV_X1 DataPath_Registers_Inst1_U17 ( .A(DataPath_Registers_Inst1_n366), 
        .ZN(DataPath_Registers_Inst1_n356) );
  INV_X1 DataPath_Registers_Inst1_U16 ( .A(DataPath_Registers_Inst1_n366), 
        .ZN(DataPath_Registers_Inst1_n359) );
  INV_X1 DataPath_Registers_Inst1_U15 ( .A(DataPath_Registers_Inst1_n366), 
        .ZN(DataPath_Registers_Inst1_n357) );
  INV_X1 DataPath_Registers_Inst1_U14 ( .A(DataPath_Registers_Inst1_n366), 
        .ZN(DataPath_Registers_Inst1_n361) );
  INV_X1 DataPath_Registers_Inst1_U13 ( .A(DataPath_Registers_Inst1_n366), 
        .ZN(DataPath_Registers_Inst1_n360) );
  INV_X2 DataPath_Registers_Inst1_U12 ( .A(DataPath_Registers_Inst1_n366), 
        .ZN(DataPath_Registers_Inst1_n363) );
  INV_X1 DataPath_Registers_Inst1_U11 ( .A(DataPath_Registers_Inst1_n366), 
        .ZN(DataPath_Registers_Inst1_n362) );
  INV_X1 DataPath_Registers_Inst1_U10 ( .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst1_n365) );
  BUF_X1 DataPath_Registers_Inst1_U9 ( .A(DataPath_Registers_Inst1_n365), .Z(
        DataPath_Registers_Inst1_n364) );
  INV_X1 DataPath_Registers_Inst1_U8 ( .A(DataPath_Registers_Inst1_n364), .ZN(
        DataPath_Registers_Inst1_n355) );
  INV_X1 DataPath_Registers_Inst1_U7 ( .A(DoSR), .ZN(
        DataPath_Registers_Inst1_n354) );
  INV_X1 DataPath_Registers_Inst1_U6 ( .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst1_n366) );
  AOI211_X1 DataPath_Registers_Inst1_U5 ( .C1(DataPath_Registers_Inst1_S11_0_), 
        .C2(DataPath_Registers_Inst1_n353), .A(DataPath_Registers_Inst1_n337), 
        .B(DataPath_Registers_Inst1_n339), .ZN(DataPath_Registers_Inst1_n497)
         );
  AOI221_X1 DataPath_Registers_Inst1_U4 ( .B1(DataPath_Registers_Inst1_in4_7_), 
        .B2(DataPath_Registers_Inst1_n338), .C1(DataPath_Registers_Inst1_n441), 
        .C2(DataPath_Registers_Inst1_n442), .A(DataPath_Registers_Inst1_n474), 
        .ZN(DataPath_Registers_Inst1_n339) );
  INV_X1 DataPath_Registers_Inst1_U3 ( .A(DataPath_Registers_Inst1_n442), .ZN(
        DataPath_Registers_Inst1_n338) );
  NOR2_X1 DataPath_Registers_Inst1_U2 ( .A1(DataPath_Registers_Inst1_n480), 
        .A2(DataPath_Registers_Inst1_n246), .ZN(DataPath_Registers_Inst1_n337)
         );
  DFF_X1 DataPath_Registers_Inst1_S3_reg_3_ ( .D(DataPath_Registers_Inst1_n289), .CK(clk), .Q(DataPath_Registers_Inst1_S3_3_), .QN(
        DataPath_Registers_Inst1_n231) );
  DFF_X1 DataPath_Registers_Inst1_S12_reg_0_ ( .D(
        DataPath_Registers_Inst1_n320), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_0_), .QN(DataPath_Registers_Inst1_n262)
         );
  DFF_X1 DataPath_Registers_Inst1_S12_reg_1_ ( .D(
        DataPath_Registers_Inst1_n319), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_1_), .QN(DataPath_Registers_Inst1_n261)
         );
  DFF_X1 DataPath_Registers_Inst1_S12_reg_2_ ( .D(
        DataPath_Registers_Inst1_n318), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_2_), .QN(DataPath_Registers_Inst1_n260)
         );
  DFF_X1 DataPath_Registers_Inst1_S12_reg_3_ ( .D(
        DataPath_Registers_Inst1_n317), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_3_), .QN(DataPath_Registers_Inst1_n259)
         );
  DFF_X1 DataPath_Registers_Inst1_S12_reg_4_ ( .D(
        DataPath_Registers_Inst1_n316), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_4_), .QN(DataPath_Registers_Inst1_n258)
         );
  DFF_X1 DataPath_Registers_Inst1_S12_reg_5_ ( .D(
        DataPath_Registers_Inst1_n315), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_5_), .QN(DataPath_Registers_Inst1_n257)
         );
  DFF_X1 DataPath_Registers_Inst1_S12_reg_7_ ( .D(
        DataPath_Registers_Inst1_n313), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_7_), .QN(DataPath_Registers_Inst1_n255)
         );
  DFF_X1 DataPath_Registers_Inst1_S8_reg_1_ ( .D(DataPath_Registers_Inst1_n312), .CK(clk), .Q(DataPath_Registers_Inst1_S8_1_), .QN(
        DataPath_Registers_Inst1_n254) );
  DFF_X1 DataPath_Registers_Inst1_S8_reg_2_ ( .D(DataPath_Registers_Inst1_n311), .CK(clk), .Q(DataPath_Registers_Inst1_S8_2_), .QN(
        DataPath_Registers_Inst1_n253) );
  DFF_X1 DataPath_Registers_Inst1_S8_reg_3_ ( .D(DataPath_Registers_Inst1_n310), .CK(clk), .Q(DataPath_Registers_Inst1_S8_3_), .QN(
        DataPath_Registers_Inst1_n252) );
  DFF_X1 DataPath_Registers_Inst1_S8_reg_4_ ( .D(DataPath_Registers_Inst1_n309), .CK(clk), .Q(DataPath_Registers_Inst1_S8_4_), .QN(
        DataPath_Registers_Inst1_n251) );
  DFF_X1 DataPath_Registers_Inst1_S8_reg_6_ ( .D(DataPath_Registers_Inst1_n307), .CK(clk), .Q(DataPath_Registers_Inst1_S8_6_), .QN(
        DataPath_Registers_Inst1_n249) );
  DFF_X1 DataPath_Registers_Inst1_S12_reg_6_ ( .D(
        DataPath_Registers_Inst1_n314), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_6_), .QN(DataPath_Registers_Inst1_n256)
         );
  DFF_X1 DataPath_Registers_Inst1_S0_reg_6_ ( .D(DataPath_Registers_Inst1_n274), .CK(clk), .Q(), .QN(DataPath_Registers_Inst1_n341) );
  DFF_X1 DataPath_Registers_Inst1_S0_reg_4_ ( .D(DataPath_Registers_Inst1_n269), .CK(clk), .Q(), .QN(DataPath_Registers_Inst1_n340) );
  DFF_X1 DataPath_Registers_Inst1_S1_reg_4_ ( .D(DataPath_Registers_Inst1_n270), .CK(clk), .Q(DataPath_Registers_Inst1_n204), .QN(
        DataPath_Registers_Inst1_n348) );
  DFF_X1 DataPath_Registers_Inst1_S2_reg_7_ ( .D(DataPath_Registers_Inst1_n271), .CK(clk), .Q(DataPath_Registers_Inst1_S2_7_), .QN(
        DataPath_Registers_Inst1_n266) );
  DFF_X1 DataPath_Registers_Inst1_S3_reg_7_ ( .D(DataPath_Registers_Inst1_n272), .CK(clk), .Q(DataPath_Registers_Inst1_S3_7_), .QN(
        DataPath_Registers_Inst1_n215) );
  DFF_X1 DataPath_Registers_Inst1_S4_reg_7_ ( .D(DataPath_Registers_Inst1_n273), .CK(clk), .Q(DataPath_Registers_Inst1_S4_7_), .QN() );
  DFF_X1 DataPath_Registers_Inst1_S1_reg_6_ ( .D(DataPath_Registers_Inst1_n275), .CK(clk), .Q(DataPath_Registers_Inst1_n206), .QN() );
  DFF_X1 DataPath_Registers_Inst1_S2_reg_6_ ( .D(DataPath_Registers_Inst1_n276), .CK(clk), .Q(DataPath_Registers_Inst1_S2_6_), .QN(
        DataPath_Registers_Inst1_n219) );
  DFF_X1 DataPath_Registers_Inst1_S3_reg_6_ ( .D(DataPath_Registers_Inst1_n277), .CK(clk), .Q(DataPath_Registers_Inst1_S3_6_), .QN(
        DataPath_Registers_Inst1_n220) );
  DFF_X1 DataPath_Registers_Inst1_S4_reg_6_ ( .D(DataPath_Registers_Inst1_n278), .CK(clk), .Q(DataPath_Registers_Inst1_S4_6_), .QN() );
  DFF_X1 DataPath_Registers_Inst1_S0_reg_5_ ( .D(DataPath_Registers_Inst1_n279), .CK(clk), .Q(), .QN(DataPath_Registers_Inst1_n342) );
  DFF_X1 DataPath_Registers_Inst1_S1_reg_5_ ( .D(DataPath_Registers_Inst1_n280), .CK(clk), .Q(DataPath_Registers_Inst1_n208), .QN() );
  DFF_X1 DataPath_Registers_Inst1_S2_reg_5_ ( .D(DataPath_Registers_Inst1_n281), .CK(clk), .Q(DataPath_Registers_Inst1_S2_5_), .QN(
        DataPath_Registers_Inst1_n224) );
  DFF_X1 DataPath_Registers_Inst1_S3_reg_5_ ( .D(DataPath_Registers_Inst1_n282), .CK(clk), .Q(DataPath_Registers_Inst1_S3_5_), .QN(
        DataPath_Registers_Inst1_n225) );
  DFF_X1 DataPath_Registers_Inst1_S4_reg_5_ ( .D(DataPath_Registers_Inst1_n283), .CK(clk), .Q(DataPath_Registers_Inst1_S4_5_), .QN() );
  DFF_X1 DataPath_Registers_Inst1_S3_reg_4_ ( .D(DataPath_Registers_Inst1_n284), .CK(clk), .Q(DataPath_Registers_Inst1_S3_4_), .QN(
        DataPath_Registers_Inst1_n263) );
  DFF_X1 DataPath_Registers_Inst1_S4_reg_4_ ( .D(DataPath_Registers_Inst1_n285), .CK(clk), .Q(DataPath_Registers_Inst1_S4_4_), .QN(
        DataPath_Registers_Inst1_n227) );
  DFF_X1 DataPath_Registers_Inst1_S0_reg_3_ ( .D(DataPath_Registers_Inst1_n286), .CK(clk), .Q(), .QN(DataPath_Registers_Inst1_n343) );
  DFF_X1 DataPath_Registers_Inst1_S1_reg_3_ ( .D(DataPath_Registers_Inst1_n287), .CK(clk), .Q(DataPath_Registers_Inst1_n210), .QN(
        DataPath_Registers_Inst1_n349) );
  DFF_X1 DataPath_Registers_Inst1_S2_reg_3_ ( .D(DataPath_Registers_Inst1_n288), .CK(clk), .Q(DataPath_Registers_Inst1_S2_3_), .QN(
        DataPath_Registers_Inst1_n230) );
  DFF_X1 DataPath_Registers_Inst1_S4_reg_3_ ( .D(DataPath_Registers_Inst1_n290), .CK(clk), .Q(DataPath_Registers_Inst1_S4_3_), .QN(
        DataPath_Registers_Inst1_n232) );
  DFF_X1 DataPath_Registers_Inst1_S0_reg_2_ ( .D(DataPath_Registers_Inst1_n291), .CK(clk), .Q(), .QN(DataPath_Registers_Inst1_n344) );
  DFF_X1 DataPath_Registers_Inst1_S1_reg_2_ ( .D(DataPath_Registers_Inst1_n292), .CK(clk), .Q(DataPath_Registers_Inst1_n212), .QN() );
  DFF_X1 DataPath_Registers_Inst1_S2_reg_2_ ( .D(DataPath_Registers_Inst1_n293), .CK(clk), .Q(DataPath_Registers_Inst1_S2_2_), .QN(
        DataPath_Registers_Inst1_n235) );
  DFF_X1 DataPath_Registers_Inst1_S3_reg_2_ ( .D(DataPath_Registers_Inst1_n294), .CK(clk), .Q(DataPath_Registers_Inst1_S3_2_), .QN(
        DataPath_Registers_Inst1_n236) );
  DFF_X1 DataPath_Registers_Inst1_S4_reg_2_ ( .D(DataPath_Registers_Inst1_n295), .CK(clk), .Q(DataPath_Registers_Inst1_S4_2_), .QN() );
  DFF_X1 DataPath_Registers_Inst1_S0_reg_1_ ( .D(DataPath_Registers_Inst1_n296), .CK(clk), .Q(), .QN(DataPath_Registers_Inst1_n345) );
  DFF_X1 DataPath_Registers_Inst1_S1_reg_1_ ( .D(DataPath_Registers_Inst1_n297), .CK(clk), .Q(DataPath_Registers_Inst1_n202), .QN(
        DataPath_Registers_Inst1_n350) );
  DFF_X1 DataPath_Registers_Inst1_S2_reg_1_ ( .D(DataPath_Registers_Inst1_n298), .CK(clk), .Q(DataPath_Registers_Inst1_S2_1_), .QN(
        DataPath_Registers_Inst1_n240) );
  DFF_X1 DataPath_Registers_Inst1_S3_reg_1_ ( .D(DataPath_Registers_Inst1_n299), .CK(clk), .Q(DataPath_Registers_Inst1_S3_1_), .QN(
        DataPath_Registers_Inst1_n241) );
  DFF_X1 DataPath_Registers_Inst1_S4_reg_1_ ( .D(DataPath_Registers_Inst1_n300), .CK(clk), .Q(DataPath_Registers_Inst1_S4_1_), .QN(
        DataPath_Registers_Inst1_n242) );
  DFF_X1 DataPath_Registers_Inst1_S0_reg_0_ ( .D(DataPath_Registers_Inst1_n301), .CK(clk), .Q(), .QN(DataPath_Registers_Inst1_n346) );
  DFF_X1 DataPath_Registers_Inst1_S1_reg_0_ ( .D(DataPath_Registers_Inst1_n6), 
        .CK(clk), .Q(DataPath_Registers_Inst1_n201), .QN() );
  DFF_X1 DataPath_Registers_Inst1_S2_reg_0_ ( .D(DataPath_Registers_Inst1_n303), .CK(clk), .Q(DataPath_Registers_Inst1_S2_0_), .QN(
        DataPath_Registers_Inst1_n245) );
  DFF_X1 DataPath_Registers_Inst1_S3_reg_0_ ( .D(DataPath_Registers_Inst1_n304), .CK(clk), .Q(DataPath_Registers_Inst1_S3_0_), .QN(
        DataPath_Registers_Inst1_n246) );
  DFF_X1 DataPath_Registers_Inst1_S4_reg_0_ ( .D(DataPath_Registers_Inst1_n305), .CK(clk), .Q(DataPath_Registers_Inst1_S4_0_), .QN() );
  DFF_X1 DataPath_Registers_Inst1_S8_reg_7_ ( .D(DataPath_Registers_Inst1_n306), .CK(clk), .Q(DataPath_Registers_Inst1_S8_7_), .QN(
        DataPath_Registers_Inst1_n248) );
  DFF_X1 DataPath_Registers_Inst1_S8_reg_5_ ( .D(DataPath_Registers_Inst1_n308), .CK(clk), .Q(DataPath_Registers_Inst1_S8_5_), .QN(
        DataPath_Registers_Inst1_n250) );
  DFF_X1 DataPath_Registers_Inst1_S2_reg_4_ ( .D(DataPath_Registers_Inst1_n321), .CK(clk), .Q(DataPath_Registers_Inst1_S2_4_), .QN(
        DataPath_Registers_Inst1_n264) );
  DFF_X1 DataPath_Registers_Inst1_S0_reg_7_ ( .D(DataPath_Registers_Inst1_n322), .CK(clk), .Q(), .QN(DataPath_Registers_Inst1_n347) );
  DFF_X1 DataPath_Registers_Inst1_S1_reg_7_ ( .D(DataPath_Registers_Inst1_n323), .CK(clk), .Q(DataPath_Registers_Inst1_n203), .QN() );
  DFF_X1 DataPath_Registers_Inst1_S8_reg_0_ ( .D(DataPath_Registers_Inst1_n324), .CK(clk), .Q(DataPath_Registers_Inst1_S8_0_), .QN(
        DataPath_Registers_Inst1_n268) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst1_n359), .B2(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_0_U3 ( .B1(
        DataPath_Registers_Inst1_n353), .B2(DataPath_Registers_Inst1_S6_0_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n9), .C2(
        DataPath_Registers_Inst1_S10_0_), .A(DataPath_Registers_Inst1_n359), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_0_U2 ( .A(
        DataPath_Registers_Inst1_n353), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S4_in[0]), .QN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_0_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst1_n359), .B2(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_1_U3 ( .B1(
        DataPath_Registers_Inst1_n353), .B2(DataPath_Registers_Inst1_S6_1_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n10), .C2(
        DataPath_Registers_Inst1_S10_1_), .A(DataPath_Registers_Inst1_n359), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_1_U2 ( .A(
        DataPath_Registers_Inst1_n353), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S4_in[1]), .QN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst1_n359), .B2(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_2_U3 ( .B1(
        DataPath_Registers_Inst1_n353), .B2(DataPath_Registers_Inst1_S6_2_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n9), .C2(
        DataPath_Registers_Inst1_S10_2_), .A(DataPath_Registers_Inst1_n359), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_2_U2 ( .A(
        DataPath_Registers_Inst1_n353), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S4_in[2]), .QN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_2_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst1_n359), .B2(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_3_U3 ( .B1(
        DataPath_Registers_Inst1_n353), .B2(DataPath_Registers_Inst1_S6_3_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n9), .C2(
        DataPath_Registers_Inst1_S10_3_), .A(DataPath_Registers_Inst1_n359), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_3_U2 ( .A(
        DataPath_Registers_Inst1_n353), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S4_in[3]), .QN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_3_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst1_n359), .B2(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_4_U3 ( .B1(
        DataPath_Registers_Inst1_n353), .B2(DataPath_Registers_Inst1_S6_4_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n9), .C2(
        DataPath_Registers_Inst1_S10_4_), .A(DataPath_Registers_Inst1_n359), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_4_U2 ( .A(
        DataPath_Registers_Inst1_n353), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S4_in[4]), .QN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_4_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst1_n359), .B2(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_5_U3 ( .B1(
        DataPath_Registers_Inst1_n353), .B2(DataPath_Registers_Inst1_S6_5_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n9), .C2(
        DataPath_Registers_Inst1_S10_5_), .A(DataPath_Registers_Inst1_n359), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_5_U2 ( .A(
        DataPath_Registers_Inst1_n353), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S4_in[5]), .QN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_5_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst1_n359), .B2(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_6_U3 ( .B1(
        DataPath_Registers_Inst1_n353), .B2(DataPath_Registers_Inst1_S6_6_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n9), .C2(
        DataPath_Registers_Inst1_S10_6_), .A(DataPath_Registers_Inst1_n359), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_6_U2 ( .A(
        DataPath_Registers_Inst1_n353), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S4_in[6]), .QN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_6_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst1_n359), .B2(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_7_U3 ( .B1(
        DataPath_Registers_Inst1_n353), .B2(DataPath_Registers_Inst1_S6_7_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n9), .C2(
        DataPath_Registers_Inst1_S10_7_), .A(DataPath_Registers_Inst1_n359), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_7_U2 ( .A(
        DataPath_Registers_Inst1_n353), .ZN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S5_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S4_in[7]), .QN(
        DataPath_Registers_Inst1_ScanFF_S5_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_0_U5 ( .B1(
        DataPath_Registers_Inst1_n362), .B2(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n10), .B2(
        DataPath_Registers_Inst1_S7_0_), .C1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n11), .C2(
        DataPath_Registers_Inst1_S15_0_), .A(DataPath_Registers_Inst1_n362), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_0_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_0_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S6_0_), .QN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_1_U5 ( .B1(
        DataPath_Registers_Inst1_n362), .B2(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n10), .B2(
        DataPath_Registers_Inst1_S7_1_), .C1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n11), .C2(
        DataPath_Registers_Inst1_S15_1_), .A(DataPath_Registers_Inst1_n362), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_1_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_1_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S6_1_), .QN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_2_U5 ( .B1(
        DataPath_Registers_Inst1_n362), .B2(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n10), .B2(
        DataPath_Registers_Inst1_S7_2_), .C1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n11), .C2(
        DataPath_Registers_Inst1_S15_2_), .A(DataPath_Registers_Inst1_n362), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_2_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_2_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S6_2_), .QN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_3_U5 ( .B1(
        DataPath_Registers_Inst1_n362), .B2(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n10), .B2(
        DataPath_Registers_Inst1_S7_3_), .C1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n11), .C2(
        DataPath_Registers_Inst1_S15_3_), .A(DataPath_Registers_Inst1_n362), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_3_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_3_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S6_3_), .QN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_4_U5 ( .B1(
        DataPath_Registers_Inst1_n362), .B2(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n10), .B2(
        DataPath_Registers_Inst1_S7_4_), .C1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n11), .C2(
        DataPath_Registers_Inst1_S15_4_), .A(DataPath_Registers_Inst1_n362), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_4_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_4_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S6_4_), .QN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst1_n362), .B2(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n10), .B2(
        DataPath_Registers_Inst1_S7_5_), .C1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n11), .C2(
        DataPath_Registers_Inst1_S15_5_), .A(DataPath_Registers_Inst1_n362), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_5_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_5_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S6_5_), .QN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_5_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst1_n362), .B2(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n10), .B2(
        DataPath_Registers_Inst1_S7_6_), .C1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n11), .C2(
        DataPath_Registers_Inst1_S15_6_), .A(DataPath_Registers_Inst1_n362), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_6_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_6_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S6_6_), .QN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_6_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst1_n362), .B2(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n10), .B2(
        DataPath_Registers_Inst1_S7_7_), .C1(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n11), .C2(
        DataPath_Registers_Inst1_S15_7_), .A(DataPath_Registers_Inst1_n362), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_7_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_7_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S6_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S6_7_), .QN(
        DataPath_Registers_Inst1_ScanFF_S6_SFF_7_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_0_U5 ( .B1(
        DataPath_Registers_Inst1_n361), .B2(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n10), .B2(
        DataPath_Registers_Inst1_S8_0_), .C1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n11), .C2(
        DataPath_Registers_Inst1_S4_0_), .A(DataPath_Registers_Inst1_n361), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_0_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_0_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S7_0_), .QN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_1_U5 ( .B1(
        DataPath_Registers_Inst1_n361), .B2(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n10), .B2(
        DataPath_Registers_Inst1_S8_1_), .C1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n11), .C2(
        DataPath_Registers_Inst1_S4_1_), .A(DataPath_Registers_Inst1_n361), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_1_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_1_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S7_1_), .QN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_2_U5 ( .B1(
        DataPath_Registers_Inst1_n361), .B2(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n10), .B2(
        DataPath_Registers_Inst1_S8_2_), .C1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n11), .C2(
        DataPath_Registers_Inst1_S4_2_), .A(DataPath_Registers_Inst1_n361), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_2_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_2_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S7_2_), .QN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst1_n361), .B2(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_3_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(DataPath_Registers_Inst1_S8_3_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n10), .C2(
        DataPath_Registers_Inst1_S4_3_), .A(DataPath_Registers_Inst1_n361), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_3_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S7_3_), .QN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_4_U5 ( .B1(
        DataPath_Registers_Inst1_n361), .B2(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n9), .B2(
        DataPath_Registers_Inst1_S8_4_), .C1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n10), .C2(
        DataPath_Registers_Inst1_S4_4_), .A(DataPath_Registers_Inst1_n361), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_4_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_4_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S7_4_), .QN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_4_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst1_n361), .B2(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n9), .B2(
        DataPath_Registers_Inst1_S8_5_), .C1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n10), .C2(
        DataPath_Registers_Inst1_S4_5_), .A(DataPath_Registers_Inst1_n361), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_5_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_5_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S7_5_), .QN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_5_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst1_n361), .B2(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n9), .B2(
        DataPath_Registers_Inst1_S8_6_), .C1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n10), .C2(
        DataPath_Registers_Inst1_S4_6_), .A(DataPath_Registers_Inst1_n361), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_6_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_6_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S7_6_), .QN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_6_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst1_n361), .B2(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n9), .B2(
        DataPath_Registers_Inst1_S8_7_), .C1(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n10), .C2(
        DataPath_Registers_Inst1_S4_7_), .A(DataPath_Registers_Inst1_n361), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_7_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_7_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S7_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S7_7_), .QN(
        DataPath_Registers_Inst1_ScanFF_S7_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_0_U5 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n10), .B2(
        DataPath_Registers_Inst1_S10_0_), .C1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n11), .C2(
        DataPath_Registers_Inst1_S14_0_), .A(DataPath_Registers_Inst1_n355), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_0_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_0_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S8_in[0]), .QN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_1_U5 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n10), .B2(
        DataPath_Registers_Inst1_S10_1_), .C1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n11), .C2(
        DataPath_Registers_Inst1_S14_1_), .A(DataPath_Registers_Inst1_n355), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_1_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_1_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S8_in[1]), .QN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_2_U5 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n10), .B2(
        DataPath_Registers_Inst1_S10_2_), .C1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n11), .C2(
        DataPath_Registers_Inst1_S14_2_), .A(DataPath_Registers_Inst1_n355), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_2_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_2_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S8_in[2]), .QN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_3_U5 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n10), .B2(
        DataPath_Registers_Inst1_S10_3_), .C1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n11), .C2(
        DataPath_Registers_Inst1_S14_3_), .A(DataPath_Registers_Inst1_n355), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_3_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_3_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S8_in[3]), .QN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_4_U5 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n10), .B2(
        DataPath_Registers_Inst1_S10_4_), .C1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n11), .C2(
        DataPath_Registers_Inst1_S14_4_), .A(DataPath_Registers_Inst1_n355), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_4_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_4_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S8_in[4]), .QN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n10), .B2(
        DataPath_Registers_Inst1_S10_5_), .C1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n11), .C2(
        DataPath_Registers_Inst1_S14_5_), .A(DataPath_Registers_Inst1_n355), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_5_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_5_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S8_in[5]), .QN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_5_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n10), .B2(
        DataPath_Registers_Inst1_S10_6_), .C1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n11), .C2(
        DataPath_Registers_Inst1_S14_6_), .A(DataPath_Registers_Inst1_n355), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_6_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_6_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S8_in[6]), .QN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_6_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n10), .B2(
        DataPath_Registers_Inst1_S10_7_), .C1(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n11), .C2(
        DataPath_Registers_Inst1_S14_7_), .A(DataPath_Registers_Inst1_n355), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_7_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_7_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S9_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S8_in[7]), .QN(
        DataPath_Registers_Inst1_ScanFF_S9_SFF_7_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst1_n360), .B2(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_0_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(DataPath_Registers_Inst1_S11_0_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n10), .C2(
        DataPath_Registers_Inst1_S3_0_), .A(DataPath_Registers_Inst1_n360), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_0_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S10_0_), .QN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst1_n360), .B2(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_1_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(DataPath_Registers_Inst1_S11_1_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n10), .C2(
        DataPath_Registers_Inst1_S3_1_), .A(DataPath_Registers_Inst1_n360), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_1_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S10_1_), .QN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst1_n360), .B2(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_2_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(DataPath_Registers_Inst1_S11_2_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n10), .C2(
        DataPath_Registers_Inst1_S3_2_), .A(DataPath_Registers_Inst1_n360), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_2_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S10_2_), .QN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst1_n360), .B2(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_3_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(DataPath_Registers_Inst1_S11_3_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n10), .C2(
        DataPath_Registers_Inst1_S3_3_), .A(DataPath_Registers_Inst1_n360), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_3_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S10_3_), .QN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst1_n360), .B2(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_4_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(DataPath_Registers_Inst1_S11_4_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n10), .C2(
        DataPath_Registers_Inst1_S3_4_), .A(DataPath_Registers_Inst1_n360), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_4_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S10_4_), .QN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst1_n360), .B2(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n9), .B2(
        DataPath_Registers_Inst1_S11_5_), .C1(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n10), .C2(
        DataPath_Registers_Inst1_S3_5_), .A(DataPath_Registers_Inst1_n360), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_5_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_5_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S10_5_), .QN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_5_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst1_n360), .B2(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n9), .B2(
        DataPath_Registers_Inst1_S11_6_), .C1(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n10), .C2(
        DataPath_Registers_Inst1_S3_6_), .A(DataPath_Registers_Inst1_n360), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_6_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_6_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S10_6_), .QN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_6_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst1_n360), .B2(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n9), .B2(
        DataPath_Registers_Inst1_S11_7_), .C1(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n10), .C2(
        DataPath_Registers_Inst1_S3_7_), .A(DataPath_Registers_Inst1_n360), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_7_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_7_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S10_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S10_7_), .QN(
        DataPath_Registers_Inst1_ScanFF_S10_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_0_U5 ( .B1(
        DataPath_Registers_Inst1_n356), .B2(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n10), .B2(
        DataPath_Registers_Inst1_S12_0_), .C1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n11), .C2(
        DataPath_Registers_Inst1_S8_0_), .A(DataPath_Registers_Inst1_n356), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_0_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_0_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S11_0_), .QN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_1_U5 ( .B1(
        DataPath_Registers_Inst1_n356), .B2(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n10), .B2(
        DataPath_Registers_Inst1_S12_1_), .C1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n11), .C2(
        DataPath_Registers_Inst1_S8_1_), .A(DataPath_Registers_Inst1_n356), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_1_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_1_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S11_1_), .QN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_2_U5 ( .B1(
        DataPath_Registers_Inst1_n356), .B2(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n10), .B2(
        DataPath_Registers_Inst1_S12_2_), .C1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n11), .C2(
        DataPath_Registers_Inst1_S8_2_), .A(DataPath_Registers_Inst1_n356), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_2_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_2_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S11_2_), .QN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_3_U5 ( .B1(
        DataPath_Registers_Inst1_n356), .B2(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n10), .B2(
        DataPath_Registers_Inst1_S12_3_), .C1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n11), .C2(
        DataPath_Registers_Inst1_S8_3_), .A(DataPath_Registers_Inst1_n356), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_3_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_3_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S11_3_), .QN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_4_U5 ( .B1(
        DataPath_Registers_Inst1_n356), .B2(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n10), .B2(
        DataPath_Registers_Inst1_S12_4_), .C1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n11), .C2(
        DataPath_Registers_Inst1_S8_4_), .A(DataPath_Registers_Inst1_n356), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_4_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_4_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S11_4_), .QN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst1_n356), .B2(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n10), .B2(
        DataPath_Registers_Inst1_S12_5_), .C1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n11), .C2(
        DataPath_Registers_Inst1_S8_5_), .A(DataPath_Registers_Inst1_n356), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_5_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_5_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S11_5_), .QN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_5_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst1_n356), .B2(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n10), .B2(
        DataPath_Registers_Inst1_S12_6_), .C1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n11), .C2(
        DataPath_Registers_Inst1_S8_6_), .A(DataPath_Registers_Inst1_n356), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_6_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_6_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S11_6_), .QN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_6_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst1_n356), .B2(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n10), .B2(
        DataPath_Registers_Inst1_S12_7_), .C1(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n11), .C2(
        DataPath_Registers_Inst1_S8_7_), .A(DataPath_Registers_Inst1_n356), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_7_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_7_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S11_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S11_7_), .QN(
        DataPath_Registers_Inst1_ScanFF_S11_SFF_7_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_0_U5 ( .B1(
        DataPath_Registers_Inst1_n363), .B2(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n10), .B2(
        DataPath_Registers_Inst1_S14_0_), .C1(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n11), .C2(
        DataPath_Registers_Inst1_S2_0_), .A(DataPath_Registers_Inst1_n363), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_0_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_0_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_in[0]), .QN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_1_U5 ( .B1(
        DataPath_Registers_Inst1_n363), .B2(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n12), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n10), .B2(
        DataPath_Registers_Inst1_S14_1_), .C1(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n11), .C2(
        DataPath_Registers_Inst1_S2_1_), .A(DataPath_Registers_Inst1_n363), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n12) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_1_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_1_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_in[1]), .QN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst1_n363), .B2(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_2_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S14_2_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n10), .C2(
        DataPath_Registers_Inst1_S2_2_), .A(DataPath_Registers_Inst1_n363), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_2_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_in[2]), .QN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst1_n363), .B2(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_3_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S14_3_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n10), .C2(
        DataPath_Registers_Inst1_S2_3_), .A(DataPath_Registers_Inst1_n363), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_3_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_in[3]), .QN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst1_n363), .B2(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_4_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S14_4_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n10), .C2(
        DataPath_Registers_Inst1_S2_4_), .A(DataPath_Registers_Inst1_n363), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_4_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_in[4]), .QN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst1_n363), .B2(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n9), .B2(
        DataPath_Registers_Inst1_S14_5_), .C1(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n10), .C2(
        DataPath_Registers_Inst1_S2_5_), .A(DataPath_Registers_Inst1_n363), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_5_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_5_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_in[5]), .QN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_5_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst1_n363), .B2(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n9), .B2(
        DataPath_Registers_Inst1_S14_6_), .C1(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n10), .C2(
        DataPath_Registers_Inst1_S2_6_), .A(DataPath_Registers_Inst1_n363), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_6_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_6_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_in[6]), .QN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_6_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst1_n363), .B2(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n9), .B2(
        DataPath_Registers_Inst1_S14_7_), .C1(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n10), .C2(
        DataPath_Registers_Inst1_S2_7_), .A(DataPath_Registers_Inst1_n363), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_7_U3 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_7_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S13_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S12_in[7]), .QN(
        DataPath_Registers_Inst1_ScanFF_S13_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst1_n357), .B2(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_0_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S15_0_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n10), .C2(
        DataPath_Registers_Inst1_S7_0_), .A(DataPath_Registers_Inst1_n357), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_0_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S14_0_), .QN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst1_n357), .B2(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_1_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S15_1_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n10), .C2(
        DataPath_Registers_Inst1_S7_1_), .A(DataPath_Registers_Inst1_n357), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_1_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S14_1_), .QN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst1_n357), .B2(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_2_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S15_2_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n10), .C2(
        DataPath_Registers_Inst1_S7_2_), .A(DataPath_Registers_Inst1_n357), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_2_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S14_2_), .QN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst1_n357), .B2(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_3_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S15_3_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n10), .C2(
        DataPath_Registers_Inst1_S7_3_), .A(DataPath_Registers_Inst1_n357), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_3_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S14_3_), .QN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst1_n357), .B2(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_4_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S15_4_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n10), .C2(
        DataPath_Registers_Inst1_S7_4_), .A(DataPath_Registers_Inst1_n357), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_4_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S14_4_), .QN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst1_n357), .B2(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_5_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S15_5_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n10), .C2(
        DataPath_Registers_Inst1_S7_5_), .A(DataPath_Registers_Inst1_n357), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_5_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S14_5_), .QN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_5_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst1_n357), .B2(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_6_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S15_6_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n10), .C2(
        DataPath_Registers_Inst1_S7_6_), .A(DataPath_Registers_Inst1_n357), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_6_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S14_6_), .QN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_6_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst1_n357), .B2(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_7_U3 ( .B1(
        DataPath_Registers_Inst1_n351), .B2(DataPath_Registers_Inst1_S15_7_), 
        .C1(DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n10), .C2(
        DataPath_Registers_Inst1_S7_7_), .A(DataPath_Registers_Inst1_n357), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_7_U2 ( .A(
        DataPath_Registers_Inst1_n351), .ZN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S14_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S14_7_), .QN(
        DataPath_Registers_Inst1_ScanFF_S14_SFF_7_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst1_n358), .B2(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_0_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(StateIn1[0]), .C1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n10), .C2(
        DataPath_Registers_Inst1_S12_0_), .A(DataPath_Registers_Inst1_n358), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_0_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S15_0_), .QN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst1_n358), .B2(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_1_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(StateIn1[1]), .C1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n10), .C2(
        DataPath_Registers_Inst1_S12_1_), .A(DataPath_Registers_Inst1_n358), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_1_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S15_1_), .QN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst1_n358), .B2(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_2_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(StateIn1[2]), .C1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n10), .C2(
        DataPath_Registers_Inst1_S12_2_), .A(DataPath_Registers_Inst1_n358), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_2_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S15_2_), .QN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst1_n358), .B2(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_3_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(StateIn1[3]), .C1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n10), .C2(
        DataPath_Registers_Inst1_S12_3_), .A(DataPath_Registers_Inst1_n358), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_3_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S15_3_), .QN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst1_n358), .B2(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n8), .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_4_U3 ( .B1(
        DataPath_Registers_Inst1_n352), .B2(StateIn1[4]), .C1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n10), .C2(
        DataPath_Registers_Inst1_S12_4_), .A(DataPath_Registers_Inst1_n358), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_4_U2 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst1_S15_4_), .QN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst1_n358), .B2(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n9), .B2(StateIn1[5]), .C1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n10), .C2(
        DataPath_Registers_Inst1_S12_5_), .A(DataPath_Registers_Inst1_n358), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_5_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_5_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S15_5_), .QN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_5_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst1_n358), .B2(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n9), .B2(StateIn1[6]), .C1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n10), .C2(
        DataPath_Registers_Inst1_S12_6_), .A(DataPath_Registers_Inst1_n358), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_6_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_6_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S15_6_), .QN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_6_n7) );
  OAI21_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst1_n358), .B2(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n7), .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n11), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n9), .B2(StateIn1[7]), .C1(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n10), .C2(
        DataPath_Registers_Inst1_S12_7_), .A(DataPath_Registers_Inst1_n358), 
        .ZN(DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_7_U3 ( .A(
        DataPath_Registers_Inst1_n352), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_7_U2 ( .A(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n10), .ZN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst1_ScanFF_S15_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst1_S15_7_), .QN(
        DataPath_Registers_Inst1_ScanFF_S15_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U68 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n64), .A(
        DataPath_Registers_Inst1_GEN_reg1_n134), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n96) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U67 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out4[7]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n134) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U66 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n63), .A(
        DataPath_Registers_Inst1_GEN_reg1_n133), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n95) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U65 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out4[6]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n133) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U64 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n62), .A(
        DataPath_Registers_Inst1_GEN_reg1_n132), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n94) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U63 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out4[5]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n132) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U62 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n61), .A(
        DataPath_Registers_Inst1_GEN_reg1_n131), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n93) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U61 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out4[4]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n131) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U60 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n60), .A(
        DataPath_Registers_Inst1_GEN_reg1_n130), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n92) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U59 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out4[3]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n130) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U58 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n59), .A(
        DataPath_Registers_Inst1_GEN_reg1_n129), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n91) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U57 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out4[2]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n129) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U56 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n58), .A(
        DataPath_Registers_Inst1_GEN_reg1_n128), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n90) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U55 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out4[1]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n128) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U54 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n57), .A(
        DataPath_Registers_Inst1_GEN_reg1_n127), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n89) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U53 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .A2(
        DataPath_Registers_Inst1_out4[0]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n127) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U52 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n56), .A(
        DataPath_Registers_Inst1_GEN_reg1_n126), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n88) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U51 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .A2(
        DataPath_Registers_Inst1_out3[7]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n126) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U50 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n55), .A(
        DataPath_Registers_Inst1_GEN_reg1_n125), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n87) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U49 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .A2(
        DataPath_Registers_Inst1_out3[6]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n125) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U48 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n54), .A(
        DataPath_Registers_Inst1_GEN_reg1_n124), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n86) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U47 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .A2(
        DataPath_Registers_Inst1_out3[5]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n124) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U46 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n53), .A(
        DataPath_Registers_Inst1_GEN_reg1_n123), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n85) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U45 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .A2(
        DataPath_Registers_Inst1_out3[4]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n123) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U44 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n52), .A(
        DataPath_Registers_Inst1_GEN_reg1_n122), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n84) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U43 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .A2(
        DataPath_Registers_Inst1_out3[3]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n122) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U42 ( .B1(
        DataPath_Registers_Inst1_n355), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n51), .A(
        DataPath_Registers_Inst1_GEN_reg1_n121), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n83) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U41 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out3[2]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n121) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U40 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n50), .A(
        DataPath_Registers_Inst1_GEN_reg1_n120), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n82) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U39 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .A2(
        DataPath_Registers_Inst1_out3[1]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n120) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U38 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n49), .A(
        DataPath_Registers_Inst1_GEN_reg1_n119), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n81) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U37 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .A2(
        DataPath_Registers_Inst1_out3[0]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n119) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U36 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n48), .A(
        DataPath_Registers_Inst1_GEN_reg1_n118), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n80) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U35 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out2[7]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n118) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U34 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n47), .A(
        DataPath_Registers_Inst1_GEN_reg1_n117), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n79) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U33 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out2[6]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n117) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U32 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n46), .A(
        DataPath_Registers_Inst1_GEN_reg1_n116), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n78) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U31 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out2[5]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n116) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U30 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n45), .A(
        DataPath_Registers_Inst1_GEN_reg1_n115), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n77) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U29 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out2[4]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n115) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U28 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n44), .A(
        DataPath_Registers_Inst1_GEN_reg1_n114), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n76) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U27 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out2[3]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n114) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U26 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n43), .A(
        DataPath_Registers_Inst1_GEN_reg1_n113), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n75) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U25 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out2[2]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n113) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U24 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n42), .A(
        DataPath_Registers_Inst1_GEN_reg1_n112), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n74) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U23 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out2[1]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n112) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U22 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n41), .A(
        DataPath_Registers_Inst1_GEN_reg1_n111), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n73) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U21 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .A2(
        DataPath_Registers_Inst1_out2[0]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n111) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U20 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n40), .A(
        DataPath_Registers_Inst1_GEN_reg1_n110), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n72) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U19 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out1[7]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n110) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U18 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n39), .A(
        DataPath_Registers_Inst1_GEN_reg1_n109), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n71) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U17 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out1[6]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n109) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U16 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n38), .A(
        DataPath_Registers_Inst1_GEN_reg1_n108), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n70) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U15 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out1[5]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n108) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U14 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n37), .A(
        DataPath_Registers_Inst1_GEN_reg1_n107), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n69) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U13 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out1[4]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n107) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U12 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n101), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n36), .A(
        DataPath_Registers_Inst1_GEN_reg1_n106), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n68) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U11 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out1[3]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n106) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U10 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n35), .A(
        DataPath_Registers_Inst1_GEN_reg1_n105), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n67) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U9 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out1[2]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n105) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U8 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n34), .A(
        DataPath_Registers_Inst1_GEN_reg1_n104), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n66) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U7 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out1[1]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n104) );
  OAI21_X1 DataPath_Registers_Inst1_GEN_reg1_U6 ( .B1(
        DataPath_Registers_Inst1_GEN_reg1_n102), .B2(
        DataPath_Registers_Inst1_GEN_reg1_n33), .A(
        DataPath_Registers_Inst1_GEN_reg1_n103), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n65) );
  NAND2_X1 DataPath_Registers_Inst1_GEN_reg1_U5 ( .A1(
        DataPath_Registers_Inst1_GEN_reg1_n100), .A2(
        DataPath_Registers_Inst1_out1[0]), .ZN(
        DataPath_Registers_Inst1_GEN_reg1_n103) );
  BUF_X1 DataPath_Registers_Inst1_GEN_reg1_U4 ( .A(
        DataPath_Registers_Inst1_n355), .Z(
        DataPath_Registers_Inst1_GEN_reg1_n102) );
  BUF_X1 DataPath_Registers_Inst1_GEN_reg1_U3 ( .A(
        DataPath_Registers_Inst1_n355), .Z(
        DataPath_Registers_Inst1_GEN_reg1_n101) );
  BUF_X1 DataPath_Registers_Inst1_GEN_reg1_U2 ( .A(
        DataPath_Registers_Inst1_n355), .Z(
        DataPath_Registers_Inst1_GEN_reg1_n100) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_0_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n65), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output1_1[0]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n33) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_1_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n66), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output1_1[1]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n34) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_2_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n67), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output1_1[2]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n35) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_3_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n68), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output1_1[3]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n36) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_4_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n69), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output1_1[4]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n37) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_5_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n70), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output1_1[5]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n38) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_6_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n71), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output1_1[6]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n39) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_7_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n72), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output1_1[7]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n40) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_8_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n73), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output2_1[0]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n41) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_9_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n74), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output2_1[1]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n42) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_10_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n75), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output2_1[2]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n43) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_11_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n76), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output2_1[3]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n44) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_12_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n77), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output2_1[4]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n45) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_13_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n78), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output2_1[5]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n46) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_14_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n79), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output2_1[6]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n47) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_15_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n80), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output2_1[7]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n48) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_16_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n81), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output3_1[0]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n49) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_17_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n82), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output3_1[1]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n50) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_18_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n83), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output3_1[2]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n51) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_19_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n84), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output3_1[3]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n52) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_20_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n85), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output3_1[4]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n53) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_21_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n86), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output3_1[5]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n54) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_22_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n87), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output3_1[6]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n55) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_23_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n88), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output3_1[7]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n56) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_24_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n89), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output4_1[0]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n57) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_25_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n90), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output4_1[1]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n58) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_26_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n91), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output4_1[2]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n59) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_27_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n92), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output4_1[3]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n60) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_28_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n93), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output4_1[4]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n61) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_29_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n94), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output4_1[5]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n62) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_30_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n95), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output4_1[6]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n63) );
  DFF_X1 DataPath_Registers_Inst1_GEN_reg1_Q_reg_31_ ( .D(
        DataPath_Registers_Inst1_GEN_reg1_n96), .CK(clk), .Q(
        DataPath_Registers_Inst1_reg_A_output4_1[7]), .QN(
        DataPath_Registers_Inst1_GEN_reg1_n64) );
  XNOR2_X1 DataPath_Registers_Inst1_A1_U11 ( .A(
        DataPath_Registers_Inst1_in1_4_), .B(DataPath_Registers_Inst1_A1_n14), 
        .ZN(DataPath_Registers_Inst1_in1_3_) );
  XNOR2_X1 DataPath_Registers_Inst1_A1_U10 ( .A(
        DataPath_Registers_Inst1_in1_5_), .B(DataPath_Registers_Inst1_A1_n13), 
        .ZN(DataPath_Registers_Inst1_in1_2_) );
  XOR2_X1 DataPath_Registers_Inst1_A1_U9 ( .A(DataPath_Registers_Inst1_in1_7_), 
        .B(DataPath_Registers_Inst1_reg_A_output1_1[2]), .Z(
        DataPath_Registers_Inst1_A1_n13) );
  XNOR2_X1 DataPath_Registers_Inst1_A1_U8 ( .A(
        DataPath_Registers_Inst1_reg_A_output1_1[6]), .B(
        DataPath_Registers_Inst1_reg_A_output1_1[0]), .ZN(
        DataPath_Registers_Inst1_in1_5_) );
  XOR2_X1 DataPath_Registers_Inst1_A1_U7 ( .A(
        DataPath_Registers_Inst1_reg_A_output1_1[1]), .B(
        DataPath_Registers_Inst1_A1_n14), .Z(DataPath_Registers_Inst1_in1_0_)
         );
  XNOR2_X1 DataPath_Registers_Inst1_A1_U6 ( .A(
        DataPath_Registers_Inst1_reg_A_output1_1[6]), .B(
        DataPath_Registers_Inst1_reg_A_output1_1[4]), .ZN(
        DataPath_Registers_Inst1_A1_n14) );
  XNOR2_X1 DataPath_Registers_Inst1_A1_U5 ( .A(
        DataPath_Registers_Inst1_reg_A_output1_1[1]), .B(
        DataPath_Registers_Inst1_A1_n12), .ZN(DataPath_Registers_Inst1_in1_1_)
         );
  XOR2_X1 DataPath_Registers_Inst1_A1_U4 ( .A(
        DataPath_Registers_Inst1_reg_A_output1_1[5]), .B(
        DataPath_Registers_Inst1_reg_A_output1_1[4]), .Z(
        DataPath_Registers_Inst1_A1_n12) );
  XNOR2_X1 DataPath_Registers_Inst1_A1_U3 ( .A(
        DataPath_Registers_Inst1_reg_A_output1_1[5]), .B(
        DataPath_Registers_Inst1_in1_6_), .ZN(DataPath_Registers_Inst1_in1_4_)
         );
  XNOR2_X1 DataPath_Registers_Inst1_A1_U2 ( .A(
        DataPath_Registers_Inst1_reg_A_output1_1[3]), .B(
        DataPath_Registers_Inst1_reg_A_output1_1[7]), .ZN(
        DataPath_Registers_Inst1_in1_6_) );
  XOR2_X1 DataPath_Registers_Inst1_A1_U1 ( .A(
        DataPath_Registers_Inst1_reg_A_output1_1[5]), .B(
        DataPath_Registers_Inst1_reg_A_output1_1[3]), .Z(
        DataPath_Registers_Inst1_in1_7_) );
  XNOR2_X1 DataPath_Registers_Inst1_A2_U11 ( .A(
        DataPath_Registers_Inst1_in2_4_), .B(DataPath_Registers_Inst1_A2_n14), 
        .ZN(DataPath_Registers_Inst1_in2_3_) );
  XNOR2_X1 DataPath_Registers_Inst1_A2_U10 ( .A(
        DataPath_Registers_Inst1_in2_5_), .B(DataPath_Registers_Inst1_A2_n13), 
        .ZN(DataPath_Registers_Inst1_in2_2_) );
  XOR2_X1 DataPath_Registers_Inst1_A2_U9 ( .A(DataPath_Registers_Inst1_in2_7_), 
        .B(DataPath_Registers_Inst1_reg_A_output2_1[2]), .Z(
        DataPath_Registers_Inst1_A2_n13) );
  XNOR2_X1 DataPath_Registers_Inst1_A2_U8 ( .A(
        DataPath_Registers_Inst1_reg_A_output2_1[6]), .B(
        DataPath_Registers_Inst1_reg_A_output2_1[0]), .ZN(
        DataPath_Registers_Inst1_in2_5_) );
  XOR2_X1 DataPath_Registers_Inst1_A2_U7 ( .A(
        DataPath_Registers_Inst1_reg_A_output2_1[1]), .B(
        DataPath_Registers_Inst1_A2_n14), .Z(DataPath_Registers_Inst1_in2_0_)
         );
  XNOR2_X1 DataPath_Registers_Inst1_A2_U6 ( .A(
        DataPath_Registers_Inst1_reg_A_output2_1[6]), .B(
        DataPath_Registers_Inst1_reg_A_output2_1[4]), .ZN(
        DataPath_Registers_Inst1_A2_n14) );
  XNOR2_X1 DataPath_Registers_Inst1_A2_U5 ( .A(
        DataPath_Registers_Inst1_reg_A_output2_1[1]), .B(
        DataPath_Registers_Inst1_A2_n12), .ZN(DataPath_Registers_Inst1_in2_1_)
         );
  XOR2_X1 DataPath_Registers_Inst1_A2_U4 ( .A(
        DataPath_Registers_Inst1_reg_A_output2_1[5]), .B(
        DataPath_Registers_Inst1_reg_A_output2_1[4]), .Z(
        DataPath_Registers_Inst1_A2_n12) );
  XNOR2_X1 DataPath_Registers_Inst1_A2_U3 ( .A(
        DataPath_Registers_Inst1_reg_A_output2_1[5]), .B(
        DataPath_Registers_Inst1_in2_6_), .ZN(DataPath_Registers_Inst1_in2_4_)
         );
  XNOR2_X1 DataPath_Registers_Inst1_A2_U2 ( .A(
        DataPath_Registers_Inst1_reg_A_output2_1[3]), .B(
        DataPath_Registers_Inst1_reg_A_output2_1[7]), .ZN(
        DataPath_Registers_Inst1_in2_6_) );
  XOR2_X1 DataPath_Registers_Inst1_A2_U1 ( .A(
        DataPath_Registers_Inst1_reg_A_output2_1[5]), .B(
        DataPath_Registers_Inst1_reg_A_output2_1[3]), .Z(
        DataPath_Registers_Inst1_in2_7_) );
  XNOR2_X1 DataPath_Registers_Inst1_A3_U11 ( .A(
        DataPath_Registers_Inst1_in3_4_), .B(DataPath_Registers_Inst1_A3_n14), 
        .ZN(DataPath_Registers_Inst1_in3_3_) );
  XNOR2_X1 DataPath_Registers_Inst1_A3_U10 ( .A(
        DataPath_Registers_Inst1_in3_5_), .B(DataPath_Registers_Inst1_A3_n13), 
        .ZN(DataPath_Registers_Inst1_in3_2_) );
  XOR2_X1 DataPath_Registers_Inst1_A3_U9 ( .A(DataPath_Registers_Inst1_in3_7_), 
        .B(DataPath_Registers_Inst1_reg_A_output3_1[2]), .Z(
        DataPath_Registers_Inst1_A3_n13) );
  XNOR2_X1 DataPath_Registers_Inst1_A3_U8 ( .A(
        DataPath_Registers_Inst1_reg_A_output3_1[6]), .B(
        DataPath_Registers_Inst1_reg_A_output3_1[0]), .ZN(
        DataPath_Registers_Inst1_in3_5_) );
  XOR2_X1 DataPath_Registers_Inst1_A3_U7 ( .A(
        DataPath_Registers_Inst1_reg_A_output3_1[1]), .B(
        DataPath_Registers_Inst1_A3_n14), .Z(DataPath_Registers_Inst1_in3_0_)
         );
  XNOR2_X1 DataPath_Registers_Inst1_A3_U6 ( .A(
        DataPath_Registers_Inst1_reg_A_output3_1[6]), .B(
        DataPath_Registers_Inst1_reg_A_output3_1[4]), .ZN(
        DataPath_Registers_Inst1_A3_n14) );
  XNOR2_X1 DataPath_Registers_Inst1_A3_U5 ( .A(
        DataPath_Registers_Inst1_reg_A_output3_1[1]), .B(
        DataPath_Registers_Inst1_A3_n12), .ZN(DataPath_Registers_Inst1_in3_1_)
         );
  XOR2_X1 DataPath_Registers_Inst1_A3_U4 ( .A(
        DataPath_Registers_Inst1_reg_A_output3_1[5]), .B(
        DataPath_Registers_Inst1_reg_A_output3_1[4]), .Z(
        DataPath_Registers_Inst1_A3_n12) );
  XNOR2_X1 DataPath_Registers_Inst1_A3_U3 ( .A(
        DataPath_Registers_Inst1_reg_A_output3_1[5]), .B(
        DataPath_Registers_Inst1_in3_6_), .ZN(DataPath_Registers_Inst1_in3_4_)
         );
  XNOR2_X1 DataPath_Registers_Inst1_A3_U2 ( .A(
        DataPath_Registers_Inst1_reg_A_output3_1[3]), .B(
        DataPath_Registers_Inst1_reg_A_output3_1[7]), .ZN(
        DataPath_Registers_Inst1_in3_6_) );
  XOR2_X1 DataPath_Registers_Inst1_A3_U1 ( .A(
        DataPath_Registers_Inst1_reg_A_output3_1[5]), .B(
        DataPath_Registers_Inst1_reg_A_output3_1[3]), .Z(
        DataPath_Registers_Inst1_in3_7_) );
  XNOR2_X1 DataPath_Registers_Inst1_A4_U11 ( .A(
        DataPath_Registers_Inst1_in4_4_), .B(DataPath_Registers_Inst1_A4_n14), 
        .ZN(DataPath_Registers_Inst1_in4_3_) );
  XNOR2_X1 DataPath_Registers_Inst1_A4_U10 ( .A(
        DataPath_Registers_Inst1_in4_5_), .B(DataPath_Registers_Inst1_A4_n13), 
        .ZN(DataPath_Registers_Inst1_in4_2_) );
  XOR2_X1 DataPath_Registers_Inst1_A4_U9 ( .A(DataPath_Registers_Inst1_in4_7_), 
        .B(DataPath_Registers_Inst1_reg_A_output4_1[2]), .Z(
        DataPath_Registers_Inst1_A4_n13) );
  XNOR2_X1 DataPath_Registers_Inst1_A4_U8 ( .A(
        DataPath_Registers_Inst1_reg_A_output4_1[6]), .B(
        DataPath_Registers_Inst1_reg_A_output4_1[0]), .ZN(
        DataPath_Registers_Inst1_in4_5_) );
  XOR2_X1 DataPath_Registers_Inst1_A4_U7 ( .A(
        DataPath_Registers_Inst1_reg_A_output4_1[1]), .B(
        DataPath_Registers_Inst1_A4_n14), .Z(DataPath_Registers_Inst1_in4_0_)
         );
  XNOR2_X1 DataPath_Registers_Inst1_A4_U6 ( .A(
        DataPath_Registers_Inst1_reg_A_output4_1[6]), .B(
        DataPath_Registers_Inst1_reg_A_output4_1[4]), .ZN(
        DataPath_Registers_Inst1_A4_n14) );
  XNOR2_X1 DataPath_Registers_Inst1_A4_U5 ( .A(
        DataPath_Registers_Inst1_reg_A_output4_1[1]), .B(
        DataPath_Registers_Inst1_A4_n12), .ZN(DataPath_Registers_Inst1_in4_1_)
         );
  XOR2_X1 DataPath_Registers_Inst1_A4_U4 ( .A(
        DataPath_Registers_Inst1_reg_A_output4_1[5]), .B(
        DataPath_Registers_Inst1_reg_A_output4_1[4]), .Z(
        DataPath_Registers_Inst1_A4_n12) );
  XNOR2_X1 DataPath_Registers_Inst1_A4_U3 ( .A(
        DataPath_Registers_Inst1_reg_A_output4_1[5]), .B(
        DataPath_Registers_Inst1_in4_6_), .ZN(DataPath_Registers_Inst1_in4_4_)
         );
  XNOR2_X1 DataPath_Registers_Inst1_A4_U2 ( .A(
        DataPath_Registers_Inst1_reg_A_output4_1[3]), .B(
        DataPath_Registers_Inst1_reg_A_output4_1[7]), .ZN(
        DataPath_Registers_Inst1_in4_6_) );
  XOR2_X1 DataPath_Registers_Inst1_A4_U1 ( .A(
        DataPath_Registers_Inst1_reg_A_output4_1[5]), .B(
        DataPath_Registers_Inst1_reg_A_output4_1[3]), .Z(
        DataPath_Registers_Inst1_in4_7_) );
  INV_X1 DataPath_Registers_Inst2_U279 ( .A(DataPath_Registers_Inst2_n529), 
        .ZN(DataPath_Registers_Inst2_n6) );
  OAI22_X1 DataPath_Registers_Inst2_U278 ( .A1(DataPath_Registers_Inst2_n365), 
        .A2(DataPath_Registers_Inst2_n528), .B1(DataPath_Registers_Inst2_n201), 
        .B2(DataPath_Registers_Inst2_n362), .ZN(DataPath_Registers_Inst2_n529)
         );
  XOR2_X1 DataPath_Registers_Inst2_U277 ( .A(DataPath_Registers_Inst2_n527), 
        .B(DataPath_Registers_Inst2_n526), .Z(DataPath_Registers_Inst2_out4[7]) );
  XOR2_X1 DataPath_Registers_Inst2_U276 ( .A(DataPath_Registers_Inst2_n525), 
        .B(DataPath_Registers_Inst2_n524), .Z(DataPath_Registers_Inst2_out4[6]) );
  XOR2_X1 DataPath_Registers_Inst2_U275 ( .A(DataPath_Registers_Inst2_n523), 
        .B(DataPath_Registers_Inst2_n522), .Z(DataPath_Registers_Inst2_out4[5]) );
  XNOR2_X1 DataPath_Registers_Inst2_U274 ( .A(DataPath_Registers_Inst2_n521), 
        .B(DataPath_Registers_Inst2_n520), .ZN(
        DataPath_Registers_Inst2_out4[4]) );
  XNOR2_X1 DataPath_Registers_Inst2_U273 ( .A(DataPath_Registers_Inst2_n519), 
        .B(DataPath_Registers_Inst2_n518), .ZN(
        DataPath_Registers_Inst2_out4[3]) );
  XOR2_X1 DataPath_Registers_Inst2_U272 ( .A(DataPath_Registers_Inst2_n517), 
        .B(DataPath_Registers_Inst2_n516), .Z(DataPath_Registers_Inst2_out4[2]) );
  XNOR2_X1 DataPath_Registers_Inst2_U271 ( .A(DataPath_Registers_Inst2_n515), 
        .B(DataPath_Registers_Inst2_n514), .ZN(
        DataPath_Registers_Inst2_out4[1]) );
  XOR2_X1 DataPath_Registers_Inst2_U270 ( .A(DataPath_Registers_Inst2_n513), 
        .B(DataPath_Registers_Inst2_n528), .Z(DataPath_Registers_Inst2_out4[0]) );
  XNOR2_X1 DataPath_Registers_Inst2_U269 ( .A(DataPath_Registers_Inst2_n512), 
        .B(DataPath_Registers_Inst2_n511), .ZN(
        DataPath_Registers_Inst2_out3[7]) );
  XNOR2_X1 DataPath_Registers_Inst2_U268 ( .A(DataPath_Registers_Inst2_n510), 
        .B(DataPath_Registers_Inst2_n509), .ZN(
        DataPath_Registers_Inst2_out3[6]) );
  XNOR2_X1 DataPath_Registers_Inst2_U267 ( .A(DataPath_Registers_Inst2_n508), 
        .B(DataPath_Registers_Inst2_n507), .ZN(
        DataPath_Registers_Inst2_out3[5]) );
  XOR2_X1 DataPath_Registers_Inst2_U266 ( .A(DataPath_Registers_Inst2_n506), 
        .B(DataPath_Registers_Inst2_n505), .Z(DataPath_Registers_Inst2_out3[4]) );
  XOR2_X1 DataPath_Registers_Inst2_U265 ( .A(DataPath_Registers_Inst2_n504), 
        .B(DataPath_Registers_Inst2_n503), .Z(DataPath_Registers_Inst2_out3[3]) );
  XNOR2_X1 DataPath_Registers_Inst2_U264 ( .A(DataPath_Registers_Inst2_n502), 
        .B(DataPath_Registers_Inst2_n501), .ZN(
        DataPath_Registers_Inst2_out3[2]) );
  XOR2_X1 DataPath_Registers_Inst2_U263 ( .A(DataPath_Registers_Inst2_n500), 
        .B(DataPath_Registers_Inst2_n499), .Z(DataPath_Registers_Inst2_out3[1]) );
  XNOR2_X1 DataPath_Registers_Inst2_U262 ( .A(DataPath_Registers_Inst2_n498), 
        .B(DataPath_Registers_Inst2_n497), .ZN(
        DataPath_Registers_Inst2_out3[0]) );
  XNOR2_X1 DataPath_Registers_Inst2_U261 ( .A(DataPath_Registers_Inst2_n496), 
        .B(DataPath_Registers_Inst2_n512), .ZN(
        DataPath_Registers_Inst2_out2[7]) );
  XNOR2_X1 DataPath_Registers_Inst2_U260 ( .A(DataPath_Registers_Inst2_n495), 
        .B(DataPath_Registers_Inst2_n526), .ZN(DataPath_Registers_Inst2_n512)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U259 ( .A(DataPath_Registers_Inst2_n494), 
        .B(DataPath_Registers_Inst2_n510), .ZN(
        DataPath_Registers_Inst2_out2[6]) );
  XNOR2_X1 DataPath_Registers_Inst2_U258 ( .A(DataPath_Registers_Inst2_n493), 
        .B(DataPath_Registers_Inst2_n524), .ZN(DataPath_Registers_Inst2_n510)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U257 ( .A(DataPath_Registers_Inst2_n492), 
        .B(DataPath_Registers_Inst2_n508), .ZN(
        DataPath_Registers_Inst2_out2[5]) );
  XNOR2_X1 DataPath_Registers_Inst2_U256 ( .A(DataPath_Registers_Inst2_n491), 
        .B(DataPath_Registers_Inst2_n522), .ZN(DataPath_Registers_Inst2_n508)
         );
  XOR2_X1 DataPath_Registers_Inst2_U255 ( .A(DataPath_Registers_Inst2_n490), 
        .B(DataPath_Registers_Inst2_n505), .Z(DataPath_Registers_Inst2_out2[4]) );
  XNOR2_X1 DataPath_Registers_Inst2_U254 ( .A(DataPath_Registers_Inst2_n489), 
        .B(DataPath_Registers_Inst2_n520), .ZN(DataPath_Registers_Inst2_n505)
         );
  XOR2_X1 DataPath_Registers_Inst2_U253 ( .A(DataPath_Registers_Inst2_n488), 
        .B(DataPath_Registers_Inst2_n503), .Z(DataPath_Registers_Inst2_out2[3]) );
  XNOR2_X1 DataPath_Registers_Inst2_U252 ( .A(DataPath_Registers_Inst2_n487), 
        .B(DataPath_Registers_Inst2_n518), .ZN(DataPath_Registers_Inst2_n503)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U251 ( .A(DataPath_Registers_Inst2_n486), 
        .B(DataPath_Registers_Inst2_n502), .ZN(
        DataPath_Registers_Inst2_out2[2]) );
  XNOR2_X1 DataPath_Registers_Inst2_U250 ( .A(DataPath_Registers_Inst2_n485), 
        .B(DataPath_Registers_Inst2_n516), .ZN(DataPath_Registers_Inst2_n502)
         );
  XOR2_X1 DataPath_Registers_Inst2_U249 ( .A(DataPath_Registers_Inst2_n484), 
        .B(DataPath_Registers_Inst2_n499), .Z(DataPath_Registers_Inst2_out2[1]) );
  XNOR2_X1 DataPath_Registers_Inst2_U248 ( .A(DataPath_Registers_Inst2_n483), 
        .B(DataPath_Registers_Inst2_n514), .ZN(DataPath_Registers_Inst2_n499)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U247 ( .A(DataPath_Registers_Inst2_n482), 
        .B(DataPath_Registers_Inst2_n498), .ZN(
        DataPath_Registers_Inst2_out2[0]) );
  XNOR2_X1 DataPath_Registers_Inst2_U246 ( .A(DataPath_Registers_Inst2_n481), 
        .B(DataPath_Registers_Inst2_n528), .ZN(DataPath_Registers_Inst2_n498)
         );
  OAI21_X1 DataPath_Registers_Inst2_U245 ( .B1(DataPath_Registers_Inst2_n245), 
        .B2(DataPath_Registers_Inst2_n480), .A(DataPath_Registers_Inst2_n479), 
        .ZN(DataPath_Registers_Inst2_n528) );
  AOI21_X1 DataPath_Registers_Inst2_U244 ( .B1(DataPath_Registers_Inst2_n353), 
        .B2(DataPath_Registers_Inst2_S6_0_), .A(DataPath_Registers_Inst2_n478), 
        .ZN(DataPath_Registers_Inst2_n479) );
  AOI221_X1 DataPath_Registers_Inst2_U243 ( .B1(
        DataPath_Registers_Inst2_in3_7_), .B2(DataPath_Registers_Inst2_n477), 
        .C1(DataPath_Registers_Inst2_n476), .C2(DataPath_Registers_Inst2_n475), 
        .A(DataPath_Registers_Inst2_n474), .ZN(DataPath_Registers_Inst2_n478)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U242 ( .A(DataPath_Registers_Inst2_n527), 
        .B(DataPath_Registers_Inst2_n495), .ZN(
        DataPath_Registers_Inst2_out1[7]) );
  XOR2_X1 DataPath_Registers_Inst2_U241 ( .A(DataPath_Registers_Inst2_n496), 
        .B(DataPath_Registers_Inst2_n511), .Z(DataPath_Registers_Inst2_n527)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U240 ( .A(DataPath_Registers_Inst2_n525), 
        .B(DataPath_Registers_Inst2_n493), .ZN(
        DataPath_Registers_Inst2_out1[6]) );
  XOR2_X1 DataPath_Registers_Inst2_U239 ( .A(DataPath_Registers_Inst2_n494), 
        .B(DataPath_Registers_Inst2_n509), .Z(DataPath_Registers_Inst2_n525)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U238 ( .A(DataPath_Registers_Inst2_n523), 
        .B(DataPath_Registers_Inst2_n491), .ZN(
        DataPath_Registers_Inst2_out1[5]) );
  XOR2_X1 DataPath_Registers_Inst2_U237 ( .A(DataPath_Registers_Inst2_n492), 
        .B(DataPath_Registers_Inst2_n507), .Z(DataPath_Registers_Inst2_n523)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U236 ( .A(DataPath_Registers_Inst2_n521), 
        .B(DataPath_Registers_Inst2_n489), .ZN(
        DataPath_Registers_Inst2_out1[4]) );
  XOR2_X1 DataPath_Registers_Inst2_U235 ( .A(DataPath_Registers_Inst2_n506), 
        .B(DataPath_Registers_Inst2_n490), .Z(DataPath_Registers_Inst2_n521)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U234 ( .A(DataPath_Registers_Inst2_n519), 
        .B(DataPath_Registers_Inst2_n487), .ZN(
        DataPath_Registers_Inst2_out1[3]) );
  XOR2_X1 DataPath_Registers_Inst2_U233 ( .A(DataPath_Registers_Inst2_n504), 
        .B(DataPath_Registers_Inst2_n488), .Z(DataPath_Registers_Inst2_n519)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U232 ( .A(DataPath_Registers_Inst2_n517), 
        .B(DataPath_Registers_Inst2_n485), .ZN(
        DataPath_Registers_Inst2_out1[2]) );
  XOR2_X1 DataPath_Registers_Inst2_U231 ( .A(DataPath_Registers_Inst2_n486), 
        .B(DataPath_Registers_Inst2_n501), .Z(DataPath_Registers_Inst2_n517)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U230 ( .A(DataPath_Registers_Inst2_n515), 
        .B(DataPath_Registers_Inst2_n483), .ZN(
        DataPath_Registers_Inst2_out1[1]) );
  XOR2_X1 DataPath_Registers_Inst2_U229 ( .A(DataPath_Registers_Inst2_n500), 
        .B(DataPath_Registers_Inst2_n484), .Z(DataPath_Registers_Inst2_n515)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U228 ( .A(DataPath_Registers_Inst2_n513), 
        .B(DataPath_Registers_Inst2_n481), .ZN(
        DataPath_Registers_Inst2_out1[0]) );
  XOR2_X1 DataPath_Registers_Inst2_U227 ( .A(DataPath_Registers_Inst2_n482), 
        .B(DataPath_Registers_Inst2_n497), .Z(DataPath_Registers_Inst2_n513)
         );
  OAI21_X1 DataPath_Registers_Inst2_U226 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n268), .A(DataPath_Registers_Inst2_n473), 
        .ZN(DataPath_Registers_Inst2_n324) );
  NAND2_X1 DataPath_Registers_Inst2_U225 ( .A1(DataPath_Registers_Inst2_n362), 
        .A2(DataPath_Registers_Inst2_S8_in[0]), .ZN(
        DataPath_Registers_Inst2_n473) );
  INV_X1 DataPath_Registers_Inst2_U224 ( .A(DataPath_Registers_Inst2_n472), 
        .ZN(DataPath_Registers_Inst2_n323) );
  OAI22_X1 DataPath_Registers_Inst2_U223 ( .A1(DataPath_Registers_Inst2_n365), 
        .A2(DataPath_Registers_Inst2_n526), .B1(DataPath_Registers_Inst2_n203), 
        .B2(DataPath_Registers_Inst2_n361), .ZN(DataPath_Registers_Inst2_n472)
         );
  OAI222_X1 DataPath_Registers_Inst2_U222 ( .A1(DataPath_Registers_Inst2_n471), 
        .A2(DataPath_Registers_Inst2_n474), .B1(DataPath_Registers_Inst2_n480), 
        .B2(DataPath_Registers_Inst2_n266), .C1(DataPath_Registers_Inst2_n354), 
        .C2(DataPath_Registers_Inst2_n470), .ZN(DataPath_Registers_Inst2_n526)
         );
  INV_X1 DataPath_Registers_Inst2_U221 ( .A(DataPath_Registers_Inst2_S6_7_), 
        .ZN(DataPath_Registers_Inst2_n470) );
  XNOR2_X1 DataPath_Registers_Inst2_U220 ( .A(DataPath_Registers_Inst2_in3_6_), 
        .B(DataPath_Registers_Inst2_n469), .ZN(DataPath_Registers_Inst2_n471)
         );
  AOI22_X1 DataPath_Registers_Inst2_U219 ( .A1(DataPath_Registers_Inst2_in2_7_), .A2(DataPath_Registers_Inst2_in2_6_), .B1(DataPath_Registers_Inst2_n468), 
        .B2(DataPath_Registers_Inst2_n467), .ZN(DataPath_Registers_Inst2_n469)
         );
  AOI22_X1 DataPath_Registers_Inst2_U218 ( .A1(DataPath_Registers_Inst2_n360), 
        .A2(DataPath_Registers_Inst2_n495), .B1(DataPath_Registers_Inst2_n347), 
        .B2(DataPath_Registers_Inst2_n364), .ZN(DataPath_Registers_Inst2_n322)
         );
  AOI22_X1 DataPath_Registers_Inst2_U217 ( .A1(DataPath_Registers_Inst2_n466), 
        .A2(DataPath_Registers_Inst2_n465), .B1(DataPath_Registers_Inst2_n203), 
        .B2(DataPath_Registers_Inst2_n474), .ZN(DataPath_Registers_Inst2_n495)
         );
  XOR2_X1 DataPath_Registers_Inst2_U216 ( .A(DataPath_Registers_Inst2_n464), 
        .B(DataPath_Registers_Inst2_n468), .Z(DataPath_Registers_Inst2_n465)
         );
  XOR2_X1 DataPath_Registers_Inst2_U215 ( .A(DataPath_Registers_Inst2_n463), 
        .B(DataPath_Registers_Inst2_in1_6_), .Z(DataPath_Registers_Inst2_n464)
         );
  AOI22_X1 DataPath_Registers_Inst2_U214 ( .A1(DataPath_Registers_Inst2_n360), 
        .A2(DataPath_Registers_Inst2_n506), .B1(DataPath_Registers_Inst2_n264), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n321)
         );
  AOI222_X1 DataPath_Registers_Inst2_U213 ( .A1(DataPath_Registers_Inst2_S3_4_), .A2(DataPath_Registers_Inst2_n462), .B1(DataPath_Registers_Inst2_n466), .B2(
        DataPath_Registers_Inst2_n461), .C1(DataPath_Registers_Inst2_n353), 
        .C2(DataPath_Registers_Inst2_S11_4_), .ZN(
        DataPath_Registers_Inst2_n506) );
  XNOR2_X1 DataPath_Registers_Inst2_U212 ( .A(DataPath_Registers_Inst2_n460), 
        .B(DataPath_Registers_Inst2_n459), .ZN(DataPath_Registers_Inst2_n461)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U211 ( .A(DataPath_Registers_Inst2_n458), 
        .B(DataPath_Registers_Inst2_in3_4_), .ZN(DataPath_Registers_Inst2_n460) );
  OAI21_X1 DataPath_Registers_Inst2_U210 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n262), .A(DataPath_Registers_Inst2_n457), 
        .ZN(DataPath_Registers_Inst2_n320) );
  NAND2_X1 DataPath_Registers_Inst2_U209 ( .A1(DataPath_Registers_Inst2_n362), 
        .A2(DataPath_Registers_Inst2_S12_in[0]), .ZN(
        DataPath_Registers_Inst2_n457) );
  OAI21_X1 DataPath_Registers_Inst2_U208 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n261), .A(DataPath_Registers_Inst2_n456), 
        .ZN(DataPath_Registers_Inst2_n319) );
  NAND2_X1 DataPath_Registers_Inst2_U207 ( .A1(DataPath_Registers_Inst2_n362), 
        .A2(DataPath_Registers_Inst2_S12_in[1]), .ZN(
        DataPath_Registers_Inst2_n456) );
  OAI21_X1 DataPath_Registers_Inst2_U206 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n260), .A(DataPath_Registers_Inst2_n455), 
        .ZN(DataPath_Registers_Inst2_n318) );
  NAND2_X1 DataPath_Registers_Inst2_U205 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S12_in[2]), .ZN(
        DataPath_Registers_Inst2_n455) );
  OAI21_X1 DataPath_Registers_Inst2_U204 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n259), .A(DataPath_Registers_Inst2_n454), 
        .ZN(DataPath_Registers_Inst2_n317) );
  NAND2_X1 DataPath_Registers_Inst2_U203 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S12_in[3]), .ZN(
        DataPath_Registers_Inst2_n454) );
  OAI21_X1 DataPath_Registers_Inst2_U202 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n258), .A(DataPath_Registers_Inst2_n453), 
        .ZN(DataPath_Registers_Inst2_n316) );
  NAND2_X1 DataPath_Registers_Inst2_U201 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S12_in[4]), .ZN(
        DataPath_Registers_Inst2_n453) );
  OAI21_X1 DataPath_Registers_Inst2_U200 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n257), .A(DataPath_Registers_Inst2_n452), 
        .ZN(DataPath_Registers_Inst2_n315) );
  NAND2_X1 DataPath_Registers_Inst2_U199 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S12_in[5]), .ZN(
        DataPath_Registers_Inst2_n452) );
  OAI21_X1 DataPath_Registers_Inst2_U198 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n256), .A(DataPath_Registers_Inst2_n451), 
        .ZN(DataPath_Registers_Inst2_n314) );
  NAND2_X1 DataPath_Registers_Inst2_U197 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S12_in[6]), .ZN(
        DataPath_Registers_Inst2_n451) );
  OAI21_X1 DataPath_Registers_Inst2_U196 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n255), .A(DataPath_Registers_Inst2_n450), 
        .ZN(DataPath_Registers_Inst2_n313) );
  NAND2_X1 DataPath_Registers_Inst2_U195 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S12_in[7]), .ZN(
        DataPath_Registers_Inst2_n450) );
  OAI21_X1 DataPath_Registers_Inst2_U194 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n254), .A(DataPath_Registers_Inst2_n449), 
        .ZN(DataPath_Registers_Inst2_n312) );
  NAND2_X1 DataPath_Registers_Inst2_U193 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S8_in[1]), .ZN(
        DataPath_Registers_Inst2_n449) );
  OAI21_X1 DataPath_Registers_Inst2_U192 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n253), .A(DataPath_Registers_Inst2_n448), 
        .ZN(DataPath_Registers_Inst2_n311) );
  NAND2_X1 DataPath_Registers_Inst2_U191 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S8_in[2]), .ZN(
        DataPath_Registers_Inst2_n448) );
  OAI21_X1 DataPath_Registers_Inst2_U190 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n252), .A(DataPath_Registers_Inst2_n447), 
        .ZN(DataPath_Registers_Inst2_n310) );
  NAND2_X1 DataPath_Registers_Inst2_U189 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S8_in[3]), .ZN(
        DataPath_Registers_Inst2_n447) );
  OAI21_X1 DataPath_Registers_Inst2_U188 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n251), .A(DataPath_Registers_Inst2_n446), 
        .ZN(DataPath_Registers_Inst2_n309) );
  NAND2_X1 DataPath_Registers_Inst2_U187 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S8_in[4]), .ZN(
        DataPath_Registers_Inst2_n446) );
  OAI21_X1 DataPath_Registers_Inst2_U186 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n250), .A(DataPath_Registers_Inst2_n445), 
        .ZN(DataPath_Registers_Inst2_n308) );
  NAND2_X1 DataPath_Registers_Inst2_U185 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S8_in[5]), .ZN(
        DataPath_Registers_Inst2_n445) );
  OAI21_X1 DataPath_Registers_Inst2_U184 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n249), .A(DataPath_Registers_Inst2_n444), 
        .ZN(DataPath_Registers_Inst2_n307) );
  NAND2_X1 DataPath_Registers_Inst2_U183 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S8_in[6]), .ZN(
        DataPath_Registers_Inst2_n444) );
  OAI21_X1 DataPath_Registers_Inst2_U182 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n248), .A(DataPath_Registers_Inst2_n443), 
        .ZN(DataPath_Registers_Inst2_n306) );
  NAND2_X1 DataPath_Registers_Inst2_U181 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S8_in[7]), .ZN(
        DataPath_Registers_Inst2_n443) );
  MUX2_X1 DataPath_Registers_Inst2_U180 ( .A(DataPath_Registers_Inst2_S4_in[0]), .B(DataPath_Registers_Inst2_S4_0_), .S(DataPath_Registers_Inst2_n366), .Z(
        DataPath_Registers_Inst2_n305) );
  AOI22_X1 DataPath_Registers_Inst2_U179 ( .A1(DataPath_Registers_Inst2_n359), 
        .A2(DataPath_Registers_Inst2_n482), .B1(DataPath_Registers_Inst2_n246), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n304)
         );
  AOI22_X1 DataPath_Registers_Inst2_U178 ( .A1(DataPath_Registers_Inst2_n352), 
        .A2(StateIn2[0]), .B1(DataPath_Registers_Inst2_S4_0_), .B2(
        DataPath_Registers_Inst2_n354), .ZN(DataPath_Registers_Inst2_n482) );
  AOI22_X1 DataPath_Registers_Inst2_U177 ( .A1(DataPath_Registers_Inst2_n361), 
        .A2(DataPath_Registers_Inst2_n497), .B1(DataPath_Registers_Inst2_n245), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n303)
         );
  AOI22_X1 DataPath_Registers_Inst2_U176 ( .A1(DataPath_Registers_Inst2_n360), 
        .A2(DataPath_Registers_Inst2_n481), .B1(DataPath_Registers_Inst2_n346), 
        .B2(DataPath_Registers_Inst2_n364), .ZN(DataPath_Registers_Inst2_n301)
         );
  AOI22_X1 DataPath_Registers_Inst2_U175 ( .A1(DataPath_Registers_Inst2_n466), 
        .A2(DataPath_Registers_Inst2_n440), .B1(DataPath_Registers_Inst2_n201), 
        .B2(DataPath_Registers_Inst2_n474), .ZN(DataPath_Registers_Inst2_n481)
         );
  AOI22_X1 DataPath_Registers_Inst2_U174 ( .A1(DataPath_Registers_Inst2_in2_7_), .A2(DataPath_Registers_Inst2_n439), .B1(DataPath_Registers_Inst2_n438), .B2(
        DataPath_Registers_Inst2_n467), .ZN(DataPath_Registers_Inst2_n440) );
  OAI21_X1 DataPath_Registers_Inst2_U173 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n242), .A(DataPath_Registers_Inst2_n437), 
        .ZN(DataPath_Registers_Inst2_n300) );
  NAND2_X1 DataPath_Registers_Inst2_U172 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S4_in[1]), .ZN(
        DataPath_Registers_Inst2_n437) );
  AOI22_X1 DataPath_Registers_Inst2_U171 ( .A1(DataPath_Registers_Inst2_n360), 
        .A2(DataPath_Registers_Inst2_n484), .B1(DataPath_Registers_Inst2_n241), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n299)
         );
  OAI22_X1 DataPath_Registers_Inst2_U170 ( .A1(DataPath_Registers_Inst2_n354), 
        .A2(StateIn2[1]), .B1(DataPath_Registers_Inst2_S4_1_), .B2(
        DataPath_Registers_Inst2_n353), .ZN(DataPath_Registers_Inst2_n484) );
  AOI22_X1 DataPath_Registers_Inst2_U169 ( .A1(DataPath_Registers_Inst2_n359), 
        .A2(DataPath_Registers_Inst2_n500), .B1(DataPath_Registers_Inst2_n240), 
        .B2(DataPath_Registers_Inst2_n364), .ZN(DataPath_Registers_Inst2_n298)
         );
  AOI222_X1 DataPath_Registers_Inst2_U168 ( .A1(DataPath_Registers_Inst2_S3_1_), .A2(DataPath_Registers_Inst2_n462), .B1(DataPath_Registers_Inst2_n466), .B2(
        DataPath_Registers_Inst2_n436), .C1(DataPath_Registers_Inst2_n353), 
        .C2(DataPath_Registers_Inst2_S11_1_), .ZN(
        DataPath_Registers_Inst2_n500) );
  XOR2_X1 DataPath_Registers_Inst2_U167 ( .A(DataPath_Registers_Inst2_n435), 
        .B(DataPath_Registers_Inst2_n434), .Z(DataPath_Registers_Inst2_n436)
         );
  XOR2_X1 DataPath_Registers_Inst2_U166 ( .A(DataPath_Registers_Inst2_in3_1_), 
        .B(DataPath_Registers_Inst2_n442), .Z(DataPath_Registers_Inst2_n435)
         );
  AOI22_X1 DataPath_Registers_Inst2_U165 ( .A1(DataPath_Registers_Inst2_n360), 
        .A2(DataPath_Registers_Inst2_n514), .B1(DataPath_Registers_Inst2_n350), 
        .B2(DataPath_Registers_Inst2_n364), .ZN(DataPath_Registers_Inst2_n297)
         );
  AOI222_X1 DataPath_Registers_Inst2_U164 ( .A1(DataPath_Registers_Inst2_S2_1_), .A2(DataPath_Registers_Inst2_n462), .B1(DataPath_Registers_Inst2_n466), .B2(
        DataPath_Registers_Inst2_n433), .C1(DataPath_Registers_Inst2_n353), 
        .C2(DataPath_Registers_Inst2_S6_1_), .ZN(DataPath_Registers_Inst2_n514) );
  XNOR2_X1 DataPath_Registers_Inst2_U163 ( .A(DataPath_Registers_Inst2_n432), 
        .B(DataPath_Registers_Inst2_in2_1_), .ZN(DataPath_Registers_Inst2_n433) );
  XOR2_X1 DataPath_Registers_Inst2_U162 ( .A(DataPath_Registers_Inst2_n442), 
        .B(DataPath_Registers_Inst2_n477), .Z(DataPath_Registers_Inst2_n432)
         );
  INV_X1 DataPath_Registers_Inst2_U161 ( .A(DataPath_Registers_Inst2_n475), 
        .ZN(DataPath_Registers_Inst2_n477) );
  XOR2_X1 DataPath_Registers_Inst2_U160 ( .A(DataPath_Registers_Inst2_n476), 
        .B(DataPath_Registers_Inst2_in3_0_), .Z(DataPath_Registers_Inst2_n442)
         );
  AOI22_X1 DataPath_Registers_Inst2_U159 ( .A1(DataPath_Registers_Inst2_n359), 
        .A2(DataPath_Registers_Inst2_n483), .B1(DataPath_Registers_Inst2_n345), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n296)
         );
  AOI22_X1 DataPath_Registers_Inst2_U158 ( .A1(DataPath_Registers_Inst2_n466), 
        .A2(DataPath_Registers_Inst2_n431), .B1(DataPath_Registers_Inst2_n202), 
        .B2(DataPath_Registers_Inst2_n474), .ZN(DataPath_Registers_Inst2_n483)
         );
  XOR2_X1 DataPath_Registers_Inst2_U157 ( .A(DataPath_Registers_Inst2_n430), 
        .B(DataPath_Registers_Inst2_n438), .Z(DataPath_Registers_Inst2_n431)
         );
  XOR2_X1 DataPath_Registers_Inst2_U156 ( .A(DataPath_Registers_Inst2_n475), 
        .B(DataPath_Registers_Inst2_in1_1_), .Z(DataPath_Registers_Inst2_n430)
         );
  XOR2_X1 DataPath_Registers_Inst2_U155 ( .A(DataPath_Registers_Inst2_n467), 
        .B(DataPath_Registers_Inst2_in2_0_), .Z(DataPath_Registers_Inst2_n475)
         );
  MUX2_X1 DataPath_Registers_Inst2_U154 ( .A(DataPath_Registers_Inst2_S4_in[2]), .B(DataPath_Registers_Inst2_S4_2_), .S(DataPath_Registers_Inst2_n366), .Z(
        DataPath_Registers_Inst2_n295) );
  AOI22_X1 DataPath_Registers_Inst2_U153 ( .A1(DataPath_Registers_Inst2_n359), 
        .A2(DataPath_Registers_Inst2_n486), .B1(DataPath_Registers_Inst2_n236), 
        .B2(DataPath_Registers_Inst2_n364), .ZN(DataPath_Registers_Inst2_n294)
         );
  AOI22_X1 DataPath_Registers_Inst2_U152 ( .A1(DataPath_Registers_Inst2_n353), 
        .A2(StateIn2[2]), .B1(DataPath_Registers_Inst2_S4_2_), .B2(
        DataPath_Registers_Inst2_n354), .ZN(DataPath_Registers_Inst2_n486) );
  AOI22_X1 DataPath_Registers_Inst2_U151 ( .A1(DataPath_Registers_Inst2_n358), 
        .A2(DataPath_Registers_Inst2_n501), .B1(DataPath_Registers_Inst2_n235), 
        .B2(DataPath_Registers_Inst2_n364), .ZN(DataPath_Registers_Inst2_n293)
         );
  AOI222_X1 DataPath_Registers_Inst2_U150 ( .A1(DataPath_Registers_Inst2_n429), 
        .A2(DataPath_Registers_Inst2_n466), .B1(DataPath_Registers_Inst2_n462), 
        .B2(DataPath_Registers_Inst2_S3_2_), .C1(DataPath_Registers_Inst2_n353), .C2(DataPath_Registers_Inst2_S11_2_), .ZN(DataPath_Registers_Inst2_n501) );
  XOR2_X1 DataPath_Registers_Inst2_U149 ( .A(DataPath_Registers_Inst2_in4_1_), 
        .B(DataPath_Registers_Inst2_n428), .Z(DataPath_Registers_Inst2_n429)
         );
  XOR2_X1 DataPath_Registers_Inst2_U148 ( .A(DataPath_Registers_Inst2_in3_1_), 
        .B(DataPath_Registers_Inst2_in3_2_), .Z(DataPath_Registers_Inst2_n428)
         );
  INV_X1 DataPath_Registers_Inst2_U147 ( .A(DataPath_Registers_Inst2_n427), 
        .ZN(DataPath_Registers_Inst2_n292) );
  OAI22_X1 DataPath_Registers_Inst2_U146 ( .A1(DataPath_Registers_Inst2_n365), 
        .A2(DataPath_Registers_Inst2_n516), .B1(DataPath_Registers_Inst2_n212), 
        .B2(DataPath_Registers_Inst2_n361), .ZN(DataPath_Registers_Inst2_n427)
         );
  OAI222_X1 DataPath_Registers_Inst2_U145 ( .A1(DataPath_Registers_Inst2_n426), 
        .A2(DataPath_Registers_Inst2_n474), .B1(DataPath_Registers_Inst2_n480), 
        .B2(DataPath_Registers_Inst2_n235), .C1(DataPath_Registers_Inst2_n354), 
        .C2(DataPath_Registers_Inst2_n425), .ZN(DataPath_Registers_Inst2_n516)
         );
  INV_X1 DataPath_Registers_Inst2_U144 ( .A(DataPath_Registers_Inst2_S6_2_), 
        .ZN(DataPath_Registers_Inst2_n425) );
  XNOR2_X1 DataPath_Registers_Inst2_U143 ( .A(DataPath_Registers_Inst2_in2_1_), 
        .B(DataPath_Registers_Inst2_n424), .ZN(DataPath_Registers_Inst2_n426)
         );
  XOR2_X1 DataPath_Registers_Inst2_U142 ( .A(DataPath_Registers_Inst2_in3_1_), 
        .B(DataPath_Registers_Inst2_in2_2_), .Z(DataPath_Registers_Inst2_n424)
         );
  AOI22_X1 DataPath_Registers_Inst2_U141 ( .A1(DataPath_Registers_Inst2_n359), 
        .A2(DataPath_Registers_Inst2_n485), .B1(DataPath_Registers_Inst2_n344), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n291)
         );
  AOI22_X1 DataPath_Registers_Inst2_U140 ( .A1(DataPath_Registers_Inst2_n466), 
        .A2(DataPath_Registers_Inst2_n423), .B1(DataPath_Registers_Inst2_n212), 
        .B2(DataPath_Registers_Inst2_n474), .ZN(DataPath_Registers_Inst2_n485)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U139 ( .A(DataPath_Registers_Inst2_n422), 
        .B(DataPath_Registers_Inst2_in2_1_), .ZN(DataPath_Registers_Inst2_n423) );
  XNOR2_X1 DataPath_Registers_Inst2_U138 ( .A(DataPath_Registers_Inst2_in1_1_), 
        .B(DataPath_Registers_Inst2_in1_2_), .ZN(DataPath_Registers_Inst2_n422) );
  OAI21_X1 DataPath_Registers_Inst2_U137 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n232), .A(DataPath_Registers_Inst2_n421), 
        .ZN(DataPath_Registers_Inst2_n290) );
  NAND2_X1 DataPath_Registers_Inst2_U136 ( .A1(DataPath_Registers_Inst2_n363), 
        .A2(DataPath_Registers_Inst2_S4_in[3]), .ZN(
        DataPath_Registers_Inst2_n421) );
  AOI22_X1 DataPath_Registers_Inst2_U135 ( .A1(DataPath_Registers_Inst2_n358), 
        .A2(DataPath_Registers_Inst2_n488), .B1(DataPath_Registers_Inst2_n231), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n289)
         );
  OAI22_X1 DataPath_Registers_Inst2_U134 ( .A1(DataPath_Registers_Inst2_n354), 
        .A2(StateIn2[3]), .B1(DataPath_Registers_Inst2_S4_3_), .B2(
        DataPath_Registers_Inst2_n353), .ZN(DataPath_Registers_Inst2_n488) );
  AOI22_X1 DataPath_Registers_Inst2_U133 ( .A1(DataPath_Registers_Inst2_n358), 
        .A2(DataPath_Registers_Inst2_n504), .B1(DataPath_Registers_Inst2_n230), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n288)
         );
  AOI222_X1 DataPath_Registers_Inst2_U132 ( .A1(DataPath_Registers_Inst2_S3_3_), .A2(DataPath_Registers_Inst2_n462), .B1(DataPath_Registers_Inst2_n466), .B2(
        DataPath_Registers_Inst2_n420), .C1(DataPath_Registers_Inst2_n353), 
        .C2(DataPath_Registers_Inst2_S11_3_), .ZN(
        DataPath_Registers_Inst2_n504) );
  XNOR2_X1 DataPath_Registers_Inst2_U131 ( .A(DataPath_Registers_Inst2_n419), 
        .B(DataPath_Registers_Inst2_n418), .ZN(DataPath_Registers_Inst2_n420)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U130 ( .A(DataPath_Registers_Inst2_n458), 
        .B(DataPath_Registers_Inst2_in3_2_), .ZN(DataPath_Registers_Inst2_n419) );
  AOI22_X1 DataPath_Registers_Inst2_U129 ( .A1(DataPath_Registers_Inst2_n358), 
        .A2(DataPath_Registers_Inst2_n518), .B1(DataPath_Registers_Inst2_n349), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n287)
         );
  AOI222_X1 DataPath_Registers_Inst2_U128 ( .A1(DataPath_Registers_Inst2_S2_3_), .A2(DataPath_Registers_Inst2_n462), .B1(DataPath_Registers_Inst2_n466), .B2(
        DataPath_Registers_Inst2_n417), .C1(DataPath_Registers_Inst2_n353), 
        .C2(DataPath_Registers_Inst2_S6_3_), .ZN(DataPath_Registers_Inst2_n518) );
  XNOR2_X1 DataPath_Registers_Inst2_U127 ( .A(DataPath_Registers_Inst2_n416), 
        .B(DataPath_Registers_Inst2_n415), .ZN(DataPath_Registers_Inst2_n417)
         );
  XOR2_X1 DataPath_Registers_Inst2_U126 ( .A(DataPath_Registers_Inst2_n476), 
        .B(DataPath_Registers_Inst2_in3_2_), .Z(DataPath_Registers_Inst2_n415)
         );
  XOR2_X1 DataPath_Registers_Inst2_U125 ( .A(DataPath_Registers_Inst2_in2_3_), 
        .B(DataPath_Registers_Inst2_n414), .Z(DataPath_Registers_Inst2_n416)
         );
  AOI22_X1 DataPath_Registers_Inst2_U124 ( .A1(DataPath_Registers_Inst2_n358), 
        .A2(DataPath_Registers_Inst2_n487), .B1(DataPath_Registers_Inst2_n343), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n286)
         );
  AOI22_X1 DataPath_Registers_Inst2_U123 ( .A1(DataPath_Registers_Inst2_n466), 
        .A2(DataPath_Registers_Inst2_n413), .B1(DataPath_Registers_Inst2_n210), 
        .B2(DataPath_Registers_Inst2_n474), .ZN(DataPath_Registers_Inst2_n487)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U122 ( .A(DataPath_Registers_Inst2_n412), 
        .B(DataPath_Registers_Inst2_in1_2_), .ZN(DataPath_Registers_Inst2_n413) );
  XNOR2_X1 DataPath_Registers_Inst2_U121 ( .A(DataPath_Registers_Inst2_n414), 
        .B(DataPath_Registers_Inst2_n411), .ZN(DataPath_Registers_Inst2_n412)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U120 ( .A(DataPath_Registers_Inst2_n467), 
        .B(DataPath_Registers_Inst2_in2_2_), .ZN(DataPath_Registers_Inst2_n414) );
  OAI21_X1 DataPath_Registers_Inst2_U119 ( .B1(DataPath_Registers_Inst2_n363), 
        .B2(DataPath_Registers_Inst2_n227), .A(DataPath_Registers_Inst2_n410), 
        .ZN(DataPath_Registers_Inst2_n285) );
  NAND2_X1 DataPath_Registers_Inst2_U118 ( .A1(DataPath_Registers_Inst2_n362), 
        .A2(DataPath_Registers_Inst2_S4_in[4]), .ZN(
        DataPath_Registers_Inst2_n410) );
  AOI22_X1 DataPath_Registers_Inst2_U117 ( .A1(DataPath_Registers_Inst2_n357), 
        .A2(DataPath_Registers_Inst2_n490), .B1(DataPath_Registers_Inst2_n263), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n284)
         );
  OAI22_X1 DataPath_Registers_Inst2_U116 ( .A1(DataPath_Registers_Inst2_n354), 
        .A2(StateIn2[4]), .B1(DataPath_Registers_Inst2_S4_4_), .B2(
        DataPath_Registers_Inst2_n353), .ZN(DataPath_Registers_Inst2_n490) );
  MUX2_X1 DataPath_Registers_Inst2_U115 ( .A(DataPath_Registers_Inst2_S4_in[5]), .B(DataPath_Registers_Inst2_S4_5_), .S(DataPath_Registers_Inst2_n366), .Z(
        DataPath_Registers_Inst2_n283) );
  AOI22_X1 DataPath_Registers_Inst2_U114 ( .A1(DataPath_Registers_Inst2_n357), 
        .A2(DataPath_Registers_Inst2_n492), .B1(DataPath_Registers_Inst2_n225), 
        .B2(DataPath_Registers_Inst2_n364), .ZN(DataPath_Registers_Inst2_n282)
         );
  AOI22_X1 DataPath_Registers_Inst2_U113 ( .A1(DataPath_Registers_Inst2_n353), 
        .A2(StateIn2[5]), .B1(DataPath_Registers_Inst2_S4_5_), .B2(
        DataPath_Registers_Inst2_n354), .ZN(DataPath_Registers_Inst2_n492) );
  AOI22_X1 DataPath_Registers_Inst2_U112 ( .A1(DataPath_Registers_Inst2_n357), 
        .A2(DataPath_Registers_Inst2_n507), .B1(DataPath_Registers_Inst2_n224), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n281)
         );
  AOI222_X1 DataPath_Registers_Inst2_U111 ( .A1(DataPath_Registers_Inst2_n409), 
        .A2(DataPath_Registers_Inst2_n466), .B1(DataPath_Registers_Inst2_n462), 
        .B2(DataPath_Registers_Inst2_S3_5_), .C1(DataPath_Registers_Inst2_n353), .C2(DataPath_Registers_Inst2_S11_5_), .ZN(DataPath_Registers_Inst2_n507) );
  XOR2_X1 DataPath_Registers_Inst2_U110 ( .A(DataPath_Registers_Inst2_in4_4_), 
        .B(DataPath_Registers_Inst2_n408), .Z(DataPath_Registers_Inst2_n409)
         );
  XOR2_X1 DataPath_Registers_Inst2_U109 ( .A(DataPath_Registers_Inst2_in3_4_), 
        .B(DataPath_Registers_Inst2_in3_5_), .Z(DataPath_Registers_Inst2_n408)
         );
  INV_X1 DataPath_Registers_Inst2_U108 ( .A(DataPath_Registers_Inst2_n407), 
        .ZN(DataPath_Registers_Inst2_n280) );
  OAI22_X1 DataPath_Registers_Inst2_U107 ( .A1(DataPath_Registers_Inst2_n365), 
        .A2(DataPath_Registers_Inst2_n522), .B1(DataPath_Registers_Inst2_n208), 
        .B2(DataPath_Registers_Inst2_n361), .ZN(DataPath_Registers_Inst2_n407)
         );
  OAI222_X1 DataPath_Registers_Inst2_U106 ( .A1(DataPath_Registers_Inst2_n406), 
        .A2(DataPath_Registers_Inst2_n474), .B1(DataPath_Registers_Inst2_n480), 
        .B2(DataPath_Registers_Inst2_n224), .C1(DataPath_Registers_Inst2_n354), 
        .C2(DataPath_Registers_Inst2_n405), .ZN(DataPath_Registers_Inst2_n522)
         );
  INV_X1 DataPath_Registers_Inst2_U105 ( .A(DataPath_Registers_Inst2_S6_5_), 
        .ZN(DataPath_Registers_Inst2_n405) );
  XNOR2_X1 DataPath_Registers_Inst2_U104 ( .A(DataPath_Registers_Inst2_in2_5_), 
        .B(DataPath_Registers_Inst2_n404), .ZN(DataPath_Registers_Inst2_n406)
         );
  XOR2_X1 DataPath_Registers_Inst2_U103 ( .A(DataPath_Registers_Inst2_in3_4_), 
        .B(DataPath_Registers_Inst2_in2_4_), .Z(DataPath_Registers_Inst2_n404)
         );
  AOI22_X1 DataPath_Registers_Inst2_U102 ( .A1(DataPath_Registers_Inst2_n357), 
        .A2(DataPath_Registers_Inst2_n491), .B1(DataPath_Registers_Inst2_n342), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n279)
         );
  AOI22_X1 DataPath_Registers_Inst2_U101 ( .A1(DataPath_Registers_Inst2_n466), 
        .A2(DataPath_Registers_Inst2_n403), .B1(DataPath_Registers_Inst2_n208), 
        .B2(DataPath_Registers_Inst2_n474), .ZN(DataPath_Registers_Inst2_n491)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U100 ( .A(DataPath_Registers_Inst2_n402), 
        .B(DataPath_Registers_Inst2_in1_5_), .ZN(DataPath_Registers_Inst2_n403) );
  XNOR2_X1 DataPath_Registers_Inst2_U99 ( .A(DataPath_Registers_Inst2_in1_4_), 
        .B(DataPath_Registers_Inst2_in2_4_), .ZN(DataPath_Registers_Inst2_n402) );
  MUX2_X1 DataPath_Registers_Inst2_U98 ( .A(DataPath_Registers_Inst2_S4_in[6]), 
        .B(DataPath_Registers_Inst2_S4_6_), .S(DataPath_Registers_Inst2_n366), 
        .Z(DataPath_Registers_Inst2_n278) );
  AOI22_X1 DataPath_Registers_Inst2_U97 ( .A1(DataPath_Registers_Inst2_n357), 
        .A2(DataPath_Registers_Inst2_n494), .B1(DataPath_Registers_Inst2_n220), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n277)
         );
  AOI22_X1 DataPath_Registers_Inst2_U96 ( .A1(DataPath_Registers_Inst2_n353), 
        .A2(StateIn2[6]), .B1(DataPath_Registers_Inst2_S4_6_), .B2(
        DataPath_Registers_Inst2_n354), .ZN(DataPath_Registers_Inst2_n494) );
  AOI22_X1 DataPath_Registers_Inst2_U95 ( .A1(DataPath_Registers_Inst2_n356), 
        .A2(DataPath_Registers_Inst2_n509), .B1(DataPath_Registers_Inst2_n219), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n276)
         );
  AOI222_X1 DataPath_Registers_Inst2_U94 ( .A1(DataPath_Registers_Inst2_n401), 
        .A2(DataPath_Registers_Inst2_n466), .B1(DataPath_Registers_Inst2_n462), 
        .B2(DataPath_Registers_Inst2_S3_6_), .C1(DataPath_Registers_Inst2_n353), .C2(DataPath_Registers_Inst2_S11_6_), .ZN(DataPath_Registers_Inst2_n509) );
  XOR2_X1 DataPath_Registers_Inst2_U93 ( .A(DataPath_Registers_Inst2_in4_5_), 
        .B(DataPath_Registers_Inst2_n400), .Z(DataPath_Registers_Inst2_n401)
         );
  XOR2_X1 DataPath_Registers_Inst2_U92 ( .A(DataPath_Registers_Inst2_in3_5_), 
        .B(DataPath_Registers_Inst2_in3_6_), .Z(DataPath_Registers_Inst2_n400)
         );
  INV_X1 DataPath_Registers_Inst2_U91 ( .A(DataPath_Registers_Inst2_n399), 
        .ZN(DataPath_Registers_Inst2_n275) );
  OAI22_X1 DataPath_Registers_Inst2_U90 ( .A1(DataPath_Registers_Inst2_n364), 
        .A2(DataPath_Registers_Inst2_n524), .B1(DataPath_Registers_Inst2_n206), 
        .B2(DataPath_Registers_Inst2_n361), .ZN(DataPath_Registers_Inst2_n399)
         );
  OAI222_X1 DataPath_Registers_Inst2_U89 ( .A1(DataPath_Registers_Inst2_n398), 
        .A2(DataPath_Registers_Inst2_n474), .B1(DataPath_Registers_Inst2_n480), 
        .B2(DataPath_Registers_Inst2_n219), .C1(DataPath_Registers_Inst2_n354), 
        .C2(DataPath_Registers_Inst2_n397), .ZN(DataPath_Registers_Inst2_n524)
         );
  INV_X1 DataPath_Registers_Inst2_U88 ( .A(DataPath_Registers_Inst2_S6_6_), 
        .ZN(DataPath_Registers_Inst2_n397) );
  XOR2_X1 DataPath_Registers_Inst2_U87 ( .A(DataPath_Registers_Inst2_n468), 
        .B(DataPath_Registers_Inst2_n396), .Z(DataPath_Registers_Inst2_n398)
         );
  XOR2_X1 DataPath_Registers_Inst2_U86 ( .A(DataPath_Registers_Inst2_in3_5_), 
        .B(DataPath_Registers_Inst2_in2_5_), .Z(DataPath_Registers_Inst2_n396)
         );
  INV_X1 DataPath_Registers_Inst2_U85 ( .A(DataPath_Registers_Inst2_in2_6_), 
        .ZN(DataPath_Registers_Inst2_n468) );
  AOI22_X1 DataPath_Registers_Inst2_U84 ( .A1(DataPath_Registers_Inst2_n356), 
        .A2(DataPath_Registers_Inst2_n493), .B1(DataPath_Registers_Inst2_n341), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n274)
         );
  AOI22_X1 DataPath_Registers_Inst2_U83 ( .A1(DataPath_Registers_Inst2_n466), 
        .A2(DataPath_Registers_Inst2_n395), .B1(DataPath_Registers_Inst2_n206), 
        .B2(DataPath_Registers_Inst2_n474), .ZN(DataPath_Registers_Inst2_n493)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U82 ( .A(DataPath_Registers_Inst2_n394), 
        .B(DataPath_Registers_Inst2_in1_6_), .ZN(DataPath_Registers_Inst2_n395) );
  XNOR2_X1 DataPath_Registers_Inst2_U81 ( .A(DataPath_Registers_Inst2_in1_5_), 
        .B(DataPath_Registers_Inst2_in2_5_), .ZN(DataPath_Registers_Inst2_n394) );
  MUX2_X1 DataPath_Registers_Inst2_U80 ( .A(DataPath_Registers_Inst2_S4_in[7]), 
        .B(DataPath_Registers_Inst2_S4_7_), .S(DataPath_Registers_Inst2_n366), 
        .Z(DataPath_Registers_Inst2_n273) );
  AOI22_X1 DataPath_Registers_Inst2_U79 ( .A1(DataPath_Registers_Inst2_n356), 
        .A2(DataPath_Registers_Inst2_n496), .B1(DataPath_Registers_Inst2_n215), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n272)
         );
  AOI22_X1 DataPath_Registers_Inst2_U78 ( .A1(DataPath_Registers_Inst2_n351), 
        .A2(StateIn2[7]), .B1(DataPath_Registers_Inst2_S4_7_), .B2(
        DataPath_Registers_Inst2_n354), .ZN(DataPath_Registers_Inst2_n496) );
  AOI22_X1 DataPath_Registers_Inst2_U77 ( .A1(DataPath_Registers_Inst2_n356), 
        .A2(DataPath_Registers_Inst2_n511), .B1(DataPath_Registers_Inst2_n266), 
        .B2(DataPath_Registers_Inst2_n364), .ZN(DataPath_Registers_Inst2_n271)
         );
  AOI222_X1 DataPath_Registers_Inst2_U76 ( .A1(DataPath_Registers_Inst2_n393), 
        .A2(DataPath_Registers_Inst2_n466), .B1(DataPath_Registers_Inst2_n462), 
        .B2(DataPath_Registers_Inst2_S3_7_), .C1(DataPath_Registers_Inst2_n353), .C2(DataPath_Registers_Inst2_S11_7_), .ZN(DataPath_Registers_Inst2_n511) );
  XOR2_X1 DataPath_Registers_Inst2_U75 ( .A(DataPath_Registers_Inst2_in3_6_), 
        .B(DataPath_Registers_Inst2_n392), .Z(DataPath_Registers_Inst2_n393)
         );
  AOI22_X1 DataPath_Registers_Inst2_U74 ( .A1(DataPath_Registers_Inst2_in3_7_), 
        .A2(DataPath_Registers_Inst2_in4_6_), .B1(
        DataPath_Registers_Inst2_n391), .B2(DataPath_Registers_Inst2_n476), 
        .ZN(DataPath_Registers_Inst2_n392) );
  AOI22_X1 DataPath_Registers_Inst2_U73 ( .A1(DataPath_Registers_Inst2_n356), 
        .A2(DataPath_Registers_Inst2_n520), .B1(DataPath_Registers_Inst2_n348), 
        .B2(DataPath_Registers_Inst2_n365), .ZN(DataPath_Registers_Inst2_n270)
         );
  AOI222_X1 DataPath_Registers_Inst2_U72 ( .A1(DataPath_Registers_Inst2_S2_4_), 
        .A2(DataPath_Registers_Inst2_n462), .B1(DataPath_Registers_Inst2_n466), 
        .B2(DataPath_Registers_Inst2_n390), .C1(DataPath_Registers_Inst2_n353), 
        .C2(DataPath_Registers_Inst2_S6_4_), .ZN(DataPath_Registers_Inst2_n520) );
  XNOR2_X1 DataPath_Registers_Inst2_U71 ( .A(DataPath_Registers_Inst2_n389), 
        .B(DataPath_Registers_Inst2_in2_4_), .ZN(DataPath_Registers_Inst2_n390) );
  XNOR2_X1 DataPath_Registers_Inst2_U70 ( .A(DataPath_Registers_Inst2_n458), 
        .B(DataPath_Registers_Inst2_n388), .ZN(DataPath_Registers_Inst2_n389)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U69 ( .A(DataPath_Registers_Inst2_n476), 
        .B(DataPath_Registers_Inst2_in3_3_), .ZN(DataPath_Registers_Inst2_n458) );
  INV_X1 DataPath_Registers_Inst2_U68 ( .A(DataPath_Registers_Inst2_in3_7_), 
        .ZN(DataPath_Registers_Inst2_n476) );
  NAND2_X1 DataPath_Registers_Inst2_U67 ( .A1(DataPath_Registers_Inst2_n354), 
        .A2(DataPath_Registers_Inst2_n387), .ZN(DataPath_Registers_Inst2_n480)
         );
  AOI22_X1 DataPath_Registers_Inst2_U66 ( .A1(DataPath_Registers_Inst2_n355), 
        .A2(DataPath_Registers_Inst2_n489), .B1(DataPath_Registers_Inst2_n340), 
        .B2(DataPath_Registers_Inst2_n364), .ZN(DataPath_Registers_Inst2_n269)
         );
  AOI22_X1 DataPath_Registers_Inst2_U65 ( .A1(DataPath_Registers_Inst2_n466), 
        .A2(DataPath_Registers_Inst2_n386), .B1(DataPath_Registers_Inst2_n204), 
        .B2(DataPath_Registers_Inst2_n474), .ZN(DataPath_Registers_Inst2_n489)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U64 ( .A(DataPath_Registers_Inst2_n385), 
        .B(DataPath_Registers_Inst2_in1_4_), .ZN(DataPath_Registers_Inst2_n386) );
  XNOR2_X1 DataPath_Registers_Inst2_U63 ( .A(DataPath_Registers_Inst2_n411), 
        .B(DataPath_Registers_Inst2_n388), .ZN(DataPath_Registers_Inst2_n385)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U62 ( .A(DataPath_Registers_Inst2_n467), 
        .B(DataPath_Registers_Inst2_in2_3_), .ZN(DataPath_Registers_Inst2_n388) );
  INV_X1 DataPath_Registers_Inst2_U61 ( .A(DataPath_Registers_Inst2_in2_7_), 
        .ZN(DataPath_Registers_Inst2_n467) );
  AOI22_X1 DataPath_Registers_Inst2_U60 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst2_n384), .B1(DataPath_Registers_Inst2_n347), 
        .B2(DataPath_Registers_Inst2_n387), .ZN(MCout_xor_SKey_2[7]) );
  XNOR2_X1 DataPath_Registers_Inst2_U59 ( .A(DataPath_Registers_Inst2_in1_6_), 
        .B(DataPath_Registers_Inst2_n383), .ZN(DataPath_Registers_Inst2_n384)
         );
  AOI22_X1 DataPath_Registers_Inst2_U58 ( .A1(DataPath_Registers_Inst2_in4_7_), 
        .A2(DataPath_Registers_Inst2_in4_6_), .B1(
        DataPath_Registers_Inst2_n391), .B2(DataPath_Registers_Inst2_n441), 
        .ZN(DataPath_Registers_Inst2_n383) );
  AOI22_X1 DataPath_Registers_Inst2_U57 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst2_n382), .B1(DataPath_Registers_Inst2_n341), 
        .B2(DataPath_Registers_Inst2_n387), .ZN(MCout_xor_SKey_2[6]) );
  XNOR2_X1 DataPath_Registers_Inst2_U56 ( .A(DataPath_Registers_Inst2_in1_5_), 
        .B(DataPath_Registers_Inst2_n381), .ZN(DataPath_Registers_Inst2_n382)
         );
  AOI22_X1 DataPath_Registers_Inst2_U55 ( .A1(DataPath_Registers_Inst2_in4_5_), 
        .A2(DataPath_Registers_Inst2_in4_6_), .B1(
        DataPath_Registers_Inst2_n391), .B2(DataPath_Registers_Inst2_n380), 
        .ZN(DataPath_Registers_Inst2_n381) );
  INV_X1 DataPath_Registers_Inst2_U54 ( .A(DataPath_Registers_Inst2_in4_6_), 
        .ZN(DataPath_Registers_Inst2_n391) );
  AOI22_X1 DataPath_Registers_Inst2_U53 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst2_n379), .B1(DataPath_Registers_Inst2_n342), 
        .B2(DataPath_Registers_Inst2_n387), .ZN(MCout_xor_SKey_2[5]) );
  XOR2_X1 DataPath_Registers_Inst2_U52 ( .A(DataPath_Registers_Inst2_n380), 
        .B(DataPath_Registers_Inst2_n378), .Z(DataPath_Registers_Inst2_n379)
         );
  XOR2_X1 DataPath_Registers_Inst2_U51 ( .A(DataPath_Registers_Inst2_in1_4_), 
        .B(DataPath_Registers_Inst2_in4_4_), .Z(DataPath_Registers_Inst2_n378)
         );
  INV_X1 DataPath_Registers_Inst2_U50 ( .A(DataPath_Registers_Inst2_in4_5_), 
        .ZN(DataPath_Registers_Inst2_n380) );
  AOI22_X1 DataPath_Registers_Inst2_U49 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst2_n377), .B1(DataPath_Registers_Inst2_n340), 
        .B2(DataPath_Registers_Inst2_n387), .ZN(MCout_xor_SKey_2[4]) );
  XNOR2_X1 DataPath_Registers_Inst2_U48 ( .A(DataPath_Registers_Inst2_in4_4_), 
        .B(DataPath_Registers_Inst2_n376), .ZN(DataPath_Registers_Inst2_n377)
         );
  XOR2_X1 DataPath_Registers_Inst2_U47 ( .A(DataPath_Registers_Inst2_n411), 
        .B(DataPath_Registers_Inst2_n459), .Z(DataPath_Registers_Inst2_n376)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U46 ( .A(DataPath_Registers_Inst2_n441), 
        .B(DataPath_Registers_Inst2_in4_3_), .ZN(DataPath_Registers_Inst2_n459) );
  XNOR2_X1 DataPath_Registers_Inst2_U45 ( .A(DataPath_Registers_Inst2_n463), 
        .B(DataPath_Registers_Inst2_in1_3_), .ZN(DataPath_Registers_Inst2_n411) );
  AOI22_X1 DataPath_Registers_Inst2_U44 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst2_n375), .B1(DataPath_Registers_Inst2_n343), 
        .B2(DataPath_Registers_Inst2_n387), .ZN(MCout_xor_SKey_2[3]) );
  XOR2_X1 DataPath_Registers_Inst2_U43 ( .A(DataPath_Registers_Inst2_n463), 
        .B(DataPath_Registers_Inst2_n374), .Z(DataPath_Registers_Inst2_n375)
         );
  XNOR2_X1 DataPath_Registers_Inst2_U42 ( .A(DataPath_Registers_Inst2_n373), 
        .B(DataPath_Registers_Inst2_in4_3_), .ZN(DataPath_Registers_Inst2_n374) );
  XNOR2_X1 DataPath_Registers_Inst2_U41 ( .A(DataPath_Registers_Inst2_n418), 
        .B(DataPath_Registers_Inst2_in1_2_), .ZN(DataPath_Registers_Inst2_n373) );
  XNOR2_X1 DataPath_Registers_Inst2_U40 ( .A(DataPath_Registers_Inst2_n441), 
        .B(DataPath_Registers_Inst2_in4_2_), .ZN(DataPath_Registers_Inst2_n418) );
  AOI22_X1 DataPath_Registers_Inst2_U39 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst2_n372), .B1(DataPath_Registers_Inst2_n344), 
        .B2(DataPath_Registers_Inst2_n387), .ZN(MCout_xor_SKey_2[2]) );
  XNOR2_X1 DataPath_Registers_Inst2_U38 ( .A(DataPath_Registers_Inst2_in4_1_), 
        .B(DataPath_Registers_Inst2_n371), .ZN(DataPath_Registers_Inst2_n372)
         );
  XOR2_X1 DataPath_Registers_Inst2_U37 ( .A(DataPath_Registers_Inst2_in1_1_), 
        .B(DataPath_Registers_Inst2_in4_2_), .Z(DataPath_Registers_Inst2_n371)
         );
  AOI22_X1 DataPath_Registers_Inst2_U36 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst2_n370), .B1(DataPath_Registers_Inst2_n345), 
        .B2(DataPath_Registers_Inst2_n387), .ZN(MCout_xor_SKey_2[1]) );
  XNOR2_X1 DataPath_Registers_Inst2_U35 ( .A(DataPath_Registers_Inst2_in4_1_), 
        .B(DataPath_Registers_Inst2_n369), .ZN(DataPath_Registers_Inst2_n370)
         );
  AOI22_X1 DataPath_Registers_Inst2_U34 ( .A1(DataPath_Registers_Inst2_n368), 
        .A2(DataPath_Registers_Inst2_n439), .B1(DataPath_Registers_Inst2_n438), 
        .B2(DataPath_Registers_Inst2_n434), .ZN(DataPath_Registers_Inst2_n369)
         );
  INV_X1 DataPath_Registers_Inst2_U33 ( .A(DataPath_Registers_Inst2_n438), 
        .ZN(DataPath_Registers_Inst2_n439) );
  XOR2_X1 DataPath_Registers_Inst2_U32 ( .A(DataPath_Registers_Inst2_n463), 
        .B(DataPath_Registers_Inst2_in1_0_), .Z(DataPath_Registers_Inst2_n438)
         );
  AOI22_X1 DataPath_Registers_Inst2_U31 ( .A1(DoMC), .A2(
        DataPath_Registers_Inst2_n367), .B1(DataPath_Registers_Inst2_n346), 
        .B2(DataPath_Registers_Inst2_n387), .ZN(MCout_xor_SKey_2[0]) );
  INV_X1 DataPath_Registers_Inst2_U30 ( .A(DoMC), .ZN(
        DataPath_Registers_Inst2_n387) );
  AOI22_X1 DataPath_Registers_Inst2_U29 ( .A1(DataPath_Registers_Inst2_n368), 
        .A2(DataPath_Registers_Inst2_n463), .B1(
        DataPath_Registers_Inst2_in1_7_), .B2(DataPath_Registers_Inst2_n434), 
        .ZN(DataPath_Registers_Inst2_n367) );
  INV_X1 DataPath_Registers_Inst2_U28 ( .A(DataPath_Registers_Inst2_in1_7_), 
        .ZN(DataPath_Registers_Inst2_n463) );
  INV_X1 DataPath_Registers_Inst2_U27 ( .A(DataPath_Registers_Inst2_n434), 
        .ZN(DataPath_Registers_Inst2_n368) );
  XOR2_X1 DataPath_Registers_Inst2_U26 ( .A(DataPath_Registers_Inst2_n441), 
        .B(DataPath_Registers_Inst2_in4_0_), .Z(DataPath_Registers_Inst2_n434)
         );
  INV_X1 DataPath_Registers_Inst2_U25 ( .A(DataPath_Registers_Inst2_in4_7_), 
        .ZN(DataPath_Registers_Inst2_n441) );
  INV_X2 DataPath_Registers_Inst2_U24 ( .A(DataPath_Registers_Inst2_n354), 
        .ZN(DataPath_Registers_Inst2_n353) );
  INV_X1 DataPath_Registers_Inst2_U23 ( .A(DataPath_Registers_Inst2_n480), 
        .ZN(DataPath_Registers_Inst2_n462) );
  NAND2_X1 DataPath_Registers_Inst2_U22 ( .A1(DataPath_Registers_Inst2_n354), 
        .A2(DoMC), .ZN(DataPath_Registers_Inst2_n474) );
  INV_X1 DataPath_Registers_Inst2_U21 ( .A(DataPath_Registers_Inst2_n474), 
        .ZN(DataPath_Registers_Inst2_n466) );
  INV_X2 DataPath_Registers_Inst2_U20 ( .A(DataPath_Registers_Inst2_n354), 
        .ZN(DataPath_Registers_Inst2_n351) );
  INV_X2 DataPath_Registers_Inst2_U19 ( .A(DataPath_Registers_Inst2_n354), 
        .ZN(DataPath_Registers_Inst2_n352) );
  INV_X1 DataPath_Registers_Inst2_U18 ( .A(DataPath_Registers_Inst2_n366), 
        .ZN(DataPath_Registers_Inst2_n360) );
  INV_X1 DataPath_Registers_Inst2_U17 ( .A(DataPath_Registers_Inst2_n366), 
        .ZN(DataPath_Registers_Inst2_n358) );
  INV_X1 DataPath_Registers_Inst2_U16 ( .A(DataPath_Registers_Inst2_n366), 
        .ZN(DataPath_Registers_Inst2_n359) );
  INV_X1 DataPath_Registers_Inst2_U15 ( .A(DataPath_Registers_Inst2_n366), 
        .ZN(DataPath_Registers_Inst2_n356) );
  INV_X1 DataPath_Registers_Inst2_U14 ( .A(DataPath_Registers_Inst2_n366), 
        .ZN(DataPath_Registers_Inst2_n357) );
  INV_X1 DataPath_Registers_Inst2_U13 ( .A(DataPath_Registers_Inst2_n366), 
        .ZN(DataPath_Registers_Inst2_n362) );
  INV_X1 DataPath_Registers_Inst2_U12 ( .A(DataPath_Registers_Inst2_n366), 
        .ZN(DataPath_Registers_Inst2_n361) );
  INV_X2 DataPath_Registers_Inst2_U11 ( .A(DataPath_Registers_Inst2_n366), 
        .ZN(DataPath_Registers_Inst2_n363) );
  INV_X1 DataPath_Registers_Inst2_U10 ( .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst2_n365) );
  BUF_X1 DataPath_Registers_Inst2_U9 ( .A(DataPath_Registers_Inst2_n365), .Z(
        DataPath_Registers_Inst2_n364) );
  INV_X1 DataPath_Registers_Inst2_U8 ( .A(DataPath_Registers_Inst2_n364), .ZN(
        DataPath_Registers_Inst2_n355) );
  INV_X1 DataPath_Registers_Inst2_U7 ( .A(DoSR), .ZN(
        DataPath_Registers_Inst2_n354) );
  INV_X1 DataPath_Registers_Inst2_U6 ( .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst2_n366) );
  AOI211_X1 DataPath_Registers_Inst2_U5 ( .C1(DataPath_Registers_Inst2_S11_0_), 
        .C2(DataPath_Registers_Inst2_n353), .A(DataPath_Registers_Inst2_n337), 
        .B(DataPath_Registers_Inst2_n339), .ZN(DataPath_Registers_Inst2_n497)
         );
  AOI221_X1 DataPath_Registers_Inst2_U4 ( .B1(DataPath_Registers_Inst2_in4_7_), 
        .B2(DataPath_Registers_Inst2_n338), .C1(DataPath_Registers_Inst2_n441), 
        .C2(DataPath_Registers_Inst2_n442), .A(DataPath_Registers_Inst2_n474), 
        .ZN(DataPath_Registers_Inst2_n339) );
  INV_X1 DataPath_Registers_Inst2_U3 ( .A(DataPath_Registers_Inst2_n442), .ZN(
        DataPath_Registers_Inst2_n338) );
  NOR2_X1 DataPath_Registers_Inst2_U2 ( .A1(DataPath_Registers_Inst2_n480), 
        .A2(DataPath_Registers_Inst2_n246), .ZN(DataPath_Registers_Inst2_n337)
         );
  DFF_X1 DataPath_Registers_Inst2_S3_reg_1_ ( .D(DataPath_Registers_Inst2_n299), .CK(clk), .Q(DataPath_Registers_Inst2_S3_1_), .QN(
        DataPath_Registers_Inst2_n241) );
  DFF_X1 DataPath_Registers_Inst2_S3_reg_3_ ( .D(DataPath_Registers_Inst2_n289), .CK(clk), .Q(DataPath_Registers_Inst2_S3_3_), .QN(
        DataPath_Registers_Inst2_n231) );
  DFF_X1 DataPath_Registers_Inst2_S3_reg_4_ ( .D(DataPath_Registers_Inst2_n284), .CK(clk), .Q(DataPath_Registers_Inst2_S3_4_), .QN(
        DataPath_Registers_Inst2_n263) );
  DFF_X1 DataPath_Registers_Inst2_S3_reg_6_ ( .D(DataPath_Registers_Inst2_n277), .CK(clk), .Q(DataPath_Registers_Inst2_S3_6_), .QN(
        DataPath_Registers_Inst2_n220) );
  DFF_X1 DataPath_Registers_Inst2_S3_reg_7_ ( .D(DataPath_Registers_Inst2_n272), .CK(clk), .Q(DataPath_Registers_Inst2_S3_7_), .QN(
        DataPath_Registers_Inst2_n215) );
  DFF_X1 DataPath_Registers_Inst2_S3_reg_2_ ( .D(DataPath_Registers_Inst2_n294), .CK(clk), .Q(DataPath_Registers_Inst2_S3_2_), .QN(
        DataPath_Registers_Inst2_n236) );
  DFF_X1 DataPath_Registers_Inst2_S3_reg_5_ ( .D(DataPath_Registers_Inst2_n282), .CK(clk), .Q(DataPath_Registers_Inst2_S3_5_), .QN(
        DataPath_Registers_Inst2_n225) );
  DFF_X1 DataPath_Registers_Inst2_S12_reg_0_ ( .D(
        DataPath_Registers_Inst2_n320), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_0_), .QN(DataPath_Registers_Inst2_n262)
         );
  DFF_X1 DataPath_Registers_Inst2_S12_reg_1_ ( .D(
        DataPath_Registers_Inst2_n319), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_1_), .QN(DataPath_Registers_Inst2_n261)
         );
  DFF_X1 DataPath_Registers_Inst2_S12_reg_2_ ( .D(
        DataPath_Registers_Inst2_n318), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_2_), .QN(DataPath_Registers_Inst2_n260)
         );
  DFF_X1 DataPath_Registers_Inst2_S12_reg_3_ ( .D(
        DataPath_Registers_Inst2_n317), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_3_), .QN(DataPath_Registers_Inst2_n259)
         );
  DFF_X1 DataPath_Registers_Inst2_S12_reg_4_ ( .D(
        DataPath_Registers_Inst2_n316), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_4_), .QN(DataPath_Registers_Inst2_n258)
         );
  DFF_X1 DataPath_Registers_Inst2_S12_reg_5_ ( .D(
        DataPath_Registers_Inst2_n315), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_5_), .QN(DataPath_Registers_Inst2_n257)
         );
  DFF_X1 DataPath_Registers_Inst2_S12_reg_7_ ( .D(
        DataPath_Registers_Inst2_n313), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_7_), .QN(DataPath_Registers_Inst2_n255)
         );
  DFF_X1 DataPath_Registers_Inst2_S8_reg_1_ ( .D(DataPath_Registers_Inst2_n312), .CK(clk), .Q(DataPath_Registers_Inst2_S8_1_), .QN(
        DataPath_Registers_Inst2_n254) );
  DFF_X1 DataPath_Registers_Inst2_S8_reg_2_ ( .D(DataPath_Registers_Inst2_n311), .CK(clk), .Q(DataPath_Registers_Inst2_S8_2_), .QN(
        DataPath_Registers_Inst2_n253) );
  DFF_X1 DataPath_Registers_Inst2_S8_reg_3_ ( .D(DataPath_Registers_Inst2_n310), .CK(clk), .Q(DataPath_Registers_Inst2_S8_3_), .QN(
        DataPath_Registers_Inst2_n252) );
  DFF_X1 DataPath_Registers_Inst2_S8_reg_4_ ( .D(DataPath_Registers_Inst2_n309), .CK(clk), .Q(DataPath_Registers_Inst2_S8_4_), .QN(
        DataPath_Registers_Inst2_n251) );
  DFF_X1 DataPath_Registers_Inst2_S8_reg_6_ ( .D(DataPath_Registers_Inst2_n307), .CK(clk), .Q(DataPath_Registers_Inst2_S8_6_), .QN(
        DataPath_Registers_Inst2_n249) );
  DFF_X1 DataPath_Registers_Inst2_S12_reg_6_ ( .D(
        DataPath_Registers_Inst2_n314), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_6_), .QN(DataPath_Registers_Inst2_n256)
         );
  DFF_X1 DataPath_Registers_Inst2_S0_reg_2_ ( .D(DataPath_Registers_Inst2_n291), .CK(clk), .Q(), .QN(DataPath_Registers_Inst2_n344) );
  DFF_X1 DataPath_Registers_Inst2_S0_reg_3_ ( .D(DataPath_Registers_Inst2_n286), .CK(clk), .Q(), .QN(DataPath_Registers_Inst2_n343) );
  DFF_X1 DataPath_Registers_Inst2_S0_reg_5_ ( .D(DataPath_Registers_Inst2_n279), .CK(clk), .Q(), .QN(DataPath_Registers_Inst2_n342) );
  DFF_X1 DataPath_Registers_Inst2_S0_reg_6_ ( .D(DataPath_Registers_Inst2_n274), .CK(clk), .Q(), .QN(DataPath_Registers_Inst2_n341) );
  DFF_X1 DataPath_Registers_Inst2_S0_reg_4_ ( .D(DataPath_Registers_Inst2_n269), .CK(clk), .Q(), .QN(DataPath_Registers_Inst2_n340) );
  DFF_X1 DataPath_Registers_Inst2_S1_reg_4_ ( .D(DataPath_Registers_Inst2_n270), .CK(clk), .Q(DataPath_Registers_Inst2_n204), .QN(
        DataPath_Registers_Inst2_n348) );
  DFF_X1 DataPath_Registers_Inst2_S2_reg_7_ ( .D(DataPath_Registers_Inst2_n271), .CK(clk), .Q(DataPath_Registers_Inst2_S2_7_), .QN(
        DataPath_Registers_Inst2_n266) );
  DFF_X1 DataPath_Registers_Inst2_S4_reg_7_ ( .D(DataPath_Registers_Inst2_n273), .CK(clk), .Q(DataPath_Registers_Inst2_S4_7_), .QN() );
  DFF_X1 DataPath_Registers_Inst2_S1_reg_6_ ( .D(DataPath_Registers_Inst2_n275), .CK(clk), .Q(DataPath_Registers_Inst2_n206), .QN() );
  DFF_X1 DataPath_Registers_Inst2_S2_reg_6_ ( .D(DataPath_Registers_Inst2_n276), .CK(clk), .Q(DataPath_Registers_Inst2_S2_6_), .QN(
        DataPath_Registers_Inst2_n219) );
  DFF_X1 DataPath_Registers_Inst2_S4_reg_6_ ( .D(DataPath_Registers_Inst2_n278), .CK(clk), .Q(DataPath_Registers_Inst2_S4_6_), .QN() );
  DFF_X1 DataPath_Registers_Inst2_S1_reg_5_ ( .D(DataPath_Registers_Inst2_n280), .CK(clk), .Q(DataPath_Registers_Inst2_n208), .QN() );
  DFF_X1 DataPath_Registers_Inst2_S2_reg_5_ ( .D(DataPath_Registers_Inst2_n281), .CK(clk), .Q(DataPath_Registers_Inst2_S2_5_), .QN(
        DataPath_Registers_Inst2_n224) );
  DFF_X1 DataPath_Registers_Inst2_S4_reg_5_ ( .D(DataPath_Registers_Inst2_n283), .CK(clk), .Q(DataPath_Registers_Inst2_S4_5_), .QN() );
  DFF_X1 DataPath_Registers_Inst2_S4_reg_4_ ( .D(DataPath_Registers_Inst2_n285), .CK(clk), .Q(DataPath_Registers_Inst2_S4_4_), .QN(
        DataPath_Registers_Inst2_n227) );
  DFF_X1 DataPath_Registers_Inst2_S1_reg_3_ ( .D(DataPath_Registers_Inst2_n287), .CK(clk), .Q(DataPath_Registers_Inst2_n210), .QN(
        DataPath_Registers_Inst2_n349) );
  DFF_X1 DataPath_Registers_Inst2_S2_reg_3_ ( .D(DataPath_Registers_Inst2_n288), .CK(clk), .Q(DataPath_Registers_Inst2_S2_3_), .QN(
        DataPath_Registers_Inst2_n230) );
  DFF_X1 DataPath_Registers_Inst2_S4_reg_3_ ( .D(DataPath_Registers_Inst2_n290), .CK(clk), .Q(DataPath_Registers_Inst2_S4_3_), .QN(
        DataPath_Registers_Inst2_n232) );
  DFF_X1 DataPath_Registers_Inst2_S1_reg_2_ ( .D(DataPath_Registers_Inst2_n292), .CK(clk), .Q(DataPath_Registers_Inst2_n212), .QN() );
  DFF_X1 DataPath_Registers_Inst2_S2_reg_2_ ( .D(DataPath_Registers_Inst2_n293), .CK(clk), .Q(DataPath_Registers_Inst2_S2_2_), .QN(
        DataPath_Registers_Inst2_n235) );
  DFF_X1 DataPath_Registers_Inst2_S4_reg_2_ ( .D(DataPath_Registers_Inst2_n295), .CK(clk), .Q(DataPath_Registers_Inst2_S4_2_), .QN() );
  DFF_X1 DataPath_Registers_Inst2_S0_reg_1_ ( .D(DataPath_Registers_Inst2_n296), .CK(clk), .Q(), .QN(DataPath_Registers_Inst2_n345) );
  DFF_X1 DataPath_Registers_Inst2_S1_reg_1_ ( .D(DataPath_Registers_Inst2_n297), .CK(clk), .Q(DataPath_Registers_Inst2_n202), .QN(
        DataPath_Registers_Inst2_n350) );
  DFF_X1 DataPath_Registers_Inst2_S2_reg_1_ ( .D(DataPath_Registers_Inst2_n298), .CK(clk), .Q(DataPath_Registers_Inst2_S2_1_), .QN(
        DataPath_Registers_Inst2_n240) );
  DFF_X1 DataPath_Registers_Inst2_S4_reg_1_ ( .D(DataPath_Registers_Inst2_n300), .CK(clk), .Q(DataPath_Registers_Inst2_S4_1_), .QN(
        DataPath_Registers_Inst2_n242) );
  DFF_X1 DataPath_Registers_Inst2_S0_reg_0_ ( .D(DataPath_Registers_Inst2_n301), .CK(clk), .Q(), .QN(DataPath_Registers_Inst2_n346) );
  DFF_X1 DataPath_Registers_Inst2_S1_reg_0_ ( .D(DataPath_Registers_Inst2_n6), 
        .CK(clk), .Q(DataPath_Registers_Inst2_n201), .QN() );
  DFF_X1 DataPath_Registers_Inst2_S2_reg_0_ ( .D(DataPath_Registers_Inst2_n303), .CK(clk), .Q(DataPath_Registers_Inst2_S2_0_), .QN(
        DataPath_Registers_Inst2_n245) );
  DFF_X1 DataPath_Registers_Inst2_S3_reg_0_ ( .D(DataPath_Registers_Inst2_n304), .CK(clk), .Q(DataPath_Registers_Inst2_S3_0_), .QN(
        DataPath_Registers_Inst2_n246) );
  DFF_X1 DataPath_Registers_Inst2_S4_reg_0_ ( .D(DataPath_Registers_Inst2_n305), .CK(clk), .Q(DataPath_Registers_Inst2_S4_0_), .QN() );
  DFF_X1 DataPath_Registers_Inst2_S8_reg_7_ ( .D(DataPath_Registers_Inst2_n306), .CK(clk), .Q(DataPath_Registers_Inst2_S8_7_), .QN(
        DataPath_Registers_Inst2_n248) );
  DFF_X1 DataPath_Registers_Inst2_S8_reg_5_ ( .D(DataPath_Registers_Inst2_n308), .CK(clk), .Q(DataPath_Registers_Inst2_S8_5_), .QN(
        DataPath_Registers_Inst2_n250) );
  DFF_X1 DataPath_Registers_Inst2_S2_reg_4_ ( .D(DataPath_Registers_Inst2_n321), .CK(clk), .Q(DataPath_Registers_Inst2_S2_4_), .QN(
        DataPath_Registers_Inst2_n264) );
  DFF_X1 DataPath_Registers_Inst2_S0_reg_7_ ( .D(DataPath_Registers_Inst2_n322), .CK(clk), .Q(), .QN(DataPath_Registers_Inst2_n347) );
  DFF_X1 DataPath_Registers_Inst2_S1_reg_7_ ( .D(DataPath_Registers_Inst2_n323), .CK(clk), .Q(DataPath_Registers_Inst2_n203), .QN() );
  DFF_X1 DataPath_Registers_Inst2_S8_reg_0_ ( .D(DataPath_Registers_Inst2_n324), .CK(clk), .Q(DataPath_Registers_Inst2_S8_0_), .QN(
        DataPath_Registers_Inst2_n268) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_0_U5 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n10), .B2(
        DataPath_Registers_Inst2_S6_0_), .C1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n11), .C2(
        DataPath_Registers_Inst2_S10_0_), .A(DataPath_Registers_Inst2_n355), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_0_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_0_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S4_in[0]), .QN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_1_U5 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n10), .B2(
        DataPath_Registers_Inst2_S6_1_), .C1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n11), .C2(
        DataPath_Registers_Inst2_S10_1_), .A(DataPath_Registers_Inst2_n355), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_1_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_1_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S4_in[1]), .QN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_2_U5 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n10), .B2(
        DataPath_Registers_Inst2_S6_2_), .C1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n11), .C2(
        DataPath_Registers_Inst2_S10_2_), .A(DataPath_Registers_Inst2_n355), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_2_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_2_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S4_in[2]), .QN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_3_U5 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n10), .B2(
        DataPath_Registers_Inst2_S6_3_), .C1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n11), .C2(
        DataPath_Registers_Inst2_S10_3_), .A(DataPath_Registers_Inst2_n355), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_3_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_3_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S4_in[3]), .QN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_4_U5 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n10), .B2(
        DataPath_Registers_Inst2_S6_4_), .C1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n11), .C2(
        DataPath_Registers_Inst2_S10_4_), .A(DataPath_Registers_Inst2_n355), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_4_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_4_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S4_in[4]), .QN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n10), .B2(
        DataPath_Registers_Inst2_S6_5_), .C1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n11), .C2(
        DataPath_Registers_Inst2_S10_5_), .A(DataPath_Registers_Inst2_n355), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_5_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_5_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S4_in[5]), .QN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_5_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n10), .B2(
        DataPath_Registers_Inst2_S6_6_), .C1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n11), .C2(
        DataPath_Registers_Inst2_S10_6_), .A(DataPath_Registers_Inst2_n355), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_6_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_6_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S4_in[6]), .QN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_6_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n10), .B2(
        DataPath_Registers_Inst2_S6_7_), .C1(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n11), .C2(
        DataPath_Registers_Inst2_S10_7_), .A(DataPath_Registers_Inst2_n355), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_7_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_7_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S5_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S4_in[7]), .QN(
        DataPath_Registers_Inst2_ScanFF_S5_SFF_7_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_0_U5 ( .B1(
        DataPath_Registers_Inst2_n358), .B2(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n10), .B2(
        DataPath_Registers_Inst2_S7_0_), .C1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n11), .C2(
        DataPath_Registers_Inst2_S15_0_), .A(DataPath_Registers_Inst2_n358), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_0_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_0_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S6_0_), .QN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_1_U5 ( .B1(
        DataPath_Registers_Inst2_n358), .B2(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n10), .B2(
        DataPath_Registers_Inst2_S7_1_), .C1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n11), .C2(
        DataPath_Registers_Inst2_S15_1_), .A(DataPath_Registers_Inst2_n358), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_1_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_1_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S6_1_), .QN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_2_U5 ( .B1(
        DataPath_Registers_Inst2_n358), .B2(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n10), .B2(
        DataPath_Registers_Inst2_S7_2_), .C1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n11), .C2(
        DataPath_Registers_Inst2_S15_2_), .A(DataPath_Registers_Inst2_n358), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_2_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_2_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S6_2_), .QN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_3_U5 ( .B1(
        DataPath_Registers_Inst2_n358), .B2(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n10), .B2(
        DataPath_Registers_Inst2_S7_3_), .C1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n11), .C2(
        DataPath_Registers_Inst2_S15_3_), .A(DataPath_Registers_Inst2_n358), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_3_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_3_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S6_3_), .QN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_4_U5 ( .B1(
        DataPath_Registers_Inst2_n358), .B2(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n9), .B2(
        DataPath_Registers_Inst2_S7_4_), .C1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n10), .C2(
        DataPath_Registers_Inst2_S15_4_), .A(DataPath_Registers_Inst2_n358), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_4_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_4_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S6_4_), .QN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_4_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst2_n358), .B2(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n9), .B2(
        DataPath_Registers_Inst2_S7_5_), .C1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n10), .C2(
        DataPath_Registers_Inst2_S15_5_), .A(DataPath_Registers_Inst2_n358), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_5_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_5_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S6_5_), .QN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_5_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst2_n358), .B2(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n9), .B2(
        DataPath_Registers_Inst2_S7_6_), .C1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n10), .C2(
        DataPath_Registers_Inst2_S15_6_), .A(DataPath_Registers_Inst2_n358), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_6_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_6_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S6_6_), .QN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_6_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst2_n358), .B2(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n9), .B2(
        DataPath_Registers_Inst2_S7_7_), .C1(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n10), .C2(
        DataPath_Registers_Inst2_S15_7_), .A(DataPath_Registers_Inst2_n358), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_7_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_7_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S6_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S6_7_), .QN(
        DataPath_Registers_Inst2_ScanFF_S6_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_0_U5 ( .B1(
        DataPath_Registers_Inst2_n356), .B2(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n10), .B2(
        DataPath_Registers_Inst2_S8_0_), .C1(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n11), .C2(
        DataPath_Registers_Inst2_S4_0_), .A(DataPath_Registers_Inst2_n356), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_0_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_0_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S7_0_), .QN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_1_U5 ( .B1(
        DataPath_Registers_Inst2_n356), .B2(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n10), .B2(
        DataPath_Registers_Inst2_S8_1_), .C1(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n11), .C2(
        DataPath_Registers_Inst2_S4_1_), .A(DataPath_Registers_Inst2_n356), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_1_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_1_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S7_1_), .QN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_2_U5 ( .B1(
        DataPath_Registers_Inst2_n356), .B2(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n10), .B2(
        DataPath_Registers_Inst2_S8_2_), .C1(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n11), .C2(
        DataPath_Registers_Inst2_S4_2_), .A(DataPath_Registers_Inst2_n356), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_2_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_2_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S7_2_), .QN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_3_U5 ( .B1(
        DataPath_Registers_Inst2_n356), .B2(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n10), .B2(
        DataPath_Registers_Inst2_S8_3_), .C1(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n11), .C2(
        DataPath_Registers_Inst2_S4_3_), .A(DataPath_Registers_Inst2_n356), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_3_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_3_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S7_3_), .QN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_4_U5 ( .B1(
        DataPath_Registers_Inst2_n356), .B2(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n12), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n10), .B2(
        DataPath_Registers_Inst2_S8_4_), .C1(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n11), .C2(
        DataPath_Registers_Inst2_S4_4_), .A(DataPath_Registers_Inst2_n356), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n12) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_4_U3 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_4_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S7_4_), .QN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst2_n356), .B2(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_5_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S8_5_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n10), .C2(
        DataPath_Registers_Inst2_S4_5_), .A(DataPath_Registers_Inst2_n356), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_5_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S7_5_), .QN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_5_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst2_n356), .B2(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_6_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S8_6_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n10), .C2(
        DataPath_Registers_Inst2_S4_6_), .A(DataPath_Registers_Inst2_n356), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_6_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S7_6_), .QN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_6_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst2_n356), .B2(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_7_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S8_7_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n10), .C2(
        DataPath_Registers_Inst2_S4_7_), .A(DataPath_Registers_Inst2_n356), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_7_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S7_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S7_7_), .QN(
        DataPath_Registers_Inst2_ScanFF_S7_SFF_7_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst2_n359), .B2(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_0_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(DataPath_Registers_Inst2_S10_0_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n10), .C2(
        DataPath_Registers_Inst2_S14_0_), .A(DataPath_Registers_Inst2_n359), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_0_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S8_in[0]), .QN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst2_n359), .B2(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_1_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(DataPath_Registers_Inst2_S10_1_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n10), .C2(
        DataPath_Registers_Inst2_S14_1_), .A(DataPath_Registers_Inst2_n359), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_1_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S8_in[1]), .QN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst2_n359), .B2(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_2_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(DataPath_Registers_Inst2_S10_2_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n10), .C2(
        DataPath_Registers_Inst2_S14_2_), .A(DataPath_Registers_Inst2_n359), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_2_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S8_in[2]), .QN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst2_n359), .B2(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_3_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(DataPath_Registers_Inst2_S10_3_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n10), .C2(
        DataPath_Registers_Inst2_S14_3_), .A(DataPath_Registers_Inst2_n359), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_3_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S8_in[3]), .QN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst2_n359), .B2(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_4_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(DataPath_Registers_Inst2_S10_4_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n10), .C2(
        DataPath_Registers_Inst2_S14_4_), .A(DataPath_Registers_Inst2_n359), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_4_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S8_in[4]), .QN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst2_n359), .B2(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n9), .B2(
        DataPath_Registers_Inst2_S10_5_), .C1(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n10), .C2(
        DataPath_Registers_Inst2_S14_5_), .A(DataPath_Registers_Inst2_n359), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_5_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_5_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S8_in[5]), .QN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_5_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst2_n359), .B2(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n9), .B2(
        DataPath_Registers_Inst2_S10_6_), .C1(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n10), .C2(
        DataPath_Registers_Inst2_S14_6_), .A(DataPath_Registers_Inst2_n359), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_6_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_6_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S8_in[6]), .QN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_6_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst2_n359), .B2(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n9), .B2(
        DataPath_Registers_Inst2_S10_7_), .C1(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n10), .C2(
        DataPath_Registers_Inst2_S14_7_), .A(DataPath_Registers_Inst2_n359), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_7_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_7_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S9_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S8_in[7]), .QN(
        DataPath_Registers_Inst2_ScanFF_S9_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_0_U4 ( .B1(state_reg_hold), 
        .B2(DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_0_U3 ( .B1(
        DataPath_Registers_Inst2_n353), .B2(DataPath_Registers_Inst2_S11_0_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n10), .C2(
        DataPath_Registers_Inst2_S3_0_), .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_0_U2 ( .A(
        DataPath_Registers_Inst2_n353), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S10_0_), .QN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_1_U4 ( .B1(state_reg_hold), 
        .B2(DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_1_U3 ( .B1(
        DataPath_Registers_Inst2_n353), .B2(DataPath_Registers_Inst2_S11_1_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n10), .C2(
        DataPath_Registers_Inst2_S3_1_), .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_1_U2 ( .A(
        DataPath_Registers_Inst2_n353), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S10_1_), .QN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_2_U4 ( .B1(state_reg_hold), 
        .B2(DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_2_U3 ( .B1(
        DataPath_Registers_Inst2_n353), .B2(DataPath_Registers_Inst2_S11_2_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n9), .C2(
        DataPath_Registers_Inst2_S3_2_), .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_2_U2 ( .A(
        DataPath_Registers_Inst2_n353), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S10_2_), .QN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_2_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_3_U4 ( .B1(state_reg_hold), 
        .B2(DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_3_U3 ( .B1(
        DataPath_Registers_Inst2_n353), .B2(DataPath_Registers_Inst2_S11_3_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n10), .C2(
        DataPath_Registers_Inst2_S3_3_), .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_3_U2 ( .A(
        DataPath_Registers_Inst2_n353), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S10_3_), .QN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_4_U4 ( .B1(state_reg_hold), 
        .B2(DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_4_U3 ( .B1(
        DataPath_Registers_Inst2_n353), .B2(DataPath_Registers_Inst2_S11_4_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n10), .C2(
        DataPath_Registers_Inst2_S3_4_), .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_4_U2 ( .A(
        DataPath_Registers_Inst2_n353), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S10_4_), .QN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_5_U4 ( .B1(state_reg_hold), 
        .B2(DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_5_U3 ( .B1(
        DataPath_Registers_Inst2_n353), .B2(DataPath_Registers_Inst2_S11_5_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n10), .C2(
        DataPath_Registers_Inst2_S3_5_), .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_5_U2 ( .A(
        DataPath_Registers_Inst2_n353), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S10_5_), .QN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_5_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_6_U4 ( .B1(state_reg_hold), 
        .B2(DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_6_U3 ( .B1(
        DataPath_Registers_Inst2_n353), .B2(DataPath_Registers_Inst2_S11_6_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n10), .C2(
        DataPath_Registers_Inst2_S3_6_), .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_6_U2 ( .A(
        DataPath_Registers_Inst2_n353), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S10_6_), .QN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_6_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_7_U4 ( .B1(state_reg_hold), 
        .B2(DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_7_U3 ( .B1(
        DataPath_Registers_Inst2_n353), .B2(DataPath_Registers_Inst2_S11_7_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n9), .C2(
        DataPath_Registers_Inst2_S3_7_), .A(state_reg_hold), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_7_U2 ( .A(
        DataPath_Registers_Inst2_n353), .ZN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S10_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S10_7_), .QN(
        DataPath_Registers_Inst2_ScanFF_S10_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_0_U5 ( .B1(
        DataPath_Registers_Inst2_n362), .B2(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n9), .B2(
        DataPath_Registers_Inst2_S12_0_), .C1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n10), .C2(
        DataPath_Registers_Inst2_S8_0_), .A(DataPath_Registers_Inst2_n362), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_0_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_0_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S11_0_), .QN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_0_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_1_U5 ( .B1(
        DataPath_Registers_Inst2_n362), .B2(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n9), .B2(
        DataPath_Registers_Inst2_S12_1_), .C1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n10), .C2(
        DataPath_Registers_Inst2_S8_1_), .A(DataPath_Registers_Inst2_n362), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_1_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_1_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S11_1_), .QN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_1_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_2_U5 ( .B1(
        DataPath_Registers_Inst2_n362), .B2(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n9), .B2(
        DataPath_Registers_Inst2_S12_2_), .C1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n10), .C2(
        DataPath_Registers_Inst2_S8_2_), .A(DataPath_Registers_Inst2_n362), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_2_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_2_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S11_2_), .QN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_2_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_3_U5 ( .B1(
        DataPath_Registers_Inst2_n362), .B2(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n9), .B2(
        DataPath_Registers_Inst2_S12_3_), .C1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n10), .C2(
        DataPath_Registers_Inst2_S8_3_), .A(DataPath_Registers_Inst2_n362), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_3_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_3_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S11_3_), .QN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_3_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_4_U5 ( .B1(
        DataPath_Registers_Inst2_n362), .B2(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n9), .B2(
        DataPath_Registers_Inst2_S12_4_), .C1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n10), .C2(
        DataPath_Registers_Inst2_S8_4_), .A(DataPath_Registers_Inst2_n362), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_4_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_4_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S11_4_), .QN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_4_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst2_n362), .B2(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n9), .B2(
        DataPath_Registers_Inst2_S12_5_), .C1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n10), .C2(
        DataPath_Registers_Inst2_S8_5_), .A(DataPath_Registers_Inst2_n362), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_5_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_5_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S11_5_), .QN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_5_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst2_n362), .B2(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n9), .B2(
        DataPath_Registers_Inst2_S12_6_), .C1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n10), .C2(
        DataPath_Registers_Inst2_S8_6_), .A(DataPath_Registers_Inst2_n362), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_6_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_6_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S11_6_), .QN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_6_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst2_n362), .B2(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n9), .B2(
        DataPath_Registers_Inst2_S12_7_), .C1(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n10), .C2(
        DataPath_Registers_Inst2_S8_7_), .A(DataPath_Registers_Inst2_n362), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_7_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_7_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S11_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S11_7_), .QN(
        DataPath_Registers_Inst2_ScanFF_S11_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst2_n357), .B2(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_0_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S14_0_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n10), .C2(
        DataPath_Registers_Inst2_S2_0_), .A(DataPath_Registers_Inst2_n357), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_0_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_in[0]), .QN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst2_n357), .B2(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_1_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S14_1_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n10), .C2(
        DataPath_Registers_Inst2_S2_1_), .A(DataPath_Registers_Inst2_n357), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_1_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_in[1]), .QN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst2_n357), .B2(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_2_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S14_2_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n10), .C2(
        DataPath_Registers_Inst2_S2_2_), .A(DataPath_Registers_Inst2_n357), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_2_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_in[2]), .QN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst2_n357), .B2(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_3_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S14_3_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n10), .C2(
        DataPath_Registers_Inst2_S2_3_), .A(DataPath_Registers_Inst2_n357), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_3_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_in[3]), .QN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst2_n357), .B2(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_4_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S14_4_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n10), .C2(
        DataPath_Registers_Inst2_S2_4_), .A(DataPath_Registers_Inst2_n357), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_4_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_in[4]), .QN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst2_n357), .B2(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_5_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S14_5_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n10), .C2(
        DataPath_Registers_Inst2_S2_5_), .A(DataPath_Registers_Inst2_n357), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_5_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_in[5]), .QN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_5_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst2_n357), .B2(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_6_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S14_6_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n10), .C2(
        DataPath_Registers_Inst2_S2_6_), .A(DataPath_Registers_Inst2_n357), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_6_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_in[6]), .QN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_6_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst2_n357), .B2(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_7_U3 ( .B1(
        DataPath_Registers_Inst2_n351), .B2(DataPath_Registers_Inst2_S14_7_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n10), .C2(
        DataPath_Registers_Inst2_S2_7_), .A(DataPath_Registers_Inst2_n357), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_7_U2 ( .A(
        DataPath_Registers_Inst2_n351), .ZN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S13_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S12_in[7]), .QN(
        DataPath_Registers_Inst2_ScanFF_S13_SFF_7_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst2_n360), .B2(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_0_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(DataPath_Registers_Inst2_S15_0_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n10), .C2(
        DataPath_Registers_Inst2_S7_0_), .A(DataPath_Registers_Inst2_n360), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_0_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S14_0_), .QN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst2_n360), .B2(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_1_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(DataPath_Registers_Inst2_S15_1_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n10), .C2(
        DataPath_Registers_Inst2_S7_1_), .A(DataPath_Registers_Inst2_n360), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_1_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S14_1_), .QN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_1_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst2_n360), .B2(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_2_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(DataPath_Registers_Inst2_S15_2_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n10), .C2(
        DataPath_Registers_Inst2_S7_2_), .A(DataPath_Registers_Inst2_n360), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_2_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S14_2_), .QN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_2_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst2_n360), .B2(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_3_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(DataPath_Registers_Inst2_S15_3_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n10), .C2(
        DataPath_Registers_Inst2_S7_3_), .A(DataPath_Registers_Inst2_n360), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_3_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S14_3_), .QN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_3_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst2_n360), .B2(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_4_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(DataPath_Registers_Inst2_S15_4_), 
        .C1(DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n10), .C2(
        DataPath_Registers_Inst2_S7_4_), .A(DataPath_Registers_Inst2_n360), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_4_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S14_4_), .QN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_4_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst2_n360), .B2(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n9), .B2(
        DataPath_Registers_Inst2_S15_5_), .C1(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n10), .C2(
        DataPath_Registers_Inst2_S7_5_), .A(DataPath_Registers_Inst2_n360), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_5_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_5_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S14_5_), .QN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_5_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst2_n360), .B2(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n9), .B2(
        DataPath_Registers_Inst2_S15_6_), .C1(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n10), .C2(
        DataPath_Registers_Inst2_S7_6_), .A(DataPath_Registers_Inst2_n360), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_6_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_6_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S14_6_), .QN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_6_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst2_n360), .B2(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n9), .B2(
        DataPath_Registers_Inst2_S15_7_), .C1(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n10), .C2(
        DataPath_Registers_Inst2_S7_7_), .A(DataPath_Registers_Inst2_n360), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_7_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_7_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S14_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S14_7_), .QN(
        DataPath_Registers_Inst2_ScanFF_S14_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_0_U4 ( .B1(
        DataPath_Registers_Inst2_n361), .B2(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n8), .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n7) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_0_U3 ( .B1(
        DataPath_Registers_Inst2_n352), .B2(StateIn2[0]), .C1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n10), .C2(
        DataPath_Registers_Inst2_S12_0_), .A(DataPath_Registers_Inst2_n361), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_0_U2 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n10) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_0_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n7), .CK(clk), .Q(
        DataPath_Registers_Inst2_S15_0_), .QN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_0_n8) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_1_U5 ( .B1(
        DataPath_Registers_Inst2_n361), .B2(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_1_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n9), .B2(StateIn2[1]), .C1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n10), .C2(
        DataPath_Registers_Inst2_S12_1_), .A(DataPath_Registers_Inst2_n361), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_1_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_1_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_1_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S15_1_), .QN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_1_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_2_U5 ( .B1(
        DataPath_Registers_Inst2_n361), .B2(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_2_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n9), .B2(StateIn2[2]), .C1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n10), .C2(
        DataPath_Registers_Inst2_S12_2_), .A(DataPath_Registers_Inst2_n361), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_2_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_2_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_2_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S15_2_), .QN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_2_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_3_U5 ( .B1(
        DataPath_Registers_Inst2_n361), .B2(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_3_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n9), .B2(StateIn2[3]), .C1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n10), .C2(
        DataPath_Registers_Inst2_S12_3_), .A(DataPath_Registers_Inst2_n361), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_3_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_3_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_3_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S15_3_), .QN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_3_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_4_U5 ( .B1(
        DataPath_Registers_Inst2_n361), .B2(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_4_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n9), .B2(StateIn2[4]), .C1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n10), .C2(
        DataPath_Registers_Inst2_S12_4_), .A(DataPath_Registers_Inst2_n361), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_4_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_4_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_4_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S15_4_), .QN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_4_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_5_U5 ( .B1(
        DataPath_Registers_Inst2_n361), .B2(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_5_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n9), .B2(StateIn2[5]), .C1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n10), .C2(
        DataPath_Registers_Inst2_S12_5_), .A(DataPath_Registers_Inst2_n361), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_5_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_5_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_5_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S15_5_), .QN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_5_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_6_U5 ( .B1(
        DataPath_Registers_Inst2_n361), .B2(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_6_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n9), .B2(StateIn2[6]), .C1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n10), .C2(
        DataPath_Registers_Inst2_S12_6_), .A(DataPath_Registers_Inst2_n361), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_6_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_6_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_6_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S15_6_), .QN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_6_n7) );
  OAI21_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_7_U5 ( .B1(
        DataPath_Registers_Inst2_n361), .B2(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n7), .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n11), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n6) );
  OAI221_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_7_U4 ( .B1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n9), .B2(StateIn2[7]), .C1(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n10), .C2(
        DataPath_Registers_Inst2_S12_7_), .A(DataPath_Registers_Inst2_n361), 
        .ZN(DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n11) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_7_U3 ( .A(
        DataPath_Registers_Inst2_n352), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n10) );
  INV_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_7_U2 ( .A(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n10), .ZN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n9) );
  DFF_X1 DataPath_Registers_Inst2_ScanFF_S15_SFF_7_Q_reg ( .D(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n6), .CK(clk), .Q(
        DataPath_Registers_Inst2_S15_7_), .QN(
        DataPath_Registers_Inst2_ScanFF_S15_SFF_7_n7) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U68 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n163), .A(
        DataPath_Registers_Inst2_GEN_reg1_n230), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n131) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U67 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out1[0]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n230) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U66 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n162), .A(
        DataPath_Registers_Inst2_GEN_reg1_n229), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n130) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U65 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out1[1]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n229) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U64 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n161), .A(
        DataPath_Registers_Inst2_GEN_reg1_n228), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n129) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U63 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out1[2]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n228) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U62 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n160), .A(
        DataPath_Registers_Inst2_GEN_reg1_n227), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n128) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U61 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out1[3]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n227) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U60 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n159), .A(
        DataPath_Registers_Inst2_GEN_reg1_n226), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n127) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U59 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out1[4]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n226) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U58 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n158), .A(
        DataPath_Registers_Inst2_GEN_reg1_n225), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n126) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U57 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out1[5]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n225) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U56 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n157), .A(
        DataPath_Registers_Inst2_GEN_reg1_n224), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n125) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U55 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out1[6]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n224) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U54 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n156), .A(
        DataPath_Registers_Inst2_GEN_reg1_n223), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n124) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U53 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .A2(
        DataPath_Registers_Inst2_out1[7]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n223) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U52 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n155), .A(
        DataPath_Registers_Inst2_GEN_reg1_n222), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n123) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U51 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .A2(
        DataPath_Registers_Inst2_out2[0]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n222) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U50 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n154), .A(
        DataPath_Registers_Inst2_GEN_reg1_n221), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n122) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U49 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .A2(
        DataPath_Registers_Inst2_out2[1]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n221) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U48 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n153), .A(
        DataPath_Registers_Inst2_GEN_reg1_n220), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n121) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U47 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .A2(
        DataPath_Registers_Inst2_out2[2]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n220) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U46 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n152), .A(
        DataPath_Registers_Inst2_GEN_reg1_n219), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n120) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U45 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .A2(
        DataPath_Registers_Inst2_out2[3]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n219) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U44 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n151), .A(
        DataPath_Registers_Inst2_GEN_reg1_n218), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n119) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U43 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .A2(
        DataPath_Registers_Inst2_out2[4]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n218) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U42 ( .B1(
        DataPath_Registers_Inst2_n355), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n150), .A(
        DataPath_Registers_Inst2_GEN_reg1_n217), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n118) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U41 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out2[5]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n217) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U40 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n149), .A(
        DataPath_Registers_Inst2_GEN_reg1_n216), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n117) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U39 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .A2(
        DataPath_Registers_Inst2_out2[6]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n216) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U38 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n148), .A(
        DataPath_Registers_Inst2_GEN_reg1_n215), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n116) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U37 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .A2(
        DataPath_Registers_Inst2_out2[7]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n215) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U36 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n147), .A(
        DataPath_Registers_Inst2_GEN_reg1_n214), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n115) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U35 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out3[0]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n214) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U34 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n146), .A(
        DataPath_Registers_Inst2_GEN_reg1_n213), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n114) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U33 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out3[1]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n213) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U32 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n145), .A(
        DataPath_Registers_Inst2_GEN_reg1_n212), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n113) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U31 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out3[2]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n212) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U30 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n144), .A(
        DataPath_Registers_Inst2_GEN_reg1_n211), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n112) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U29 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out3[3]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n211) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U28 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n143), .A(
        DataPath_Registers_Inst2_GEN_reg1_n210), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n111) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U27 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out3[4]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n210) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U26 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n142), .A(
        DataPath_Registers_Inst2_GEN_reg1_n209), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n110) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U25 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out3[5]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n209) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U24 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n141), .A(
        DataPath_Registers_Inst2_GEN_reg1_n208), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n109) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U23 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out3[6]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n208) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U22 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n140), .A(
        DataPath_Registers_Inst2_GEN_reg1_n207), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n108) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U21 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .A2(
        DataPath_Registers_Inst2_out3[7]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n207) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U20 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n139), .A(
        DataPath_Registers_Inst2_GEN_reg1_n206), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n107) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U19 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out4[0]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n206) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U18 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n138), .A(
        DataPath_Registers_Inst2_GEN_reg1_n205), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n106) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U17 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out4[1]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n205) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U16 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n137), .A(
        DataPath_Registers_Inst2_GEN_reg1_n204), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n105) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U15 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out4[2]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n204) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U14 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n136), .A(
        DataPath_Registers_Inst2_GEN_reg1_n203), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n104) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U13 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out4[3]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n203) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U12 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n197), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n135), .A(
        DataPath_Registers_Inst2_GEN_reg1_n202), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n103) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U11 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out4[4]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n202) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U10 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n134), .A(
        DataPath_Registers_Inst2_GEN_reg1_n201), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n102) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U9 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out4[5]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n201) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U8 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n133), .A(
        DataPath_Registers_Inst2_GEN_reg1_n200), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n101) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U7 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out4[6]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n200) );
  OAI21_X1 DataPath_Registers_Inst2_GEN_reg1_U6 ( .B1(
        DataPath_Registers_Inst2_GEN_reg1_n198), .B2(
        DataPath_Registers_Inst2_GEN_reg1_n132), .A(
        DataPath_Registers_Inst2_GEN_reg1_n199), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n100) );
  NAND2_X1 DataPath_Registers_Inst2_GEN_reg1_U5 ( .A1(
        DataPath_Registers_Inst2_GEN_reg1_n196), .A2(
        DataPath_Registers_Inst2_out4[7]), .ZN(
        DataPath_Registers_Inst2_GEN_reg1_n199) );
  BUF_X1 DataPath_Registers_Inst2_GEN_reg1_U4 ( .A(
        DataPath_Registers_Inst2_n355), .Z(
        DataPath_Registers_Inst2_GEN_reg1_n197) );
  BUF_X1 DataPath_Registers_Inst2_GEN_reg1_U3 ( .A(
        DataPath_Registers_Inst2_n355), .Z(
        DataPath_Registers_Inst2_GEN_reg1_n198) );
  BUF_X1 DataPath_Registers_Inst2_GEN_reg1_U2 ( .A(
        DataPath_Registers_Inst2_n355), .Z(
        DataPath_Registers_Inst2_GEN_reg1_n196) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_0_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n131), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output1_1[0]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n163) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_1_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n130), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output1_1[1]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n162) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_2_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n129), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output1_1[2]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n161) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_3_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n128), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output1_1[3]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n160) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_4_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n127), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output1_1[4]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n159) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_5_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n126), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output1_1[5]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n158) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_6_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n125), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output1_1[6]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n157) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_7_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n124), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output1_1[7]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n156) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_8_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n123), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output2_1[0]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n155) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_9_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n122), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output2_1[1]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n154) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_10_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n121), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output2_1[2]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n153) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_11_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n120), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output2_1[3]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n152) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_12_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n119), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output2_1[4]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n151) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_13_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n118), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output2_1[5]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n150) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_14_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n117), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output2_1[6]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n149) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_15_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n116), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output2_1[7]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n148) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_16_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n115), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output3_1[0]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n147) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_17_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n114), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output3_1[1]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n146) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_18_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n113), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output3_1[2]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n145) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_19_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n112), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output3_1[3]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n144) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_20_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n111), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output3_1[4]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n143) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_21_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n110), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output3_1[5]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n142) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_22_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n109), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output3_1[6]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n141) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_23_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n108), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output3_1[7]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n140) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_24_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n107), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output4_1[0]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n139) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_25_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n106), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output4_1[1]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n138) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_26_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n105), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output4_1[2]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n137) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_27_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n104), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output4_1[3]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n136) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_28_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n103), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output4_1[4]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n135) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_29_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n102), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output4_1[5]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n134) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_30_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n101), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output4_1[6]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n133) );
  DFF_X1 DataPath_Registers_Inst2_GEN_reg1_Q_reg_31_ ( .D(
        DataPath_Registers_Inst2_GEN_reg1_n100), .CK(clk), .Q(
        DataPath_Registers_Inst2_reg_A_output4_1[7]), .QN(
        DataPath_Registers_Inst2_GEN_reg1_n132) );
  XNOR2_X1 DataPath_Registers_Inst2_A1_U11 ( .A(
        DataPath_Registers_Inst2_in1_4_), .B(DataPath_Registers_Inst2_A1_n12), 
        .ZN(DataPath_Registers_Inst2_in1_3_) );
  XNOR2_X1 DataPath_Registers_Inst2_A1_U10 ( .A(
        DataPath_Registers_Inst2_A1_n11), .B(DataPath_Registers_Inst2_in1_5_), 
        .ZN(DataPath_Registers_Inst2_in1_2_) );
  XNOR2_X1 DataPath_Registers_Inst2_A1_U9 ( .A(DataPath_Registers_Inst2_in1_7_), .B(DataPath_Registers_Inst2_reg_A_output1_1[2]), .ZN(
        DataPath_Registers_Inst2_A1_n11) );
  XOR2_X1 DataPath_Registers_Inst2_A1_U8 ( .A(
        DataPath_Registers_Inst2_reg_A_output1_1[6]), .B(
        DataPath_Registers_Inst2_reg_A_output1_1[0]), .Z(
        DataPath_Registers_Inst2_in1_5_) );
  XNOR2_X1 DataPath_Registers_Inst2_A1_U7 ( .A(DataPath_Registers_Inst2_A1_n10), .B(DataPath_Registers_Inst2_reg_A_output1_1[1]), .ZN(
        DataPath_Registers_Inst2_in1_1_) );
  XNOR2_X1 DataPath_Registers_Inst2_A1_U6 ( .A(
        DataPath_Registers_Inst2_reg_A_output1_1[5]), .B(
        DataPath_Registers_Inst2_reg_A_output1_1[4]), .ZN(
        DataPath_Registers_Inst2_A1_n10) );
  XNOR2_X1 DataPath_Registers_Inst2_A1_U5 ( .A(
        DataPath_Registers_Inst2_reg_A_output1_1[1]), .B(
        DataPath_Registers_Inst2_A1_n12), .ZN(DataPath_Registers_Inst2_in1_0_)
         );
  XNOR2_X1 DataPath_Registers_Inst2_A1_U4 ( .A(
        DataPath_Registers_Inst2_reg_A_output1_1[6]), .B(
        DataPath_Registers_Inst2_reg_A_output1_1[4]), .ZN(
        DataPath_Registers_Inst2_A1_n12) );
  XOR2_X1 DataPath_Registers_Inst2_A1_U3 ( .A(
        DataPath_Registers_Inst2_reg_A_output1_1[5]), .B(
        DataPath_Registers_Inst2_in1_6_), .Z(DataPath_Registers_Inst2_in1_4_)
         );
  XOR2_X1 DataPath_Registers_Inst2_A1_U2 ( .A(
        DataPath_Registers_Inst2_reg_A_output1_1[3]), .B(
        DataPath_Registers_Inst2_reg_A_output1_1[7]), .Z(
        DataPath_Registers_Inst2_in1_6_) );
  XOR2_X1 DataPath_Registers_Inst2_A1_U1 ( .A(
        DataPath_Registers_Inst2_reg_A_output1_1[5]), .B(
        DataPath_Registers_Inst2_reg_A_output1_1[3]), .Z(
        DataPath_Registers_Inst2_in1_7_) );
  XNOR2_X1 DataPath_Registers_Inst2_A2_U11 ( .A(
        DataPath_Registers_Inst2_in2_4_), .B(DataPath_Registers_Inst2_A2_n12), 
        .ZN(DataPath_Registers_Inst2_in2_3_) );
  XNOR2_X1 DataPath_Registers_Inst2_A2_U10 ( .A(
        DataPath_Registers_Inst2_A2_n11), .B(DataPath_Registers_Inst2_in2_5_), 
        .ZN(DataPath_Registers_Inst2_in2_2_) );
  XNOR2_X1 DataPath_Registers_Inst2_A2_U9 ( .A(DataPath_Registers_Inst2_in2_7_), .B(DataPath_Registers_Inst2_reg_A_output2_1[2]), .ZN(
        DataPath_Registers_Inst2_A2_n11) );
  XOR2_X1 DataPath_Registers_Inst2_A2_U8 ( .A(
        DataPath_Registers_Inst2_reg_A_output2_1[6]), .B(
        DataPath_Registers_Inst2_reg_A_output2_1[0]), .Z(
        DataPath_Registers_Inst2_in2_5_) );
  XNOR2_X1 DataPath_Registers_Inst2_A2_U7 ( .A(DataPath_Registers_Inst2_A2_n10), .B(DataPath_Registers_Inst2_reg_A_output2_1[1]), .ZN(
        DataPath_Registers_Inst2_in2_1_) );
  XNOR2_X1 DataPath_Registers_Inst2_A2_U6 ( .A(
        DataPath_Registers_Inst2_reg_A_output2_1[5]), .B(
        DataPath_Registers_Inst2_reg_A_output2_1[4]), .ZN(
        DataPath_Registers_Inst2_A2_n10) );
  XNOR2_X1 DataPath_Registers_Inst2_A2_U5 ( .A(
        DataPath_Registers_Inst2_reg_A_output2_1[1]), .B(
        DataPath_Registers_Inst2_A2_n12), .ZN(DataPath_Registers_Inst2_in2_0_)
         );
  XNOR2_X1 DataPath_Registers_Inst2_A2_U4 ( .A(
        DataPath_Registers_Inst2_reg_A_output2_1[6]), .B(
        DataPath_Registers_Inst2_reg_A_output2_1[4]), .ZN(
        DataPath_Registers_Inst2_A2_n12) );
  XOR2_X1 DataPath_Registers_Inst2_A2_U3 ( .A(
        DataPath_Registers_Inst2_reg_A_output2_1[5]), .B(
        DataPath_Registers_Inst2_in2_6_), .Z(DataPath_Registers_Inst2_in2_4_)
         );
  XOR2_X1 DataPath_Registers_Inst2_A2_U2 ( .A(
        DataPath_Registers_Inst2_reg_A_output2_1[3]), .B(
        DataPath_Registers_Inst2_reg_A_output2_1[7]), .Z(
        DataPath_Registers_Inst2_in2_6_) );
  XOR2_X1 DataPath_Registers_Inst2_A2_U1 ( .A(
        DataPath_Registers_Inst2_reg_A_output2_1[5]), .B(
        DataPath_Registers_Inst2_reg_A_output2_1[3]), .Z(
        DataPath_Registers_Inst2_in2_7_) );
  XNOR2_X1 DataPath_Registers_Inst2_A3_U11 ( .A(
        DataPath_Registers_Inst2_in3_4_), .B(DataPath_Registers_Inst2_A3_n12), 
        .ZN(DataPath_Registers_Inst2_in3_3_) );
  XNOR2_X1 DataPath_Registers_Inst2_A3_U10 ( .A(
        DataPath_Registers_Inst2_A3_n11), .B(DataPath_Registers_Inst2_in3_5_), 
        .ZN(DataPath_Registers_Inst2_in3_2_) );
  XNOR2_X1 DataPath_Registers_Inst2_A3_U9 ( .A(DataPath_Registers_Inst2_in3_7_), .B(DataPath_Registers_Inst2_reg_A_output3_1[2]), .ZN(
        DataPath_Registers_Inst2_A3_n11) );
  XOR2_X1 DataPath_Registers_Inst2_A3_U8 ( .A(
        DataPath_Registers_Inst2_reg_A_output3_1[6]), .B(
        DataPath_Registers_Inst2_reg_A_output3_1[0]), .Z(
        DataPath_Registers_Inst2_in3_5_) );
  XNOR2_X1 DataPath_Registers_Inst2_A3_U7 ( .A(DataPath_Registers_Inst2_A3_n10), .B(DataPath_Registers_Inst2_reg_A_output3_1[1]), .ZN(
        DataPath_Registers_Inst2_in3_1_) );
  XNOR2_X1 DataPath_Registers_Inst2_A3_U6 ( .A(
        DataPath_Registers_Inst2_reg_A_output3_1[5]), .B(
        DataPath_Registers_Inst2_reg_A_output3_1[4]), .ZN(
        DataPath_Registers_Inst2_A3_n10) );
  XNOR2_X1 DataPath_Registers_Inst2_A3_U5 ( .A(
        DataPath_Registers_Inst2_reg_A_output3_1[1]), .B(
        DataPath_Registers_Inst2_A3_n12), .ZN(DataPath_Registers_Inst2_in3_0_)
         );
  XNOR2_X1 DataPath_Registers_Inst2_A3_U4 ( .A(
        DataPath_Registers_Inst2_reg_A_output3_1[6]), .B(
        DataPath_Registers_Inst2_reg_A_output3_1[4]), .ZN(
        DataPath_Registers_Inst2_A3_n12) );
  XOR2_X1 DataPath_Registers_Inst2_A3_U3 ( .A(
        DataPath_Registers_Inst2_reg_A_output3_1[5]), .B(
        DataPath_Registers_Inst2_in3_6_), .Z(DataPath_Registers_Inst2_in3_4_)
         );
  XOR2_X1 DataPath_Registers_Inst2_A3_U2 ( .A(
        DataPath_Registers_Inst2_reg_A_output3_1[3]), .B(
        DataPath_Registers_Inst2_reg_A_output3_1[7]), .Z(
        DataPath_Registers_Inst2_in3_6_) );
  XOR2_X1 DataPath_Registers_Inst2_A3_U1 ( .A(
        DataPath_Registers_Inst2_reg_A_output3_1[5]), .B(
        DataPath_Registers_Inst2_reg_A_output3_1[3]), .Z(
        DataPath_Registers_Inst2_in3_7_) );
  XNOR2_X1 DataPath_Registers_Inst2_A4_U11 ( .A(
        DataPath_Registers_Inst2_in4_4_), .B(DataPath_Registers_Inst2_A4_n12), 
        .ZN(DataPath_Registers_Inst2_in4_3_) );
  XNOR2_X1 DataPath_Registers_Inst2_A4_U10 ( .A(
        DataPath_Registers_Inst2_A4_n11), .B(DataPath_Registers_Inst2_in4_5_), 
        .ZN(DataPath_Registers_Inst2_in4_2_) );
  XNOR2_X1 DataPath_Registers_Inst2_A4_U9 ( .A(DataPath_Registers_Inst2_in4_7_), .B(DataPath_Registers_Inst2_reg_A_output4_1[2]), .ZN(
        DataPath_Registers_Inst2_A4_n11) );
  XOR2_X1 DataPath_Registers_Inst2_A4_U8 ( .A(
        DataPath_Registers_Inst2_reg_A_output4_1[6]), .B(
        DataPath_Registers_Inst2_reg_A_output4_1[0]), .Z(
        DataPath_Registers_Inst2_in4_5_) );
  XNOR2_X1 DataPath_Registers_Inst2_A4_U7 ( .A(DataPath_Registers_Inst2_A4_n10), .B(DataPath_Registers_Inst2_reg_A_output4_1[1]), .ZN(
        DataPath_Registers_Inst2_in4_1_) );
  XNOR2_X1 DataPath_Registers_Inst2_A4_U6 ( .A(
        DataPath_Registers_Inst2_reg_A_output4_1[5]), .B(
        DataPath_Registers_Inst2_reg_A_output4_1[4]), .ZN(
        DataPath_Registers_Inst2_A4_n10) );
  XNOR2_X1 DataPath_Registers_Inst2_A4_U5 ( .A(
        DataPath_Registers_Inst2_reg_A_output4_1[1]), .B(
        DataPath_Registers_Inst2_A4_n12), .ZN(DataPath_Registers_Inst2_in4_0_)
         );
  XNOR2_X1 DataPath_Registers_Inst2_A4_U4 ( .A(
        DataPath_Registers_Inst2_reg_A_output4_1[6]), .B(
        DataPath_Registers_Inst2_reg_A_output4_1[4]), .ZN(
        DataPath_Registers_Inst2_A4_n12) );
  XOR2_X1 DataPath_Registers_Inst2_A4_U3 ( .A(
        DataPath_Registers_Inst2_reg_A_output4_1[5]), .B(
        DataPath_Registers_Inst2_in4_6_), .Z(DataPath_Registers_Inst2_in4_4_)
         );
  XOR2_X1 DataPath_Registers_Inst2_A4_U2 ( .A(
        DataPath_Registers_Inst2_reg_A_output4_1[3]), .B(
        DataPath_Registers_Inst2_reg_A_output4_1[7]), .Z(
        DataPath_Registers_Inst2_in4_6_) );
  XOR2_X1 DataPath_Registers_Inst2_A4_U1 ( .A(
        DataPath_Registers_Inst2_reg_A_output4_1[5]), .B(
        DataPath_Registers_Inst2_reg_A_output4_1[3]), .Z(
        DataPath_Registers_Inst2_in4_7_) );
  AOI22_X1 Key_Registers_INST1_U124 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n282), .B1(Key_Registers_INST1_n130), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n226) );
  AOI22_X1 Key_Registers_INST1_U123 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n130), .B1(Key_Registers_INST1_n128), .B2(
        Key_Registers_INST1_n285), .ZN(Key_Registers_INST1_n225) );
  MUX2_X1 Key_Registers_INST1_U122 ( .A(Key_Registers_INST1_S14_in[0]), .B(
        Key_Registers_INST1_n249), .S(Key_Registers_INST1_n283), .Z(
        Key_Registers_INST1_n224) );
  MUX2_X1 Key_Registers_INST1_U121 ( .A(Key_Registers_INST1_S14_in[1]), .B(
        Key_Registers_INST1_n242), .S(Key_Registers_INST1_n283), .Z(
        Key_Registers_INST1_n223) );
  AOI22_X1 Key_Registers_INST1_U120 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n281), .B1(Key_Registers_INST1_n126), .B2(
        Key_Registers_INST1_n285), .ZN(Key_Registers_INST1_n222) );
  AOI22_X1 Key_Registers_INST1_U119 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n126), .B1(Key_Registers_INST1_n125), .B2(
        Key_Registers_INST1_n285), .ZN(Key_Registers_INST1_n221) );
  MUX2_X1 Key_Registers_INST1_U118 ( .A(Key_Registers_INST1_S14_in[2]), .B(
        Key_Registers_INST1_n241), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n220) );
  AOI22_X1 Key_Registers_INST1_U117 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n280), .B1(Key_Registers_INST1_n123), .B2(
        Key_Registers_INST1_n285), .ZN(Key_Registers_INST1_n219) );
  AOI22_X1 Key_Registers_INST1_U116 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n123), .B1(Key_Registers_INST1_n122), .B2(
        Key_Registers_INST1_n285), .ZN(Key_Registers_INST1_n218) );
  MUX2_X1 Key_Registers_INST1_U115 ( .A(Key_Registers_INST1_S14_in[3]), .B(
        Key_Registers_INST1_n240), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n217) );
  AOI22_X1 Key_Registers_INST1_U114 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n279), .B1(Key_Registers_INST1_n120), .B2(
        Key_Registers_INST1_n285), .ZN(Key_Registers_INST1_n216) );
  AOI22_X1 Key_Registers_INST1_U113 ( .A1(Key_Registers_INST1_n317), .A2(
        Key_Registers_INST1_n120), .B1(Key_Registers_INST1_n119), .B2(
        Key_Registers_INST1_n285), .ZN(Key_Registers_INST1_n215) );
  MUX2_X1 Key_Registers_INST1_U112 ( .A(Key_Registers_INST1_S14_in[4]), .B(
        Key_Registers_INST1_n239), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n214) );
  AOI22_X1 Key_Registers_INST1_U111 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n278), .B1(Key_Registers_INST1_n117), .B2(
        Key_Registers_INST1_n285), .ZN(Key_Registers_INST1_n213) );
  AOI22_X1 Key_Registers_INST1_U110 ( .A1(Key_Registers_INST1_n317), .A2(
        Key_Registers_INST1_n117), .B1(Key_Registers_INST1_n116), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n212) );
  MUX2_X1 Key_Registers_INST1_U109 ( .A(Key_Registers_INST1_S14_in[5]), .B(
        Key_Registers_INST1_n238), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n211) );
  AOI22_X1 Key_Registers_INST1_U108 ( .A1(Key_Registers_INST1_n317), .A2(
        Key_Registers_INST1_n277), .B1(Key_Registers_INST1_n114), .B2(
        Key_Registers_INST1_n285), .ZN(Key_Registers_INST1_n210) );
  AOI22_X1 Key_Registers_INST1_U107 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n114), .B1(Key_Registers_INST1_n113), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n209) );
  MUX2_X1 Key_Registers_INST1_U106 ( .A(Key_Registers_INST1_S14_in[6]), .B(
        Key_Registers_INST1_n237), .S(Key_Registers_INST1_n285), .Z(
        Key_Registers_INST1_n208) );
  AOI22_X1 Key_Registers_INST1_U105 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n276), .B1(Key_Registers_INST1_n111), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n207) );
  AOI22_X1 Key_Registers_INST1_U104 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n111), .B1(Key_Registers_INST1_n110), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n206) );
  MUX2_X1 Key_Registers_INST1_U103 ( .A(Key_Registers_INST1_S14_in[7]), .B(
        Key_Registers_INST1_n236), .S(Key_Registers_INST1_n285), .Z(
        Key_Registers_INST1_n205) );
  AOI22_X1 Key_Registers_INST1_U102 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n275), .B1(Key_Registers_INST1_n108), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n204) );
  AOI22_X1 Key_Registers_INST1_U101 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n108), .B1(Key_Registers_INST1_n107), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n203) );
  MUX2_X1 Key_Registers_INST1_U100 ( .A(Key_Registers_INST1_S10_in[0]), .B(
        Key_Registers_INST1_n235), .S(Key_Registers_INST1_n285), .Z(
        Key_Registers_INST1_n202) );
  INV_X1 Key_Registers_INST1_U99 ( .A(Key_Registers_INST1_n316), .ZN(
        Key_Registers_INST1_n201) );
  OAI22_X1 Key_Registers_INST1_U98 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n235), .B1(Key_Registers_INST1_n234), .B2(
        Key_Registers_INST1_n288), .ZN(Key_Registers_INST1_n316) );
  AOI22_X1 Key_Registers_INST1_U97 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n274), .B1(Key_Registers_INST1_n104), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n200) );
  MUX2_X1 Key_Registers_INST1_U96 ( .A(Key_Registers_INST1_S10_in[1]), .B(
        Key_Registers_INST1_n233), .S(Key_Registers_INST1_n285), .Z(
        Key_Registers_INST1_n199) );
  INV_X1 Key_Registers_INST1_U95 ( .A(Key_Registers_INST1_n315), .ZN(
        Key_Registers_INST1_n198) );
  OAI22_X1 Key_Registers_INST1_U94 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n233), .B1(Key_Registers_INST1_n232), .B2(
        Key_Registers_INST1_n317), .ZN(Key_Registers_INST1_n315) );
  AOI22_X1 Key_Registers_INST1_U93 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n273), .B1(Key_Registers_INST1_n101), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n197) );
  MUX2_X1 Key_Registers_INST1_U92 ( .A(Key_Registers_INST1_S10_in[2]), .B(
        Key_Registers_INST1_n231), .S(Key_Registers_INST1_n285), .Z(
        Key_Registers_INST1_n196) );
  INV_X1 Key_Registers_INST1_U91 ( .A(Key_Registers_INST1_n314), .ZN(
        Key_Registers_INST1_n195) );
  OAI22_X1 Key_Registers_INST1_U90 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n231), .B1(Key_Registers_INST1_n230), .B2(
        Key_Registers_INST1_n287), .ZN(Key_Registers_INST1_n314) );
  AOI22_X1 Key_Registers_INST1_U89 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n272), .B1(Key_Registers_INST1_n98), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n194) );
  MUX2_X1 Key_Registers_INST1_U88 ( .A(Key_Registers_INST1_S10_in[3]), .B(
        Key_Registers_INST1_n229), .S(Key_Registers_INST1_n285), .Z(
        Key_Registers_INST1_n193) );
  INV_X1 Key_Registers_INST1_U87 ( .A(Key_Registers_INST1_n313), .ZN(
        Key_Registers_INST1_n192) );
  OAI22_X1 Key_Registers_INST1_U86 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n229), .B1(Key_Registers_INST1_n228), .B2(
        Key_Registers_INST1_n288), .ZN(Key_Registers_INST1_n313) );
  AOI22_X1 Key_Registers_INST1_U85 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n271), .B1(Key_Registers_INST1_n95), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n191) );
  MUX2_X1 Key_Registers_INST1_U84 ( .A(Key_Registers_INST1_S10_in[4]), .B(
        Key_Registers_INST1_n227), .S(Key_Registers_INST1_n285), .Z(
        Key_Registers_INST1_n190) );
  INV_X1 Key_Registers_INST1_U83 ( .A(Key_Registers_INST1_n312), .ZN(
        Key_Registers_INST1_n189) );
  OAI22_X1 Key_Registers_INST1_U82 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n227), .B1(Key_Registers_INST1_n129), .B2(
        Key_Registers_INST1_n288), .ZN(Key_Registers_INST1_n312) );
  AOI22_X1 Key_Registers_INST1_U81 ( .A1(Key_Registers_INST1_n317), .A2(
        Key_Registers_INST1_n270), .B1(Key_Registers_INST1_n92), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n188) );
  MUX2_X1 Key_Registers_INST1_U80 ( .A(Key_Registers_INST1_S10_in[5]), .B(
        Key_Registers_INST1_n127), .S(Key_Registers_INST1_n285), .Z(
        Key_Registers_INST1_n187) );
  INV_X1 Key_Registers_INST1_U79 ( .A(Key_Registers_INST1_n311), .ZN(
        Key_Registers_INST1_n186) );
  OAI22_X1 Key_Registers_INST1_U78 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n127), .B1(Key_Registers_INST1_n124), .B2(
        Key_Registers_INST1_n317), .ZN(Key_Registers_INST1_n311) );
  AOI22_X1 Key_Registers_INST1_U77 ( .A1(Key_Registers_INST1_n317), .A2(
        Key_Registers_INST1_n269), .B1(Key_Registers_INST1_n89), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n185) );
  MUX2_X1 Key_Registers_INST1_U76 ( .A(Key_Registers_INST1_S10_in[6]), .B(
        Key_Registers_INST1_n121), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n184) );
  INV_X1 Key_Registers_INST1_U75 ( .A(Key_Registers_INST1_n310), .ZN(
        Key_Registers_INST1_n183) );
  OAI22_X1 Key_Registers_INST1_U74 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n121), .B1(Key_Registers_INST1_n118), .B2(
        Key_Registers_INST1_n317), .ZN(Key_Registers_INST1_n310) );
  AOI22_X1 Key_Registers_INST1_U73 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n268), .B1(Key_Registers_INST1_n86), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n182) );
  MUX2_X1 Key_Registers_INST1_U72 ( .A(Key_Registers_INST1_S10_in[7]), .B(
        Key_Registers_INST1_n115), .S(Key_Registers_INST1_n285), .Z(
        Key_Registers_INST1_n181) );
  INV_X1 Key_Registers_INST1_U71 ( .A(Key_Registers_INST1_n309), .ZN(
        Key_Registers_INST1_n180) );
  OAI22_X1 Key_Registers_INST1_U70 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n115), .B1(Key_Registers_INST1_n112), .B2(
        Key_Registers_INST1_n288), .ZN(Key_Registers_INST1_n309) );
  AOI22_X1 Key_Registers_INST1_U69 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n267), .B1(Key_Registers_INST1_n83), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n179) );
  MUX2_X1 Key_Registers_INST1_U68 ( .A(Key_Registers_INST1_S6_in[0]), .B(
        Key_Registers_INST1_n109), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n178) );
  INV_X1 Key_Registers_INST1_U67 ( .A(Key_Registers_INST1_n308), .ZN(
        Key_Registers_INST1_n177) );
  OAI22_X1 Key_Registers_INST1_U66 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n109), .B1(Key_Registers_INST1_n106), .B2(
        Key_Registers_INST1_n287), .ZN(Key_Registers_INST1_n308) );
  AOI22_X1 Key_Registers_INST1_U65 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n266), .B1(Key_Registers_INST1_n80), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n176) );
  MUX2_X1 Key_Registers_INST1_U64 ( .A(Key_Registers_INST1_S6_in[1]), .B(
        Key_Registers_INST1_n105), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n175) );
  INV_X1 Key_Registers_INST1_U63 ( .A(Key_Registers_INST1_n307), .ZN(
        Key_Registers_INST1_n174) );
  OAI22_X1 Key_Registers_INST1_U62 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n105), .B1(Key_Registers_INST1_n103), .B2(
        Key_Registers_INST1_n287), .ZN(Key_Registers_INST1_n307) );
  AOI22_X1 Key_Registers_INST1_U61 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n265), .B1(Key_Registers_INST1_n77), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n173) );
  MUX2_X1 Key_Registers_INST1_U60 ( .A(Key_Registers_INST1_S6_in[2]), .B(
        Key_Registers_INST1_n102), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n172) );
  INV_X1 Key_Registers_INST1_U59 ( .A(Key_Registers_INST1_n306), .ZN(
        Key_Registers_INST1_n171) );
  OAI22_X1 Key_Registers_INST1_U58 ( .A1(Key_Registers_INST1_n284), .A2(
        Key_Registers_INST1_n102), .B1(Key_Registers_INST1_n100), .B2(
        Key_Registers_INST1_n317), .ZN(Key_Registers_INST1_n306) );
  AOI22_X1 Key_Registers_INST1_U57 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n264), .B1(Key_Registers_INST1_n74), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n170) );
  MUX2_X1 Key_Registers_INST1_U56 ( .A(Key_Registers_INST1_S6_in[3]), .B(
        Key_Registers_INST1_n99), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n169) );
  INV_X1 Key_Registers_INST1_U55 ( .A(Key_Registers_INST1_n305), .ZN(
        Key_Registers_INST1_n168) );
  OAI22_X1 Key_Registers_INST1_U54 ( .A1(Key_Registers_INST1_n286), .A2(
        Key_Registers_INST1_n99), .B1(Key_Registers_INST1_n97), .B2(
        Key_Registers_INST1_n288), .ZN(Key_Registers_INST1_n305) );
  AOI22_X1 Key_Registers_INST1_U53 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n263), .B1(Key_Registers_INST1_n71), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n167) );
  MUX2_X1 Key_Registers_INST1_U52 ( .A(Key_Registers_INST1_S6_in[4]), .B(
        Key_Registers_INST1_n96), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n166) );
  INV_X1 Key_Registers_INST1_U51 ( .A(Key_Registers_INST1_n304), .ZN(
        Key_Registers_INST1_n165) );
  OAI22_X1 Key_Registers_INST1_U50 ( .A1(Key_Registers_INST1_n285), .A2(
        Key_Registers_INST1_n96), .B1(Key_Registers_INST1_n94), .B2(
        Key_Registers_INST1_n287), .ZN(Key_Registers_INST1_n304) );
  AOI22_X1 Key_Registers_INST1_U49 ( .A1(Key_Registers_INST1_n287), .A2(
        Key_Registers_INST1_n262), .B1(Key_Registers_INST1_n68), .B2(
        Key_Registers_INST1_n286), .ZN(Key_Registers_INST1_n164) );
  MUX2_X1 Key_Registers_INST1_U48 ( .A(Key_Registers_INST1_S6_in[5]), .B(
        Key_Registers_INST1_n79), .S(Key_Registers_INST1_n284), .Z(
        Key_Registers_INST1_n163) );
  INV_X1 Key_Registers_INST1_U47 ( .A(Key_Registers_INST1_n303), .ZN(
        Key_Registers_INST1_n162) );
  OAI22_X1 Key_Registers_INST1_U46 ( .A1(Key_Registers_INST1_n286), .A2(
        Key_Registers_INST1_n79), .B1(Key_Registers_INST1_n78), .B2(
        Key_Registers_INST1_n287), .ZN(Key_Registers_INST1_n303) );
  AOI22_X1 Key_Registers_INST1_U45 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n261), .B1(Key_Registers_INST1_n65), .B2(
        Key_Registers_INST1_n284), .ZN(Key_Registers_INST1_n161) );
  MUX2_X1 Key_Registers_INST1_U44 ( .A(Key_Registers_INST1_S6_in[6]), .B(
        Key_Registers_INST1_n76), .S(Key_Registers_INST1_n283), .Z(
        Key_Registers_INST1_n160) );
  INV_X1 Key_Registers_INST1_U43 ( .A(Key_Registers_INST1_n302), .ZN(
        Key_Registers_INST1_n159) );
  OAI22_X1 Key_Registers_INST1_U42 ( .A1(Key_Registers_INST1_n285), .A2(
        Key_Registers_INST1_n76), .B1(Key_Registers_INST1_n75), .B2(
        Key_Registers_INST1_n288), .ZN(Key_Registers_INST1_n302) );
  AOI22_X1 Key_Registers_INST1_U41 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n260), .B1(Key_Registers_INST1_n62), .B2(
        Key_Registers_INST1_n284), .ZN(Key_Registers_INST1_n158) );
  MUX2_X1 Key_Registers_INST1_U40 ( .A(Key_Registers_INST1_S6_in[7]), .B(
        Key_Registers_INST1_n73), .S(Key_Registers_INST1_n283), .Z(
        Key_Registers_INST1_n157) );
  INV_X1 Key_Registers_INST1_U39 ( .A(Key_Registers_INST1_n301), .ZN(
        Key_Registers_INST1_n156) );
  OAI22_X1 Key_Registers_INST1_U38 ( .A1(Key_Registers_INST1_n286), .A2(
        Key_Registers_INST1_n73), .B1(Key_Registers_INST1_n72), .B2(
        Key_Registers_INST1_n288), .ZN(Key_Registers_INST1_n301) );
  AOI22_X1 Key_Registers_INST1_U37 ( .A1(Key_Registers_INST1_n288), .A2(
        Key_Registers_INST1_n259), .B1(Key_Registers_INST1_n59), .B2(
        Key_Registers_INST1_n285), .ZN(Key_Registers_INST1_n155) );
  MUX2_X1 Key_Registers_INST1_U36 ( .A(Key_Registers_INST1_S2_in[0]), .B(
        Key_Registers_INST1_n93), .S(Key_Registers_INST1_n292), .Z(
        Key_Registers_INST1_n154) );
  OAI22_X1 Key_Registers_INST1_U35 ( .A1(Key_Registers_INST1_n292), .A2(
        Key_Registers_INST1_n93), .B1(Key_Registers_INST1_n91), .B2(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_n300) );
  AOI22_X1 Key_Registers_INST1_U34 ( .A1(Key_Registers_INST1_n290), .A2(
        Key_Registers_INST1_n258), .B1(Key_Registers_INST1_n56), .B2(
        Key_Registers_INST1_n292), .ZN(Key_Registers_INST1_n152) );
  MUX2_X1 Key_Registers_INST1_U33 ( .A(Key_Registers_INST1_S2_in[1]), .B(
        Key_Registers_INST1_n90), .S(Key_Registers_INST1_n292), .Z(
        Key_Registers_INST1_n151) );
  OAI22_X1 Key_Registers_INST1_U32 ( .A1(Key_Registers_INST1_n292), .A2(
        Key_Registers_INST1_n90), .B1(Key_Registers_INST1_n88), .B2(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_n299) );
  AOI22_X1 Key_Registers_INST1_U31 ( .A1(Key_Registers_INST1_n290), .A2(
        Key_Registers_INST1_n257), .B1(Key_Registers_INST1_n53), .B2(
        Key_Registers_INST1_n292), .ZN(Key_Registers_INST1_n149) );
  MUX2_X1 Key_Registers_INST1_U30 ( .A(Key_Registers_INST1_S2_in[2]), .B(
        Key_Registers_INST1_n87), .S(Key_Registers_INST1_n292), .Z(
        Key_Registers_INST1_n148) );
  OAI22_X1 Key_Registers_INST1_U29 ( .A1(Key_Registers_INST1_n292), .A2(
        Key_Registers_INST1_n87), .B1(Key_Registers_INST1_n85), .B2(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_n298) );
  AOI22_X1 Key_Registers_INST1_U28 ( .A1(Key_Registers_INST1_n290), .A2(
        Key_Registers_INST1_n256), .B1(Key_Registers_INST1_n50), .B2(
        Key_Registers_INST1_n291), .ZN(Key_Registers_INST1_n146) );
  MUX2_X1 Key_Registers_INST1_U27 ( .A(Key_Registers_INST1_S2_in[3]), .B(
        Key_Registers_INST1_n84), .S(Key_Registers_INST1_n292), .Z(
        Key_Registers_INST1_n145) );
  OAI22_X1 Key_Registers_INST1_U26 ( .A1(Key_Registers_INST1_n292), .A2(
        Key_Registers_INST1_n84), .B1(Key_Registers_INST1_n82), .B2(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_n297) );
  AOI22_X1 Key_Registers_INST1_U25 ( .A1(Key_Registers_INST1_n290), .A2(
        Key_Registers_INST1_n255), .B1(Key_Registers_INST1_n47), .B2(
        Key_Registers_INST1_n291), .ZN(Key_Registers_INST1_n143) );
  MUX2_X1 Key_Registers_INST1_U24 ( .A(Key_Registers_INST1_S2_in[4]), .B(
        Key_Registers_INST1_n250), .S(Key_Registers_INST1_n292), .Z(
        Key_Registers_INST1_n142) );
  OAI22_X1 Key_Registers_INST1_U23 ( .A1(Key_Registers_INST1_n292), .A2(
        Key_Registers_INST1_n250), .B1(Key_Registers_INST1_n248), .B2(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_n296) );
  AOI22_X1 Key_Registers_INST1_U22 ( .A1(Key_Registers_INST1_n290), .A2(
        Key_Registers_INST1_n254), .B1(Key_Registers_INST1_n44), .B2(
        Key_Registers_INST1_n291), .ZN(Key_Registers_INST1_n140) );
  MUX2_X1 Key_Registers_INST1_U21 ( .A(Key_Registers_INST1_S2_in[5]), .B(
        Key_Registers_INST1_n81), .S(Key_Registers_INST1_n292), .Z(
        Key_Registers_INST1_n139) );
  OAI22_X1 Key_Registers_INST1_U20 ( .A1(Key_Registers_INST1_n292), .A2(
        Key_Registers_INST1_n81), .B1(Key_Registers_INST1_n247), .B2(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_n295) );
  AOI22_X1 Key_Registers_INST1_U19 ( .A1(Key_Registers_INST1_n290), .A2(
        Key_Registers_INST1_n253), .B1(Key_Registers_INST1_n41), .B2(
        Key_Registers_INST1_n291), .ZN(Key_Registers_INST1_n137) );
  MUX2_X1 Key_Registers_INST1_U18 ( .A(Key_Registers_INST1_S2_in[6]), .B(
        Key_Registers_INST1_n246), .S(Key_Registers_INST1_n292), .Z(
        Key_Registers_INST1_n136) );
  OAI22_X1 Key_Registers_INST1_U17 ( .A1(Key_Registers_INST1_n292), .A2(
        Key_Registers_INST1_n246), .B1(Key_Registers_INST1_n245), .B2(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_n294) );
  AOI22_X1 Key_Registers_INST1_U16 ( .A1(Key_Registers_INST1_n290), .A2(
        Key_Registers_INST1_n252), .B1(Key_Registers_INST1_n38), .B2(
        Key_Registers_INST1_n292), .ZN(Key_Registers_INST1_n134) );
  MUX2_X1 Key_Registers_INST1_U15 ( .A(Key_Registers_INST1_S2_in[7]), .B(
        Key_Registers_INST1_n244), .S(Key_Registers_INST1_n292), .Z(
        Key_Registers_INST1_n133) );
  OAI22_X1 Key_Registers_INST1_U14 ( .A1(Key_Registers_INST1_n292), .A2(
        Key_Registers_INST1_n244), .B1(Key_Registers_INST1_n243), .B2(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_n293) );
  AOI22_X1 Key_Registers_INST1_U13 ( .A1(Key_Registers_INST1_n290), .A2(
        Key_Registers_INST1_n251), .B1(Key_Registers_INST1_n35), .B2(
        Key_Registers_INST1_n292), .ZN(Key_Registers_INST1_n131) );
  BUF_X2 Key_Registers_INST1_U12 ( .A(DoKeySbox), .Z(Key_Registers_INST1_n289)
         );
  INV_X2 Key_Registers_INST1_U11 ( .A(Key_Registers_INST1_n291), .ZN(
        Key_Registers_INST1_n290) );
  INV_X2 Key_Registers_INST1_U10 ( .A(Key_Registers_INST1_n288), .ZN(
        Key_Registers_INST1_n284) );
  INV_X1 Key_Registers_INST1_U9 ( .A(key_reg_hold), .ZN(
        Key_Registers_INST1_n292) );
  BUF_X1 Key_Registers_INST1_U8 ( .A(Key_Registers_INST1_n292), .Z(
        Key_Registers_INST1_n291) );
  NOR2_X1 Key_Registers_INST1_U7 ( .A1(JustFirstColShift), .A2(
        Key_Registers_INST1_n291), .ZN(Key_Registers_INST1_n317) );
  BUF_X1 Key_Registers_INST1_U6 ( .A(Key_Registers_INST1_n317), .Z(
        Key_Registers_INST1_n287) );
  INV_X1 Key_Registers_INST1_U5 ( .A(Key_Registers_INST1_n287), .ZN(
        Key_Registers_INST1_n285) );
  BUF_X1 Key_Registers_INST1_U4 ( .A(Key_Registers_INST1_n317), .Z(
        Key_Registers_INST1_n288) );
  INV_X1 Key_Registers_INST1_U3 ( .A(Key_Registers_INST1_n288), .ZN(
        Key_Registers_INST1_n283) );
  INV_X1 Key_Registers_INST1_U2 ( .A(Key_Registers_INST1_n287), .ZN(
        Key_Registers_INST1_n286) );
  DFF_X1 Key_Registers_INST1_S1_reg_0_ ( .D(Key_Registers_INST1_n300), .CK(clk), .Q(Key_Registers_INST1_n258), .QN(Key_Registers_INST1_n91) );
  DFF_X1 Key_Registers_INST1_S1_reg_1_ ( .D(Key_Registers_INST1_n299), .CK(clk), .Q(Key_Registers_INST1_n257), .QN(Key_Registers_INST1_n88) );
  DFF_X1 Key_Registers_INST1_S1_reg_2_ ( .D(Key_Registers_INST1_n298), .CK(clk), .Q(Key_Registers_INST1_n256), .QN(Key_Registers_INST1_n85) );
  DFF_X1 Key_Registers_INST1_S1_reg_3_ ( .D(Key_Registers_INST1_n297), .CK(clk), .Q(Key_Registers_INST1_n255), .QN(Key_Registers_INST1_n82) );
  DFF_X1 Key_Registers_INST1_S1_reg_4_ ( .D(Key_Registers_INST1_n296), .CK(clk), .Q(Key_Registers_INST1_n254), .QN(Key_Registers_INST1_n248) );
  DFF_X1 Key_Registers_INST1_S1_reg_5_ ( .D(Key_Registers_INST1_n295), .CK(clk), .Q(Key_Registers_INST1_n253), .QN(Key_Registers_INST1_n247) );
  DFF_X1 Key_Registers_INST1_S1_reg_6_ ( .D(Key_Registers_INST1_n294), .CK(clk), .Q(Key_Registers_INST1_n252), .QN(Key_Registers_INST1_n245) );
  DFF_X1 Key_Registers_INST1_S1_reg_7_ ( .D(Key_Registers_INST1_n293), .CK(clk), .Q(Key_Registers_INST1_n251), .QN(Key_Registers_INST1_n243) );
  DFF_X1 Key_Registers_INST1_S0_reg_0_ ( .D(Key_Registers_INST1_n152), .CK(clk), .Q(KeyOut1[0]), .QN(Key_Registers_INST1_n56) );
  DFF_X1 Key_Registers_INST1_S0_reg_1_ ( .D(Key_Registers_INST1_n149), .CK(clk), .Q(KeyOut1[1]), .QN(Key_Registers_INST1_n53) );
  DFF_X1 Key_Registers_INST1_S0_reg_6_ ( .D(Key_Registers_INST1_n134), .CK(clk), .Q(KeyOut1[6]), .QN(Key_Registers_INST1_n38) );
  DFF_X1 Key_Registers_INST1_S0_reg_7_ ( .D(Key_Registers_INST1_n131), .CK(clk), .Q(KeyOut1[7]), .QN(Key_Registers_INST1_n35) );
  DFF_X1 Key_Registers_INST1_S0_reg_2_ ( .D(Key_Registers_INST1_n146), .CK(clk), .Q(KeyOut1[2]), .QN(Key_Registers_INST1_n50) );
  DFF_X1 Key_Registers_INST1_S0_reg_3_ ( .D(Key_Registers_INST1_n143), .CK(clk), .Q(KeyOut1[3]), .QN(Key_Registers_INST1_n47) );
  DFF_X1 Key_Registers_INST1_S0_reg_4_ ( .D(Key_Registers_INST1_n140), .CK(clk), .Q(KeyOut1[4]), .QN(Key_Registers_INST1_n44) );
  DFF_X1 Key_Registers_INST1_S0_reg_5_ ( .D(Key_Registers_INST1_n137), .CK(clk), .Q(KeyOut1[5]), .QN(Key_Registers_INST1_n41) );
  DFF_X1 Key_Registers_INST1_S13_reg_1_ ( .D(Key_Registers_INST1_n222), .CK(
        clk), .Q(KeyToSbox1[1]), .QN(Key_Registers_INST1_n126) );
  DFF_X1 Key_Registers_INST1_S13_reg_2_ ( .D(Key_Registers_INST1_n219), .CK(
        clk), .Q(KeyToSbox1[2]), .QN(Key_Registers_INST1_n123) );
  DFF_X1 Key_Registers_INST1_S13_reg_3_ ( .D(Key_Registers_INST1_n216), .CK(
        clk), .Q(KeyToSbox1[3]), .QN(Key_Registers_INST1_n120) );
  DFF_X1 Key_Registers_INST1_S13_reg_4_ ( .D(Key_Registers_INST1_n213), .CK(
        clk), .Q(KeyToSbox1[4]), .QN(Key_Registers_INST1_n117) );
  DFF_X1 Key_Registers_INST1_S13_reg_5_ ( .D(Key_Registers_INST1_n210), .CK(
        clk), .Q(KeyToSbox1[5]), .QN(Key_Registers_INST1_n114) );
  DFF_X1 Key_Registers_INST1_S13_reg_6_ ( .D(Key_Registers_INST1_n207), .CK(
        clk), .Q(KeyToSbox1[6]), .QN(Key_Registers_INST1_n111) );
  DFF_X1 Key_Registers_INST1_S13_reg_7_ ( .D(Key_Registers_INST1_n204), .CK(
        clk), .Q(KeyToSbox1[7]), .QN(Key_Registers_INST1_n108) );
  DFF_X1 Key_Registers_INST1_S12_reg_0_ ( .D(Key_Registers_INST1_n225), .CK(
        clk), .Q(KeyForSchedule1[0]), .QN(Key_Registers_INST1_n128) );
  DFF_X1 Key_Registers_INST1_S13_reg_0_ ( .D(Key_Registers_INST1_n226), .CK(
        clk), .Q(KeyToSbox1[0]), .QN(Key_Registers_INST1_n130) );
  DFF_X1 Key_Registers_INST1_S5_reg_7_ ( .D(Key_Registers_INST1_n156), .CK(clk), .Q(Key_Registers_INST1_n72), .QN(Key_Registers_INST1_n259) );
  DFF_X1 Key_Registers_INST1_S6_reg_7_ ( .D(Key_Registers_INST1_n157), .CK(clk), .Q(Key_Registers_INST1_n73), .QN() );
  DFF_X1 Key_Registers_INST1_S5_reg_5_ ( .D(Key_Registers_INST1_n162), .CK(clk), .Q(Key_Registers_INST1_n78), .QN(Key_Registers_INST1_n261) );
  DFF_X1 Key_Registers_INST1_S5_reg_6_ ( .D(Key_Registers_INST1_n159), .CK(clk), .Q(Key_Registers_INST1_n75), .QN(Key_Registers_INST1_n260) );
  DFF_X1 Key_Registers_INST1_S6_reg_5_ ( .D(Key_Registers_INST1_n163), .CK(clk), .Q(Key_Registers_INST1_n79), .QN() );
  DFF_X1 Key_Registers_INST1_S6_reg_6_ ( .D(Key_Registers_INST1_n160), .CK(clk), .Q(Key_Registers_INST1_n76), .QN() );
  DFF_X1 Key_Registers_INST1_S5_reg_0_ ( .D(Key_Registers_INST1_n177), .CK(clk), .Q(Key_Registers_INST1_n106), .QN(Key_Registers_INST1_n266) );
  DFF_X1 Key_Registers_INST1_S5_reg_1_ ( .D(Key_Registers_INST1_n174), .CK(clk), .Q(Key_Registers_INST1_n103), .QN(Key_Registers_INST1_n265) );
  DFF_X1 Key_Registers_INST1_S5_reg_2_ ( .D(Key_Registers_INST1_n171), .CK(clk), .Q(Key_Registers_INST1_n100), .QN(Key_Registers_INST1_n264) );
  DFF_X1 Key_Registers_INST1_S5_reg_3_ ( .D(Key_Registers_INST1_n168), .CK(clk), .Q(Key_Registers_INST1_n97), .QN(Key_Registers_INST1_n263) );
  DFF_X1 Key_Registers_INST1_S5_reg_4_ ( .D(Key_Registers_INST1_n165), .CK(clk), .Q(Key_Registers_INST1_n94), .QN(Key_Registers_INST1_n262) );
  DFF_X1 Key_Registers_INST1_S6_reg_0_ ( .D(Key_Registers_INST1_n178), .CK(clk), .Q(Key_Registers_INST1_n109), .QN() );
  DFF_X1 Key_Registers_INST1_S6_reg_1_ ( .D(Key_Registers_INST1_n175), .CK(clk), .Q(Key_Registers_INST1_n105), .QN() );
  DFF_X1 Key_Registers_INST1_S6_reg_2_ ( .D(Key_Registers_INST1_n172), .CK(clk), .Q(Key_Registers_INST1_n102), .QN() );
  DFF_X1 Key_Registers_INST1_S6_reg_3_ ( .D(Key_Registers_INST1_n169), .CK(clk), .Q(Key_Registers_INST1_n99), .QN() );
  DFF_X1 Key_Registers_INST1_S6_reg_4_ ( .D(Key_Registers_INST1_n166), .CK(clk), .Q(Key_Registers_INST1_n96), .QN() );
  DFF_X1 Key_Registers_INST1_S9_reg_0_ ( .D(Key_Registers_INST1_n201), .CK(clk), .Q(Key_Registers_INST1_n234), .QN(Key_Registers_INST1_n274) );
  DFF_X1 Key_Registers_INST1_S9_reg_1_ ( .D(Key_Registers_INST1_n198), .CK(clk), .Q(Key_Registers_INST1_n232), .QN(Key_Registers_INST1_n273) );
  DFF_X1 Key_Registers_INST1_S9_reg_2_ ( .D(Key_Registers_INST1_n195), .CK(clk), .Q(Key_Registers_INST1_n230), .QN(Key_Registers_INST1_n272) );
  DFF_X1 Key_Registers_INST1_S9_reg_3_ ( .D(Key_Registers_INST1_n192), .CK(clk), .Q(Key_Registers_INST1_n228), .QN(Key_Registers_INST1_n271) );
  DFF_X1 Key_Registers_INST1_S9_reg_4_ ( .D(Key_Registers_INST1_n189), .CK(clk), .Q(Key_Registers_INST1_n129), .QN(Key_Registers_INST1_n270) );
  DFF_X1 Key_Registers_INST1_S9_reg_5_ ( .D(Key_Registers_INST1_n186), .CK(clk), .Q(Key_Registers_INST1_n124), .QN(Key_Registers_INST1_n269) );
  DFF_X1 Key_Registers_INST1_S9_reg_6_ ( .D(Key_Registers_INST1_n183), .CK(clk), .Q(Key_Registers_INST1_n118), .QN(Key_Registers_INST1_n268) );
  DFF_X1 Key_Registers_INST1_S9_reg_7_ ( .D(Key_Registers_INST1_n180), .CK(clk), .Q(Key_Registers_INST1_n112), .QN(Key_Registers_INST1_n267) );
  DFF_X1 Key_Registers_INST1_S10_reg_0_ ( .D(Key_Registers_INST1_n202), .CK(
        clk), .Q(Key_Registers_INST1_n235), .QN() );
  DFF_X1 Key_Registers_INST1_S10_reg_1_ ( .D(Key_Registers_INST1_n199), .CK(
        clk), .Q(Key_Registers_INST1_n233), .QN() );
  DFF_X1 Key_Registers_INST1_S10_reg_2_ ( .D(Key_Registers_INST1_n196), .CK(
        clk), .Q(Key_Registers_INST1_n231), .QN() );
  DFF_X1 Key_Registers_INST1_S10_reg_3_ ( .D(Key_Registers_INST1_n193), .CK(
        clk), .Q(Key_Registers_INST1_n229), .QN() );
  DFF_X1 Key_Registers_INST1_S10_reg_4_ ( .D(Key_Registers_INST1_n190), .CK(
        clk), .Q(Key_Registers_INST1_n227), .QN() );
  DFF_X1 Key_Registers_INST1_S10_reg_5_ ( .D(Key_Registers_INST1_n187), .CK(
        clk), .Q(Key_Registers_INST1_n127), .QN() );
  DFF_X1 Key_Registers_INST1_S10_reg_6_ ( .D(Key_Registers_INST1_n184), .CK(
        clk), .Q(Key_Registers_INST1_n121), .QN() );
  DFF_X1 Key_Registers_INST1_S10_reg_7_ ( .D(Key_Registers_INST1_n181), .CK(
        clk), .Q(Key_Registers_INST1_n115), .QN() );
  DFF_X1 Key_Registers_INST1_S14_reg_0_ ( .D(Key_Registers_INST1_n224), .CK(
        clk), .Q(Key_Registers_INST1_n249), .QN(Key_Registers_INST1_n282) );
  DFF_X1 Key_Registers_INST1_S14_reg_1_ ( .D(Key_Registers_INST1_n223), .CK(
        clk), .Q(Key_Registers_INST1_n242), .QN(Key_Registers_INST1_n281) );
  DFF_X1 Key_Registers_INST1_S14_reg_2_ ( .D(Key_Registers_INST1_n220), .CK(
        clk), .Q(Key_Registers_INST1_n241), .QN(Key_Registers_INST1_n280) );
  DFF_X1 Key_Registers_INST1_S14_reg_3_ ( .D(Key_Registers_INST1_n217), .CK(
        clk), .Q(Key_Registers_INST1_n240), .QN(Key_Registers_INST1_n279) );
  DFF_X1 Key_Registers_INST1_S14_reg_4_ ( .D(Key_Registers_INST1_n214), .CK(
        clk), .Q(Key_Registers_INST1_n239), .QN(Key_Registers_INST1_n278) );
  DFF_X1 Key_Registers_INST1_S14_reg_5_ ( .D(Key_Registers_INST1_n211), .CK(
        clk), .Q(Key_Registers_INST1_n238), .QN(Key_Registers_INST1_n277) );
  DFF_X1 Key_Registers_INST1_S14_reg_6_ ( .D(Key_Registers_INST1_n208), .CK(
        clk), .Q(Key_Registers_INST1_n237), .QN(Key_Registers_INST1_n276) );
  DFF_X1 Key_Registers_INST1_S14_reg_7_ ( .D(Key_Registers_INST1_n205), .CK(
        clk), .Q(Key_Registers_INST1_n236), .QN(Key_Registers_INST1_n275) );
  DFF_X1 Key_Registers_INST1_S2_reg_0_ ( .D(Key_Registers_INST1_n154), .CK(clk), .Q(Key_Registers_INST1_n93), .QN() );
  DFF_X1 Key_Registers_INST1_S2_reg_1_ ( .D(Key_Registers_INST1_n151), .CK(clk), .Q(Key_Registers_INST1_n90), .QN() );
  DFF_X1 Key_Registers_INST1_S2_reg_2_ ( .D(Key_Registers_INST1_n148), .CK(clk), .Q(Key_Registers_INST1_n87), .QN() );
  DFF_X1 Key_Registers_INST1_S2_reg_3_ ( .D(Key_Registers_INST1_n145), .CK(clk), .Q(Key_Registers_INST1_n84), .QN() );
  DFF_X1 Key_Registers_INST1_S2_reg_5_ ( .D(Key_Registers_INST1_n139), .CK(clk), .Q(Key_Registers_INST1_n81), .QN() );
  DFF_X1 Key_Registers_INST1_S2_reg_6_ ( .D(Key_Registers_INST1_n136), .CK(clk), .Q(Key_Registers_INST1_n246), .QN() );
  DFF_X1 Key_Registers_INST1_S2_reg_7_ ( .D(Key_Registers_INST1_n133), .CK(clk), .Q(Key_Registers_INST1_n244), .QN() );
  DFF_X1 Key_Registers_INST1_S2_reg_4_ ( .D(Key_Registers_INST1_n142), .CK(clk), .Q(Key_Registers_INST1_n250), .QN() );
  DFF_X1 Key_Registers_INST1_S4_reg_7_ ( .D(Key_Registers_INST1_n155), .CK(clk), .Q(Key_Registers_INST1_S4_7_), .QN(Key_Registers_INST1_n59) );
  DFF_X1 Key_Registers_INST1_S4_reg_6_ ( .D(Key_Registers_INST1_n158), .CK(clk), .Q(Key_Registers_INST1_S4_6_), .QN(Key_Registers_INST1_n62) );
  DFF_X1 Key_Registers_INST1_S4_reg_5_ ( .D(Key_Registers_INST1_n161), .CK(clk), .Q(Key_Registers_INST1_S4_5_), .QN(Key_Registers_INST1_n65) );
  DFF_X1 Key_Registers_INST1_S4_reg_4_ ( .D(Key_Registers_INST1_n164), .CK(clk), .Q(Key_Registers_INST1_S4_4_), .QN(Key_Registers_INST1_n68) );
  DFF_X1 Key_Registers_INST1_S4_reg_3_ ( .D(Key_Registers_INST1_n167), .CK(clk), .Q(Key_Registers_INST1_S4_3_), .QN(Key_Registers_INST1_n71) );
  DFF_X1 Key_Registers_INST1_S4_reg_2_ ( .D(Key_Registers_INST1_n170), .CK(clk), .Q(Key_Registers_INST1_S4_2_), .QN(Key_Registers_INST1_n74) );
  DFF_X1 Key_Registers_INST1_S4_reg_1_ ( .D(Key_Registers_INST1_n173), .CK(clk), .Q(Key_Registers_INST1_S4_1_), .QN(Key_Registers_INST1_n77) );
  DFF_X1 Key_Registers_INST1_S4_reg_0_ ( .D(Key_Registers_INST1_n176), .CK(clk), .Q(Key_Registers_INST1_S4_0_), .QN(Key_Registers_INST1_n80) );
  DFF_X1 Key_Registers_INST1_S8_reg_7_ ( .D(Key_Registers_INST1_n179), .CK(clk), .Q(Key_Registers_INST1_S8_7_), .QN(Key_Registers_INST1_n83) );
  DFF_X1 Key_Registers_INST1_S8_reg_6_ ( .D(Key_Registers_INST1_n182), .CK(clk), .Q(Key_Registers_INST1_S8_6_), .QN(Key_Registers_INST1_n86) );
  DFF_X1 Key_Registers_INST1_S8_reg_5_ ( .D(Key_Registers_INST1_n185), .CK(clk), .Q(Key_Registers_INST1_S8_5_), .QN(Key_Registers_INST1_n89) );
  DFF_X1 Key_Registers_INST1_S8_reg_4_ ( .D(Key_Registers_INST1_n188), .CK(clk), .Q(Key_Registers_INST1_S8_4_), .QN(Key_Registers_INST1_n92) );
  DFF_X1 Key_Registers_INST1_S8_reg_3_ ( .D(Key_Registers_INST1_n191), .CK(clk), .Q(Key_Registers_INST1_S8_3_), .QN(Key_Registers_INST1_n95) );
  DFF_X1 Key_Registers_INST1_S8_reg_2_ ( .D(Key_Registers_INST1_n194), .CK(clk), .Q(Key_Registers_INST1_S8_2_), .QN(Key_Registers_INST1_n98) );
  DFF_X1 Key_Registers_INST1_S8_reg_1_ ( .D(Key_Registers_INST1_n197), .CK(clk), .Q(Key_Registers_INST1_S8_1_), .QN(Key_Registers_INST1_n101) );
  DFF_X1 Key_Registers_INST1_S8_reg_0_ ( .D(Key_Registers_INST1_n200), .CK(clk), .Q(Key_Registers_INST1_S8_0_), .QN(Key_Registers_INST1_n104) );
  DFF_X1 Key_Registers_INST1_S12_reg_7_ ( .D(Key_Registers_INST1_n203), .CK(
        clk), .Q(KeyForSchedule1[7]), .QN(Key_Registers_INST1_n107) );
  DFF_X1 Key_Registers_INST1_S12_reg_6_ ( .D(Key_Registers_INST1_n206), .CK(
        clk), .Q(KeyForSchedule1[6]), .QN(Key_Registers_INST1_n110) );
  DFF_X1 Key_Registers_INST1_S12_reg_5_ ( .D(Key_Registers_INST1_n209), .CK(
        clk), .Q(KeyForSchedule1[5]), .QN(Key_Registers_INST1_n113) );
  DFF_X1 Key_Registers_INST1_S12_reg_4_ ( .D(Key_Registers_INST1_n212), .CK(
        clk), .Q(KeyForSchedule1[4]), .QN(Key_Registers_INST1_n116) );
  DFF_X1 Key_Registers_INST1_S12_reg_3_ ( .D(Key_Registers_INST1_n215), .CK(
        clk), .Q(KeyForSchedule1[3]), .QN(Key_Registers_INST1_n119) );
  DFF_X1 Key_Registers_INST1_S12_reg_2_ ( .D(Key_Registers_INST1_n218), .CK(
        clk), .Q(KeyForSchedule1[2]), .QN(Key_Registers_INST1_n122) );
  DFF_X1 Key_Registers_INST1_S12_reg_1_ ( .D(Key_Registers_INST1_n221), .CK(
        clk), .Q(KeyForSchedule1[1]), .QN(Key_Registers_INST1_n125) );
  OAI21_X1 Key_Registers_INST1_ScanFF_S3_SFF_0_U4 ( .B1(
        Key_Registers_INST1_n290), .B2(Key_Registers_INST1_ScanFF_S3_SFF_0_n8), 
        .A(Key_Registers_INST1_ScanFF_S3_SFF_0_n11), .ZN(
        Key_Registers_INST1_ScanFF_S3_SFF_0_n7) );
  OAI221_X1 Key_Registers_INST1_ScanFF_S3_SFF_0_U3 ( .B1(
        Key_Registers_INST1_n289), .B2(Key_Registers_INST1_S4_0_), .C1(
        Key_Registers_INST1_ScanFF_S3_SFF_0_n10), .C2(KeyOut1[0]), .A(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_ScanFF_S3_SFF_0_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S3_SFF_0_U2 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S3_SFF_0_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S3_SFF_0_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S3_SFF_0_n7), .CK(clk), .Q(
        Key_Registers_INST1_S2_in[0]), .QN(
        Key_Registers_INST1_ScanFF_S3_SFF_0_n8) );
  OAI21_X1 Key_Registers_INST1_ScanFF_S3_SFF_1_U4 ( .B1(
        Key_Registers_INST1_n290), .B2(Key_Registers_INST1_ScanFF_S3_SFF_1_n7), 
        .A(Key_Registers_INST1_ScanFF_S3_SFF_1_n10), .ZN(
        Key_Registers_INST1_ScanFF_S3_SFF_1_n6) );
  OAI221_X1 Key_Registers_INST1_ScanFF_S3_SFF_1_U3 ( .B1(
        Key_Registers_INST1_n289), .B2(Key_Registers_INST1_S4_1_), .C1(
        Key_Registers_INST1_ScanFF_S3_SFF_1_n9), .C2(KeyOut1[1]), .A(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_ScanFF_S3_SFF_1_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S3_SFF_1_U2 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S3_SFF_1_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S3_SFF_1_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S3_SFF_1_n6), .CK(clk), .Q(
        Key_Registers_INST1_S2_in[1]), .QN(
        Key_Registers_INST1_ScanFF_S3_SFF_1_n7) );
  OAI21_X1 Key_Registers_INST1_ScanFF_S3_SFF_2_U4 ( .B1(
        Key_Registers_INST1_n290), .B2(Key_Registers_INST1_ScanFF_S3_SFF_2_n7), 
        .A(Key_Registers_INST1_ScanFF_S3_SFF_2_n10), .ZN(
        Key_Registers_INST1_ScanFF_S3_SFF_2_n6) );
  OAI221_X1 Key_Registers_INST1_ScanFF_S3_SFF_2_U3 ( .B1(
        Key_Registers_INST1_n289), .B2(Key_Registers_INST1_S4_2_), .C1(
        Key_Registers_INST1_ScanFF_S3_SFF_2_n9), .C2(KeyOut1[2]), .A(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_ScanFF_S3_SFF_2_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S3_SFF_2_U2 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S3_SFF_2_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S3_SFF_2_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S3_SFF_2_n6), .CK(clk), .Q(
        Key_Registers_INST1_S2_in[2]), .QN(
        Key_Registers_INST1_ScanFF_S3_SFF_2_n7) );
  OAI21_X1 Key_Registers_INST1_ScanFF_S3_SFF_3_U4 ( .B1(
        Key_Registers_INST1_n290), .B2(Key_Registers_INST1_ScanFF_S3_SFF_3_n7), 
        .A(Key_Registers_INST1_ScanFF_S3_SFF_3_n10), .ZN(
        Key_Registers_INST1_ScanFF_S3_SFF_3_n6) );
  OAI221_X1 Key_Registers_INST1_ScanFF_S3_SFF_3_U3 ( .B1(
        Key_Registers_INST1_n289), .B2(Key_Registers_INST1_S4_3_), .C1(
        Key_Registers_INST1_ScanFF_S3_SFF_3_n9), .C2(KeyOut1[3]), .A(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_ScanFF_S3_SFF_3_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S3_SFF_3_U2 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S3_SFF_3_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S3_SFF_3_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S3_SFF_3_n6), .CK(clk), .Q(
        Key_Registers_INST1_S2_in[3]), .QN(
        Key_Registers_INST1_ScanFF_S3_SFF_3_n7) );
  OAI21_X1 Key_Registers_INST1_ScanFF_S3_SFF_4_U4 ( .B1(
        Key_Registers_INST1_n290), .B2(Key_Registers_INST1_ScanFF_S3_SFF_4_n7), 
        .A(Key_Registers_INST1_ScanFF_S3_SFF_4_n10), .ZN(
        Key_Registers_INST1_ScanFF_S3_SFF_4_n6) );
  OAI221_X1 Key_Registers_INST1_ScanFF_S3_SFF_4_U3 ( .B1(
        Key_Registers_INST1_n289), .B2(Key_Registers_INST1_S4_4_), .C1(
        Key_Registers_INST1_ScanFF_S3_SFF_4_n9), .C2(KeyOut1[4]), .A(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_ScanFF_S3_SFF_4_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S3_SFF_4_U2 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S3_SFF_4_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S3_SFF_4_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S3_SFF_4_n6), .CK(clk), .Q(
        Key_Registers_INST1_S2_in[4]), .QN(
        Key_Registers_INST1_ScanFF_S3_SFF_4_n7) );
  OAI21_X1 Key_Registers_INST1_ScanFF_S3_SFF_5_U4 ( .B1(
        Key_Registers_INST1_n290), .B2(Key_Registers_INST1_ScanFF_S3_SFF_5_n7), 
        .A(Key_Registers_INST1_ScanFF_S3_SFF_5_n10), .ZN(
        Key_Registers_INST1_ScanFF_S3_SFF_5_n6) );
  OAI221_X1 Key_Registers_INST1_ScanFF_S3_SFF_5_U3 ( .B1(
        Key_Registers_INST1_n289), .B2(Key_Registers_INST1_S4_5_), .C1(
        Key_Registers_INST1_ScanFF_S3_SFF_5_n9), .C2(KeyOut1[5]), .A(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_ScanFF_S3_SFF_5_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S3_SFF_5_U2 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S3_SFF_5_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S3_SFF_5_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S3_SFF_5_n6), .CK(clk), .Q(
        Key_Registers_INST1_S2_in[5]), .QN(
        Key_Registers_INST1_ScanFF_S3_SFF_5_n7) );
  OAI21_X1 Key_Registers_INST1_ScanFF_S3_SFF_6_U4 ( .B1(
        Key_Registers_INST1_n290), .B2(Key_Registers_INST1_ScanFF_S3_SFF_6_n7), 
        .A(Key_Registers_INST1_ScanFF_S3_SFF_6_n10), .ZN(
        Key_Registers_INST1_ScanFF_S3_SFF_6_n6) );
  OAI221_X1 Key_Registers_INST1_ScanFF_S3_SFF_6_U3 ( .B1(
        Key_Registers_INST1_n289), .B2(Key_Registers_INST1_S4_6_), .C1(
        Key_Registers_INST1_ScanFF_S3_SFF_6_n9), .C2(KeyOut1[6]), .A(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_ScanFF_S3_SFF_6_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S3_SFF_6_U2 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S3_SFF_6_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S3_SFF_6_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S3_SFF_6_n6), .CK(clk), .Q(
        Key_Registers_INST1_S2_in[6]), .QN(
        Key_Registers_INST1_ScanFF_S3_SFF_6_n7) );
  OAI21_X1 Key_Registers_INST1_ScanFF_S3_SFF_7_U4 ( .B1(
        Key_Registers_INST1_n290), .B2(Key_Registers_INST1_ScanFF_S3_SFF_7_n7), 
        .A(Key_Registers_INST1_ScanFF_S3_SFF_7_n10), .ZN(
        Key_Registers_INST1_ScanFF_S3_SFF_7_n6) );
  OAI221_X1 Key_Registers_INST1_ScanFF_S3_SFF_7_U3 ( .B1(
        Key_Registers_INST1_n289), .B2(Key_Registers_INST1_S4_7_), .C1(
        Key_Registers_INST1_ScanFF_S3_SFF_7_n9), .C2(KeyOut1[7]), .A(
        Key_Registers_INST1_n290), .ZN(Key_Registers_INST1_ScanFF_S3_SFF_7_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S3_SFF_7_U2 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S3_SFF_7_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S3_SFF_7_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S3_SFF_7_n6), .CK(clk), .Q(
        Key_Registers_INST1_S2_in[7]), .QN(
        Key_Registers_INST1_ScanFF_S3_SFF_7_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_0_U5 ( .A1(
        Key_Registers_INST1_n284), .A2(Key_Registers_INST1_ScanFF_S7_SFF_0_n8), 
        .B1(Key_Registers_INST1_ScanFF_S7_SFF_0_n12), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_0_n10), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_0_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_0_U4 ( .A1(
        Key_Registers_INST1_n289), .A2(Key_Registers_INST1_S4_0_), .B1(
        Key_Registers_INST1_S8_0_), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_0_n11), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_0_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_0_U3 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_0_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_0_U2 ( .A(Key_Registers_INST1_n284), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_0_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S7_SFF_0_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S7_SFF_0_n7), .CK(clk), .Q(
        Key_Registers_INST1_S6_in[0]), .QN(
        Key_Registers_INST1_ScanFF_S7_SFF_0_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_1_U6 ( .A1(
        Key_Registers_INST1_n284), .A2(Key_Registers_INST1_ScanFF_S7_SFF_1_n8), 
        .B1(Key_Registers_INST1_ScanFF_S7_SFF_1_n13), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_1_n10), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_1_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_1_U5 ( .A1(
        Key_Registers_INST1_ScanFF_S7_SFF_1_n11), .A2(
        Key_Registers_INST1_S4_1_), .B1(Key_Registers_INST1_S8_1_), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_1_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_1_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_1_U4 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_1_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_1_U3 ( .A(
        Key_Registers_INST1_ScanFF_S7_SFF_1_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_1_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_1_U2 ( .A(Key_Registers_INST1_n284), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_1_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S7_SFF_1_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S7_SFF_1_n7), .CK(clk), .Q(
        Key_Registers_INST1_S6_in[1]), .QN(
        Key_Registers_INST1_ScanFF_S7_SFF_1_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_2_U6 ( .A1(
        Key_Registers_INST1_n284), .A2(Key_Registers_INST1_ScanFF_S7_SFF_2_n8), 
        .B1(Key_Registers_INST1_ScanFF_S7_SFF_2_n13), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_2_n10), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_2_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_2_U5 ( .A1(
        Key_Registers_INST1_ScanFF_S7_SFF_2_n11), .A2(
        Key_Registers_INST1_S4_2_), .B1(Key_Registers_INST1_S8_2_), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_2_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_2_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_2_U4 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_2_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_2_U3 ( .A(
        Key_Registers_INST1_ScanFF_S7_SFF_2_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_2_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_2_U2 ( .A(Key_Registers_INST1_n284), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_2_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S7_SFF_2_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S7_SFF_2_n7), .CK(clk), .Q(
        Key_Registers_INST1_S6_in[2]), .QN(
        Key_Registers_INST1_ScanFF_S7_SFF_2_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_3_U6 ( .A1(
        Key_Registers_INST1_n284), .A2(Key_Registers_INST1_ScanFF_S7_SFF_3_n8), 
        .B1(Key_Registers_INST1_ScanFF_S7_SFF_3_n13), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_3_n10), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_3_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_3_U5 ( .A1(
        Key_Registers_INST1_ScanFF_S7_SFF_3_n11), .A2(
        Key_Registers_INST1_S4_3_), .B1(Key_Registers_INST1_S8_3_), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_3_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_3_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_3_U4 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_3_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_3_U3 ( .A(
        Key_Registers_INST1_ScanFF_S7_SFF_3_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_3_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_3_U2 ( .A(Key_Registers_INST1_n284), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_3_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S7_SFF_3_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S7_SFF_3_n7), .CK(clk), .Q(
        Key_Registers_INST1_S6_in[3]), .QN(
        Key_Registers_INST1_ScanFF_S7_SFF_3_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_4_U6 ( .A1(
        Key_Registers_INST1_n284), .A2(Key_Registers_INST1_ScanFF_S7_SFF_4_n8), 
        .B1(Key_Registers_INST1_ScanFF_S7_SFF_4_n13), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_4_n10), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_4_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_4_U5 ( .A1(
        Key_Registers_INST1_ScanFF_S7_SFF_4_n11), .A2(
        Key_Registers_INST1_S4_4_), .B1(Key_Registers_INST1_S8_4_), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_4_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_4_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_4_U4 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_4_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_4_U3 ( .A(
        Key_Registers_INST1_ScanFF_S7_SFF_4_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_4_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_4_U2 ( .A(Key_Registers_INST1_n284), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_4_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S7_SFF_4_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S7_SFF_4_n7), .CK(clk), .Q(
        Key_Registers_INST1_S6_in[4]), .QN(
        Key_Registers_INST1_ScanFF_S7_SFF_4_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_5_U6 ( .A1(
        Key_Registers_INST1_n284), .A2(Key_Registers_INST1_ScanFF_S7_SFF_5_n8), 
        .B1(Key_Registers_INST1_ScanFF_S7_SFF_5_n13), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_5_n10), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_5_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_5_U5 ( .A1(
        Key_Registers_INST1_ScanFF_S7_SFF_5_n11), .A2(
        Key_Registers_INST1_S4_5_), .B1(Key_Registers_INST1_S8_5_), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_5_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_5_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_5_U4 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_5_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_5_U3 ( .A(
        Key_Registers_INST1_ScanFF_S7_SFF_5_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_5_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_5_U2 ( .A(Key_Registers_INST1_n284), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_5_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S7_SFF_5_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S7_SFF_5_n7), .CK(clk), .Q(
        Key_Registers_INST1_S6_in[5]), .QN(
        Key_Registers_INST1_ScanFF_S7_SFF_5_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_6_U6 ( .A1(
        Key_Registers_INST1_n284), .A2(Key_Registers_INST1_ScanFF_S7_SFF_6_n8), 
        .B1(Key_Registers_INST1_ScanFF_S7_SFF_6_n13), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_6_n10), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_6_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_6_U5 ( .A1(
        Key_Registers_INST1_ScanFF_S7_SFF_6_n11), .A2(
        Key_Registers_INST1_S4_6_), .B1(Key_Registers_INST1_S8_6_), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_6_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_6_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_6_U4 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_6_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_6_U3 ( .A(
        Key_Registers_INST1_ScanFF_S7_SFF_6_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_6_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_6_U2 ( .A(Key_Registers_INST1_n284), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_6_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S7_SFF_6_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S7_SFF_6_n7), .CK(clk), .Q(
        Key_Registers_INST1_S6_in[6]), .QN(
        Key_Registers_INST1_ScanFF_S7_SFF_6_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_7_U6 ( .A1(
        Key_Registers_INST1_n284), .A2(Key_Registers_INST1_ScanFF_S7_SFF_7_n8), 
        .B1(Key_Registers_INST1_ScanFF_S7_SFF_7_n13), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_7_n10), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_7_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S7_SFF_7_U5 ( .A1(
        Key_Registers_INST1_ScanFF_S7_SFF_7_n11), .A2(
        Key_Registers_INST1_S4_7_), .B1(Key_Registers_INST1_S8_7_), .B2(
        Key_Registers_INST1_ScanFF_S7_SFF_7_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_7_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_7_U4 ( .A(Key_Registers_INST1_n289), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_7_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_7_U3 ( .A(
        Key_Registers_INST1_ScanFF_S7_SFF_7_n12), .ZN(
        Key_Registers_INST1_ScanFF_S7_SFF_7_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S7_SFF_7_U2 ( .A(Key_Registers_INST1_n284), 
        .ZN(Key_Registers_INST1_ScanFF_S7_SFF_7_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S7_SFF_7_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S7_SFF_7_n7), .CK(clk), .Q(
        Key_Registers_INST1_S6_in[7]), .QN(
        Key_Registers_INST1_ScanFF_S7_SFF_7_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_0_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n10), .A2(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n8), .B1(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n14), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n11), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_0_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n12), .A2(
        Key_Registers_INST1_S8_0_), .B1(KeyForSchedule1[0]), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n13), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n14) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_0_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_0_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_0_U4 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n13), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_0_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_0_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_0_U2 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n11), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S11_SFF_0_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n7), .CK(clk), .Q(
        Key_Registers_INST1_S10_in[0]), .QN(
        Key_Registers_INST1_ScanFF_S11_SFF_0_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_1_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n10), .A2(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n8), .B1(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n14), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n11), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_1_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n12), .A2(
        Key_Registers_INST1_S8_1_), .B1(KeyForSchedule1[1]), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n13), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n14) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_1_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_1_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_1_U4 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n13), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_1_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_1_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_1_U2 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n11), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S11_SFF_1_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n7), .CK(clk), .Q(
        Key_Registers_INST1_S10_in[1]), .QN(
        Key_Registers_INST1_ScanFF_S11_SFF_1_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_2_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n10), .A2(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n8), .B1(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n14), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n11), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_2_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n12), .A2(
        Key_Registers_INST1_S8_2_), .B1(KeyForSchedule1[2]), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n13), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n14) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_2_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_2_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_2_U4 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n13), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_2_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_2_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_2_U2 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n11), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S11_SFF_2_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n7), .CK(clk), .Q(
        Key_Registers_INST1_S10_in[2]), .QN(
        Key_Registers_INST1_ScanFF_S11_SFF_2_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_3_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n10), .A2(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n8), .B1(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n14), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n11), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_3_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n12), .A2(
        Key_Registers_INST1_S8_3_), .B1(KeyForSchedule1[3]), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n13), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n14) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_3_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_3_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_3_U4 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n13), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_3_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_3_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_3_U2 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n11), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S11_SFF_3_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n7), .CK(clk), .Q(
        Key_Registers_INST1_S10_in[3]), .QN(
        Key_Registers_INST1_ScanFF_S11_SFF_3_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_4_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n10), .A2(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n8), .B1(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n14), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n11), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_4_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n12), .A2(
        Key_Registers_INST1_S8_4_), .B1(KeyForSchedule1[4]), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n13), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n14) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_4_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_4_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_4_U4 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n13), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_4_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_4_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_4_U2 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n11), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S11_SFF_4_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n7), .CK(clk), .Q(
        Key_Registers_INST1_S10_in[4]), .QN(
        Key_Registers_INST1_ScanFF_S11_SFF_4_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_5_U5 ( .A1(
        Key_Registers_INST1_n283), .A2(Key_Registers_INST1_ScanFF_S11_SFF_5_n7), .B1(Key_Registers_INST1_ScanFF_S11_SFF_5_n11), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_5_n9), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_5_n6) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_5_U4 ( .A1(
        Key_Registers_INST1_n289), .A2(Key_Registers_INST1_S8_5_), .B1(
        KeyForSchedule1[5]), .B2(Key_Registers_INST1_ScanFF_S11_SFF_5_n10), 
        .ZN(Key_Registers_INST1_ScanFF_S11_SFF_5_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_5_U3 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_5_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_5_U2 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_5_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S11_SFF_5_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S11_SFF_5_n6), .CK(clk), .Q(
        Key_Registers_INST1_S10_in[5]), .QN(
        Key_Registers_INST1_ScanFF_S11_SFF_5_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_6_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n9), .A2(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n7), .B1(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n13), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n10), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n6) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_6_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n11), .A2(
        Key_Registers_INST1_S8_6_), .B1(KeyForSchedule1[6]), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n12), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_6_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_6_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_6_U4 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n12), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_6_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_6_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_6_U2 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n10), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S11_SFF_6_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n6), .CK(clk), .Q(
        Key_Registers_INST1_S10_in[6]), .QN(
        Key_Registers_INST1_ScanFF_S11_SFF_6_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_7_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n9), .A2(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n7), .B1(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n13), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n10), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n6) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S11_SFF_7_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n11), .A2(
        Key_Registers_INST1_S8_7_), .B1(KeyForSchedule1[7]), .B2(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n12), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_7_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_7_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_7_U4 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n12), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_7_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S11_SFF_7_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S11_SFF_7_U2 ( .A(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n10), .ZN(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S11_SFF_7_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n6), .CK(clk), .Q(
        Key_Registers_INST1_S10_in[7]), .QN(
        Key_Registers_INST1_ScanFF_S11_SFF_7_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_0_U5 ( .A1(
        Key_Registers_INST1_n283), .A2(Key_Registers_INST1_ScanFF_S15_SFF_0_n8), .B1(Key_Registers_INST1_ScanFF_S15_SFF_0_n12), .B2(
        Key_Registers_INST1_ScanFF_S15_SFF_0_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_0_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_0_U4 ( .A1(
        Key_Registers_INST1_n289), .A2(KeyForSchedule1[0]), .B1(KeyIn1[0]), 
        .B2(Key_Registers_INST1_ScanFF_S15_SFF_0_n11), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_0_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_0_U3 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_0_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_0_U2 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_0_n10) );
  DFF_X1 Key_Registers_INST1_ScanFF_S15_SFF_0_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S15_SFF_0_n7), .CK(clk), .Q(
        Key_Registers_INST1_S14_in[0]), .QN(
        Key_Registers_INST1_ScanFF_S15_SFF_0_n8) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_1_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n9), .A2(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n7), .B1(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n13), .B2(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n6) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_1_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n11), .A2(KeyForSchedule1[1]), 
        .B1(KeyIn1[1]), .B2(Key_Registers_INST1_ScanFF_S15_SFF_1_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_1_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_1_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_1_U4 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_1_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_1_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_1_U2 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S15_SFF_1_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n6), .CK(clk), .Q(
        Key_Registers_INST1_S14_in[1]), .QN(
        Key_Registers_INST1_ScanFF_S15_SFF_1_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_2_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n9), .A2(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n7), .B1(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n13), .B2(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n6) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_2_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n11), .A2(KeyForSchedule1[2]), 
        .B1(KeyIn1[2]), .B2(Key_Registers_INST1_ScanFF_S15_SFF_2_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_2_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_2_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_2_U4 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_2_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_2_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_2_U2 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S15_SFF_2_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n6), .CK(clk), .Q(
        Key_Registers_INST1_S14_in[2]), .QN(
        Key_Registers_INST1_ScanFF_S15_SFF_2_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_3_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n9), .A2(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n7), .B1(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n13), .B2(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n6) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_3_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n11), .A2(KeyForSchedule1[3]), 
        .B1(KeyIn1[3]), .B2(Key_Registers_INST1_ScanFF_S15_SFF_3_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_3_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_3_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_3_U4 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_3_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_3_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_3_U2 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S15_SFF_3_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n6), .CK(clk), .Q(
        Key_Registers_INST1_S14_in[3]), .QN(
        Key_Registers_INST1_ScanFF_S15_SFF_3_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_4_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n9), .A2(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n7), .B1(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n13), .B2(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n6) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_4_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n11), .A2(KeyForSchedule1[4]), 
        .B1(KeyIn1[4]), .B2(Key_Registers_INST1_ScanFF_S15_SFF_4_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_4_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_4_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_4_U4 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_4_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_4_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_4_U2 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S15_SFF_4_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n6), .CK(clk), .Q(
        Key_Registers_INST1_S14_in[4]), .QN(
        Key_Registers_INST1_ScanFF_S15_SFF_4_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_5_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n9), .A2(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n7), .B1(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n13), .B2(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n6) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_5_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n11), .A2(KeyForSchedule1[5]), 
        .B1(KeyIn1[5]), .B2(Key_Registers_INST1_ScanFF_S15_SFF_5_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_5_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_5_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_5_U4 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_5_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_5_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_5_U2 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S15_SFF_5_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n6), .CK(clk), .Q(
        Key_Registers_INST1_S14_in[5]), .QN(
        Key_Registers_INST1_ScanFF_S15_SFF_5_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_6_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n9), .A2(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n7), .B1(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n13), .B2(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n6) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_6_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n11), .A2(KeyForSchedule1[6]), 
        .B1(KeyIn1[6]), .B2(Key_Registers_INST1_ScanFF_S15_SFF_6_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_6_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_6_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_6_U4 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_6_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_6_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_6_U2 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S15_SFF_6_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n6), .CK(clk), .Q(
        Key_Registers_INST1_S14_in[6]), .QN(
        Key_Registers_INST1_ScanFF_S15_SFF_6_n7) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_7_U7 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n9), .A2(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n7), .B1(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n13), .B2(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n6) );
  AOI22_X1 Key_Registers_INST1_ScanFF_S15_SFF_7_U6 ( .A1(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n11), .A2(KeyForSchedule1[7]), 
        .B1(KeyIn1[7]), .B2(Key_Registers_INST1_ScanFF_S15_SFF_7_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n13) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_7_U5 ( .A(Key_Registers_INST1_n289), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_7_n12) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_7_U4 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n12), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n11) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_7_U3 ( .A(Key_Registers_INST1_n283), .ZN(Key_Registers_INST1_ScanFF_S15_SFF_7_n10) );
  INV_X1 Key_Registers_INST1_ScanFF_S15_SFF_7_U2 ( .A(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n10), .ZN(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n9) );
  DFF_X1 Key_Registers_INST1_ScanFF_S15_SFF_7_Q_reg ( .D(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n6), .CK(clk), .Q(
        Key_Registers_INST1_S14_in[7]), .QN(
        Key_Registers_INST1_ScanFF_S15_SFF_7_n7) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U14 ( .A(SboxIn1[4]), .B(
        GF256Inv_o_InputAffine_Inst1_inv_input1[1]), .Z(
        GF256Inv_o_InputAffine_Inst1_inv_input1[6]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U13 ( .A(SboxIn1[1]), .B(
        GF256Inv_o_InputAffine_Inst1_inv_input1[1]), .Z(
        GF256Inv_o_InputAffine_Inst1_inv_input1[5]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U12 ( .A(SboxIn1[1]), .B(
        GF256Inv_o_InputAffine_Inst1_A1_n9), .Z(
        GF256Inv_o_InputAffine_Inst1_inv_input1[3]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U11 ( .A(
        GF256Inv_o_InputAffine_Inst1_A1_n8), .B(
        GF256Inv_o_InputAffine_Inst1_A1_n7), .ZN(
        GF256Inv_o_InputAffine_Inst1_A1_n9) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U10 ( .A(
        GF256Inv_o_InputAffine_Inst1_inv_input1[2]), .B(SboxIn1[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_A1_n7) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U9 ( .A(SboxIn1[4]), .B(SboxIn1[3]), 
        .Z(GF256Inv_o_InputAffine_Inst1_A1_n8) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U8 ( .A(
        GF256Inv_o_InputAffine_Inst1_A1_n6), .B(SboxIn1[3]), .Z(
        GF256Inv_o_InputAffine_Inst1_inv_input1[0]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U7 ( .A(
        GF256Inv_o_InputAffine_Inst1_A1_n5), .B(
        GF256Inv_o_InputAffine_Inst1_A1_n4), .ZN(
        GF256Inv_o_InputAffine_Inst1_inv_input1[4]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U6 ( .A(
        GF256Inv_o_InputAffine_Inst1_A1_n6), .B(
        GF256Inv_o_InputAffine_Inst1_A1_n4), .ZN(
        GF256Inv_o_InputAffine_Inst1_inv_input1[7]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U5 ( .A(SboxIn1[5]), .B(SboxIn1[7]), 
        .ZN(GF256Inv_o_InputAffine_Inst1_A1_n4) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U4 ( .A(
        GF256Inv_o_InputAffine_Inst1_A1_n3), .B(SboxIn1[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_A1_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U3 ( .A(
        GF256Inv_o_InputAffine_Inst1_A1_n5), .B(SboxIn1[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_A1_n3) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U2 ( .A(
        GF256Inv_o_InputAffine_Inst1_A1_n5), .B(SboxIn1[5]), .Z(
        GF256Inv_o_InputAffine_Inst1_inv_input1[1]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A1_U1 ( .A(
        GF256Inv_o_InputAffine_Inst1_inv_input1[2]), .B(SboxIn1[6]), .Z(
        GF256Inv_o_InputAffine_Inst1_A1_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U14 ( .A(n167), .B(
        GF256Inv_o_InputAffine_Inst1_inv_input2[1]), .Z(
        GF256Inv_o_InputAffine_Inst1_inv_input2[6]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U13 ( .A(n164), .B(
        GF256Inv_o_InputAffine_Inst1_inv_input2[1]), .Z(
        GF256Inv_o_InputAffine_Inst1_inv_input2[5]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U12 ( .A(n164), .B(
        GF256Inv_o_InputAffine_Inst1_A2_n28), .Z(
        GF256Inv_o_InputAffine_Inst1_inv_input2[3]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U11 ( .A(
        GF256Inv_o_InputAffine_Inst1_A2_n27), .B(
        GF256Inv_o_InputAffine_Inst1_A2_n26), .ZN(
        GF256Inv_o_InputAffine_Inst1_A2_n28) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U10 ( .A(
        GF256Inv_o_InputAffine_Inst1_inv_input2[2]), .B(n170), .ZN(
        GF256Inv_o_InputAffine_Inst1_A2_n26) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U9 ( .A(n167), .B(n166), .Z(
        GF256Inv_o_InputAffine_Inst1_A2_n27) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U8 ( .A(
        GF256Inv_o_InputAffine_Inst1_A2_n25), .B(n166), .Z(
        GF256Inv_o_InputAffine_Inst1_inv_input2[0]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U7 ( .A(
        GF256Inv_o_InputAffine_Inst1_A2_n24), .B(
        GF256Inv_o_InputAffine_Inst1_A2_n23), .ZN(
        GF256Inv_o_InputAffine_Inst1_inv_input2[4]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U6 ( .A(
        GF256Inv_o_InputAffine_Inst1_A2_n25), .B(
        GF256Inv_o_InputAffine_Inst1_A2_n23), .ZN(
        GF256Inv_o_InputAffine_Inst1_inv_input2[7]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U5 ( .A(n168), .B(n170), .ZN(
        GF256Inv_o_InputAffine_Inst1_A2_n23) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U4 ( .A(
        GF256Inv_o_InputAffine_Inst1_A2_n22), .B(n165), .ZN(
        GF256Inv_o_InputAffine_Inst1_A2_n25) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U3 ( .A(
        GF256Inv_o_InputAffine_Inst1_A2_n24), .B(n164), .ZN(
        GF256Inv_o_InputAffine_Inst1_A2_n22) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U2 ( .A(
        GF256Inv_o_InputAffine_Inst1_A2_n24), .B(n168), .Z(
        GF256Inv_o_InputAffine_Inst1_inv_input2[1]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_A2_U1 ( .A(
        GF256Inv_o_InputAffine_Inst1_inv_input2[2]), .B(n169), .Z(
        GF256Inv_o_InputAffine_Inst1_A2_n24) );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_0_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input1[0]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_1_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input1[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_2_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input1[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_3_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input1[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_4_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input1[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_5_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input1[5]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_6_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input1[6]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_7_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input1[7]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_8_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input2[0]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_9_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input2[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_10_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input2[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_11_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input2[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_12_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input2[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_13_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input2[5]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_14_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input2[6]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_GEN_reg1_s_current_state_reg_15_ ( .D(
        GF256Inv_o_InputAffine_Inst1_inv_input2[7]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg1_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg1[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg1_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg1[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg1_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg1[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg1_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg1[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg1_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg1[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg1_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg1[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg1_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg1[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg1_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg1[3]), .QN() );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U51 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n81), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n80), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu[1]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U50 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n79), .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n78), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n80) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U49 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n78) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U48 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n81), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n77), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd[1]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U47 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n76), .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n75), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n77) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U46 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n76) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U45 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n74), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n73), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n81) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U44 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n72), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n71), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n74) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U43 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n70), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n69), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu[1]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U42 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n68), .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n67), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n69) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U41 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n66), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n70), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd[1]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U40 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n65), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n64), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n70) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U39 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n63), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n62), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n65) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U38 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n62) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U37 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n71), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n61), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n63) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U36 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n60), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n59), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n71) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U35 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n58), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n57), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n59) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U34 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n57) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U33 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n58) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U32 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n56), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n55), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n60) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U31 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n55) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U30 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n56) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U29 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n54), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n66) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U28 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n53), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n52), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu[1]) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U27 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n52) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U26 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n72), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n61), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n53) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U25 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n51), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n54), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n72) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U24 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n54) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U23 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n50), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n49), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n51) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U22 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n75), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n68), .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n49) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U21 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n68) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U20 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n64), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n48), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n50) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U19 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n48) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U18 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n67), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n79), .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n64) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U17 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n67) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U16 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n47), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U15 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n47), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td[1]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U14 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n73), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n46), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n47) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U13 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n45), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n44), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n46) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U12 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n79), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n75), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n44) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U11 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n75) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U10 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n79) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U9 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n61), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n43), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n45) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U8 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .C1(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .C2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n42), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n43) );
  OAI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U7 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .B1(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n42) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n41), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n40), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n61) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U5 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n40) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U4 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n41) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n39), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n38), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n73) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U2 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n38) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U1 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n39) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U60 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n59), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n58), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu[2]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U59 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n57), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n58) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U58 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n56), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n55), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd[3]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U57 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n57), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n55) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U56 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n54), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n53), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n57) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U55 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n52), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n51), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n54) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U54 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n50), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n49), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n52) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U53 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n48), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n47), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n56) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U52 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n46), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n45), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n48) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U51 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n44), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n43), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n45) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U50 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n42), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n46) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U49 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n47), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n41), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U48 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n41), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n40), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd[3]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U47 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n39), .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n38), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n40) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U46 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n37), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n36), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n41) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U45 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n35), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n34), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n36) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U44 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n33), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n32), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n35) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U43 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n50), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n31), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n37) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U42 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n30), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n29), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n50) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U41 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n29) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U40 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n28), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n27), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n30) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U39 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n26), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n25), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n27) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U38 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n25) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U37 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n26) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U36 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n24), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n23), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu[2]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U35 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n22), .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n43), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n23) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U34 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n24), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n59), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd[3]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U33 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n28), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n59) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U32 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n28) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U31 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n21), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n53), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n24) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U30 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n20), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n19), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n53) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U29 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n33), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n18), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n19) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U28 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n18) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U27 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n33) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U26 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n31), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n17), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n20) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U25 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n17) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U24 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n44), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n22), .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n31) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U23 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n44) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U22 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n16), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U21 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n47), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n16), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td[3]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U20 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n21), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n15), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n16) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U19 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n15) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U18 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U17 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n51), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U16 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n22), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n38), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n43), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U15 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n43) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U14 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n38) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U13 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n11), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n10), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n51) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U12 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n10) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U11 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n11) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U10 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n9), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n49), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n21) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U9 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n49) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U8 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n34), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n8), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n9) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U7 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n42), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n32), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n8) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U6 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n32) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U5 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n42) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U4 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n34) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U3 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n39), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n22), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n47) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U2 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n22) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U1 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n39) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U61 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n61), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n60), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu[3]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U60 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n59), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n58), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n57), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n60) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U59 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n56), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n55), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n61) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U58 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n55), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U57 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n54), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n53), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n55) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U56 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n52), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n51), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n53) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U55 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n50), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n49), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n51) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U54 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n58), .A2(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n49) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U53 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n48), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n47), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n50) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U52 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n46), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n45), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n52) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U51 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n44), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n59), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu[3]) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U50 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n58), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n59) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U49 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n43), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n42), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n58) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U48 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n44), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n41), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U47 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n40), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n39), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n44) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U46 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n38), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n37), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n40) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U45 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n36), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n47), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n37) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U44 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n35), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n34), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n47) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U43 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n33), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n32), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n34) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U42 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n31), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n30), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n32) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U41 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n30) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U40 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n31) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U39 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n43), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n29), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n35) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U38 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n57), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n28), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n38) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U37 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n27), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n26), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd[2]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U36 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n29), .B1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n26) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U35 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n41), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu[3]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U34 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n43), .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n41) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U33 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U32 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n43), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U31 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U30 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n56), .A2(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U29 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n29), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n56) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U28 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U27 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U26 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n17), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U25 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n16), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n45), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U24 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n45) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U23 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n28), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n42), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n16) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U22 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n29), .B1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n15), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n28) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U21 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n15), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n14), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n57), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U20 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n15) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U19 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n27), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n46), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu[3]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U18 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n33), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n46) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U17 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n33) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U16 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n13), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n48), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n27) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U15 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n57), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n42), .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n48) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U14 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n42) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U13 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n12), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n17), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n13) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U12 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n36), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n11), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n17) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U11 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n11) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U10 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n36) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U9 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n54), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n10), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n12) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U8 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n57), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n43), .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n10) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U7 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n57) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n39), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n54) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U5 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U4 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n29), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n14), .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n39) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U3 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n14) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U2 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n29) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U1 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n43) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U58 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n98), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n97), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu[4]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U57 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n96), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n95), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n98) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U56 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n94), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n97), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd[4]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U55 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n93), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n92), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n97) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U54 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n91), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n90), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n93) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U53 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n90) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U52 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n89), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n88), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n91) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U51 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n87), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n86), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n88) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U50 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n85), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n84), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n86) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U49 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n83), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n82), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n85) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U48 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n81), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n82) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U47 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n80), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n83) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U46 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n79), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n78), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n87) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U45 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n77), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n78), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu[4]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U44 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n76), .B1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n75), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n78) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U43 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n77), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n74), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd[4]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U42 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n79), .B1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n95), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n74) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U41 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n79) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U40 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n73), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n72), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n77) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U39 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n71), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n92), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n73) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U38 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n70), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n69), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n92) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U37 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n70) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U36 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n68), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n69), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu[4]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U35 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n67), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n66), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n69) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U34 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n66) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U33 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n80), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n75), .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n67) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U32 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n65), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n68) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U31 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U30 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n89), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n65) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U29 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n61), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U28 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n59), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n61) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U27 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n59) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U26 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n80), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n96), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U25 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n96) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U24 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n80) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U23 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U22 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n95), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n76), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n89) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U21 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n76) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U20 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n95) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U19 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n71), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n56), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu[4]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U18 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n54), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n56) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U17 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n94), .A2(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n54) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U16 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n84), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n53), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U15 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n52), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n53) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U14 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .B2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n72), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U13 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n72) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U12 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n52) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U11 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n51), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n50), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n84) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U10 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n50) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U9 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n51) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U8 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n49), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n71) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U7 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n48), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n47), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U6 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n47) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U5 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n48) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U4 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n94), .A2(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n49) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U3 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n75), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n81), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n94) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U2 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n81) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U1 ( 
        .A(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n75) );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_0_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_1_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_2_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_3_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_4_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_5_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_6_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_7_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_8_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_9_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_10_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_11_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_12_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_13_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_14_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_15_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_0_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_1_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_2_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_3_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_4_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_5_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_6_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_7_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_8_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_9_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_10_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_11_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_12_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_13_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_14_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_GEN_reg01_s_current_state_reg_15_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td_reg[4]), .QN() );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L1_XORInst0_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu_reg[2]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1[1]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L1_XORInst1_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xu_reg[4]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2[1]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L1_XORInst2_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu_reg[2]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1[2]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L1_XORInst3_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yu_reg[4]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2[2]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L1_XORInst4_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu_reg[2]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1[3]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L1_XORInst5_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zu_reg[4]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2[3]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L1_XORInst6_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu_reg[2]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1[4]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L1_XORInst7_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_tu_reg[4]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2[4]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L2_XORInst0_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd_reg[2]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1[1]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L2_XORInst1_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_xd_reg[4]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2[1]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L2_XORInst2_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd_reg[2]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1[2]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L2_XORInst3_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_yd_reg[4]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2[2]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L2_XORInst4_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd_reg[2]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1[3]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L2_XORInst5_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_zd_reg[4]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2[3]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L2_XORInst6_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td_reg[2]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1[4]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L2_XORInst7_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf6_sq_scl_mul_Canright_td_reg[4]), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2[4]) );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg2_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg1[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg2_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[5]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg1[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg2_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[6]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg1[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg2_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input1_reg[7]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg1[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg2_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg1[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg2_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[5]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg1[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg2_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[6]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg1[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg2_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_inv_input2_reg[7]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg1[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg3_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg1[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg2[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg3_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg1[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg2[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg3_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg1[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg2[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg3_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg1[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg2[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg3_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg1[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg2[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg3_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg1[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg2[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg3_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg1[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg2[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg3_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg1[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg2[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4u_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4u_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4u_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4u_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4u_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4u_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4u_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4u_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4d_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4d_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4d_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4d_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4d_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4d_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4d_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg4d_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg5_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg1[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg2[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg5_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg1[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg2[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg5_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg1[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg2[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg5_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg1[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg2[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg5_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg1[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg2[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg5_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg1[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg2[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg5_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg1[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg2[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg5_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg1[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg2[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg6_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg2[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg3[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg6_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg2[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg3[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg6_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg2[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg3[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg6_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg2[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg3[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg6_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg2[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg3[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg6_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg2[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg3[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg6_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg2[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg3[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg6_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg2[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg3[3]), .QN() );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_U4 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n7), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[1]) );
  OAI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_U3 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n7) );
  AND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9) );
  OAI33_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_U4 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14), .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .B3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[2])
         );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U12 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[3]) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U11 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U10 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U9 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[3]) );
  OAI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U8 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U7 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[3])
         );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U5 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U4 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U3 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[3]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U2 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_U1 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U14 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n61), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[4]) );
  NAND3_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U13 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n61) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U12 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n59), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[4]) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U11 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n59) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U10 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n56), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[4]) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U9 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n56) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U8 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U7 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U6 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[4]) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U5 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U4 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_U4 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_n8), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_n6), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[5]) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_U3 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_n6) );
  AND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F5_n8) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U12 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40), .C1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n39), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n38), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[5]) );
  NOR3_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U11 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n39), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n38) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U10 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n37), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n39) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U9 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n36), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[5]) );
  OAI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U8 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n35), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n36) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U7 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n37) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U6 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n35), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[6]) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U5 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n35) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U4 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40) );
  NOR3_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n33), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[5]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_U1 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n37), .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F6_n33) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_U10 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n25), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[7]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_U9 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n25) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_U8 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n24), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n23), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[7]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_U7 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n24), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n23) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n24) );
  NOR3_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_U5 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n22), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[7]) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_U4 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n22) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n21), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n20), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[7]) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n20) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_U1 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F7_n21) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U11 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n28), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[8]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U10 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n28) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U9 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n27), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[8]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U8 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n26), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n27) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U7 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n25), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n24), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[8]) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U6 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n25), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n23), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n24) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U5 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n25) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U4 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n23), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n26), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n22), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[8]) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n22) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n23), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n26) );
  AND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_U1 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F8_n23) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_U8 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n20), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[1]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_U7 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n20) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_U6 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n19), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n18), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[1]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_U5 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n19), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n18) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_U4 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n19) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_U3 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n16), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n17), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[1]) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n16), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n17) );
  AND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_U1 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F9_n16) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_U8 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n17), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[2]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_U7 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n17) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_U6 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n16), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[2]) );
  OAI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_U5 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n16) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_U4 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n15), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n14), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n13), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[2]) );
  NAND3_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_U3 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n15), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[1]), 
        .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n13) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n14) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_U1 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F10_n15) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U11 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n24), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n23), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n22), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[6]) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U10 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n22) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U9 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n21), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n24), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n20), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[6])
         );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U8 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n21), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n20) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U7 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n23), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n21) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n23) );
  OAI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U5 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n19), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n18), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n17), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[6]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U4 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n19), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n17) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U3 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n24), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n18) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n24) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_sq_scl_mul_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_N_F11_n19) );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_0_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_1_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_2_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_3_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_4_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[5]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[5]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_5_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[6]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[6]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_6_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[7]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[7]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_7_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x[8]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[8]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_8_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_9_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_10_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_11_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_12_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[5]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[5]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_13_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[6]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[6]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_14_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[7]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[7]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_15_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y[8]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[8]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_16_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_17_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_18_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_19_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_20_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[5]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[5]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_21_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[6]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[6]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_22_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[7]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[7]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_23_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z[8]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[8]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_24_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_25_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_26_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_27_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_28_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[5]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[5]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_29_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[6]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[6]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_30_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[7]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[7]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_GEN_reg_s_current_state_reg_31_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t[8]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[8]), .QN() );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1[0]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[3]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[1]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2[0]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[7]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[8]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[5]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_x_reg[6]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[3]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[1]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[7]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[8]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[5]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_y_reg[6]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[3]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[1]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[7]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[8]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[5]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_z_reg[6]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1[3]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[3]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[1]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2[3]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[7]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[8]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[5]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_t_reg[6]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_u_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n6) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_U4 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n7), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[1]) );
  OAI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_U3 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n7) );
  AND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9) );
  OAI33_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_U4 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14), .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .B3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[2])
         );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U12 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[3]) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U11 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U10 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U9 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[3]) );
  OAI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U8 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U7 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[3])
         );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U5 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U4 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U3 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[3]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U2 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_U1 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U14 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n61), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[4]) );
  NAND3_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U13 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n61) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U12 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n59), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[4]) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U11 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n59) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U10 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n56), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[4]) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U9 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n56) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U8 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n62) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U7 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n57) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U6 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[4]) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U5 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n63) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U4 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n64) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n58) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n55) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F4_n60) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_U4 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_n8), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_n6), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[5]) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_U3 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_n6) );
  AND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F5_n8) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U12 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40), .C1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n39), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n38), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[5]) );
  NOR3_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U11 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n39), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n38) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U10 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n37), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n39) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U9 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n36), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[5]) );
  OAI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U8 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n35), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n36) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U7 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n37) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U6 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n35), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[6]) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U5 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n35) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U4 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40) );
  NOR3_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n33), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[5]) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_U1 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n37), .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n40), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F6_n33) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_U10 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n25), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[7]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_U9 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n25) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_U8 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n24), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n23), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[7]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_U7 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n24), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n23) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n24) );
  NOR3_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_U5 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n22), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[7]) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_U4 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n22) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n21), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n20), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[7]) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n20) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_U1 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F7_n21) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U11 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n28), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[8]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U10 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n28) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U9 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n27), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[8]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U8 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n26), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n27) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U7 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n25), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n24), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[8]) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U6 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n25), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n23), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n24) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U5 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n25) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U4 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n23), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n26), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n22), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[8]) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n22) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n23), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n26) );
  AND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_U1 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F8_n23) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_U8 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n20), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[1]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_U7 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n20) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_U6 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n19), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n18), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[1]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_U5 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n19), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n18) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_U4 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n19) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_U3 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n16), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n17), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[1]) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_U2 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n16), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n17) );
  AND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_U1 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F9_n16) );
  AOI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_U8 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n17), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[2]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_U7 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n17) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_U6 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n16), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[2]) );
  OAI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_U5 ( 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n16) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_U4 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n15), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n14), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n13), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[2]) );
  NAND3_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_U3 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n15), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[1]), 
        .A3(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n13) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n14) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_U1 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F10_n15) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U11 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n24), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n23), .C2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n22), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[6]) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U10 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n22) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U9 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n21), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n24), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n20), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[6])
         );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U8 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n21), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n20) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U7 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n23), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n21) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n23) );
  OAI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U5 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n19), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n18), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n17), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[6]) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U4 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n19), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n17) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U3 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[2]), 
        .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n24), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n18) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n24) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_sq_scl_mul_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_N_F11_n19) );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_0_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_1_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_2_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_3_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_4_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[5]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[5]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_5_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[6]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[6]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_6_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[7]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[7]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_7_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x[8]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[8]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_8_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_9_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_10_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_11_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_12_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[5]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[5]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_13_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[6]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[6]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_14_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[7]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[7]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_15_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y[8]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[8]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_16_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_17_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_18_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_19_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_20_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[5]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[5]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_21_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[6]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[6]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_22_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[7]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[7]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_23_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z[8]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[8]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_24_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_25_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_26_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_27_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[4]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_28_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[5]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[5]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_29_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[6]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[6]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_30_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[7]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[7]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_GEN_reg_s_current_state_reg_31_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t[8]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[8]), .QN() );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1[0]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[3]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[1]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2[0]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[7]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[8]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[5]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_x_reg[6]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[3]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[1]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[7]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[8]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[5]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_y_reg[6]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[3]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[1]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[7]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[8]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[5]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_z_reg[6]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1[3]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[3]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[4]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[1]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n6) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n6), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n5), .ZN(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2[3]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[7]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[8]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n5) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[5]), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_t_reg[6]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_GF16_inv_282_d_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n6) );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg7_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg2[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg3[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg7_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg2[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg3[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg7_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg2[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg3[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg7_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg2[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg3[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg7_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg2[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg3[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg7_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg2[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg3[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg7_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg2[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg3[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg7_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg2[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg3[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg8_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg3[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg8_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg3[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg8_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg3[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg8_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg3[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg8_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg3[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg8_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg3[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg8_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg3[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg8_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg3[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9u_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1[0]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9u_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9u_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9u_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9u_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2[0]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9u_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9u_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[2]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9u_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[3]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9d_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1[0]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9d_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9d_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9d_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9d_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2[0]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9d_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2[1]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9d_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2[2]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[2]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg9d_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2[3]), 
        .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[3]), 
        .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg10_s_current_state_reg_0_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg3[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg10_s_current_state_reg_1_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg3[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg10_s_current_state_reg_2_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg3[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg10_s_current_state_reg_3_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg3[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg10_s_current_state_reg_4_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg3[0]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[0]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg10_s_current_state_reg_5_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg3[1]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg10_s_current_state_reg_6_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg3[2]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_GEN_reg10_s_current_state_reg_7_ ( 
        .D(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg3[3]), .CK(clk), .Q(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .QN() );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U47 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n133), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n132), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U46 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n131), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n130), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n133) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U45 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n130) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U44 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n129), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n131) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U43 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n128), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n129) );
  OAI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U42 ( 
        .C1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U41 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U40 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U39 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U38 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U37 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U36 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U35 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U34 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U33 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U32 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U31 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U30 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U29 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n132), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U28 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n132) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U27 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U26 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U25 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U24 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U23 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U22 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U21 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U20 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U19 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U18 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U17 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U16 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U15 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U14 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U13 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n128), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U12 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n128) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U11 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U10 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U9 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U8 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U7 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U5 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U4 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U3 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U1 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U44 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z[2]) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U43 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U42 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U41 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U40 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U39 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U38 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U37 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U36 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U35 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U34 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U33 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U32 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U31 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U30 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U29 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U28 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U27 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U26 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U25 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U24 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U23 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U22 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U21 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U20 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[3]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U19 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U18 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U17 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U16 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U15 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U14 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U13 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U12 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U11 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[2]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U10 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U9 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U8 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U7 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U6 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U5 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n100), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U4 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[2]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[1]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n100) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U3 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U2 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U1 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U43 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z[3]) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U42 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U41 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U40 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U39 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U38 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U37 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U36 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y[3]) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U35 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U34 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U33 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U32 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U31 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U30 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U29 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U28 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U27 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U26 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x[3]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U25 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U24 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U23 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[0]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U22 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U21 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U20 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n110), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n109), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U19 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n109) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U18 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[0]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U17 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n110) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U16 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n108), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U15 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n107), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n106), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t[3]) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U14 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n106) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U13 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U12 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n105), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n107) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U11 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n104), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n103), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n105) );
  MUX2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U10 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .S(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n103) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U9 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U8 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U7 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n108), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n104) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U6 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n108) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U5 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U4 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n102), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n101), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U2 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n101) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U1 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n102) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U46 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y[4]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U45 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U44 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U43 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U42 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U41 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U40 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x[4]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U39 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U38 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U37 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[0]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U36 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U35 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U34 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U33 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[3]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U32 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U31 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U30 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U29 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U28 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U27 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[3]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U26 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U25 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U24 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t[4]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U23 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U22 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U21 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U20 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U19 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110) );
  MUX2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U18 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .S(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U17 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U16 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U15 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U14 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U13 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U12 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U11 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U10 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z[4]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U9 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U8 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[1]), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[2]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U7 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U5 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_dcba2_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U4 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U3 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[2]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U2 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[3]), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n98), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U1 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_u_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n98) );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_0_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_1_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_2_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_3_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_4_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_5_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_6_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_7_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_8_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_9_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_10_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_11_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_12_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_13_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_14_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_15_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t_reg[4]), .QN() );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst0_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x_reg[2]), .Z(StateIn1[4]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_x_reg[4]), .Z(StateIn2[4]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y_reg[2]), .Z(StateIn1[5]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_y_reg[4]), .Z(StateIn2[5]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z_reg[2]), .Z(StateIn1[6]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_z_reg[4]), .Z(StateIn2[6]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t_reg[2]), .Z(StateIn1[7]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright1_t_reg[4]), .Z(StateIn2[7]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U47 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n133), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n132), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U46 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n131), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n130), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n133) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U45 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n130) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U44 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n129), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n131) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U43 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n128), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n129) );
  OAI211_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U42 ( 
        .C1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U41 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U40 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U39 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U38 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U37 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U36 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U35 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U34 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U33 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U32 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U31 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U30 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U29 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n132), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U28 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n132) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U27 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U26 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U25 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U24 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U23 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U22 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U21 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U20 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U19 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U18 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U17 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t[1]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U16 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U15 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U14 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U13 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n128), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U12 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n128) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U11 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U10 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U9 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U8 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U7 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U5 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U4 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U3 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U2 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U1 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U44 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z[2]) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U43 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U42 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U41 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U40 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U39 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U38 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U37 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128) );
  NOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U36 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U35 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U34 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U33 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U32 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U31 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U30 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U29 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U28 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U27 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U26 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U25 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U24 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U23 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U22 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110) );
  OAI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U21 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U20 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[3]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U19 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U18 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U17 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t[2]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U16 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U15 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U14 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U13 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U12 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U11 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[2]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U10 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U9 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U8 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U7 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U6 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U5 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n100), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U4 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[2]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[1]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n100) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U3 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U2 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U1 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe1_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U43 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z[3]) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U42 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U41 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U40 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U39 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U38 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U37 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U36 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y[3]) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U35 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U34 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U33 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U32 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[0]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U31 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U30 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U29 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U28 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U27 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U26 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x[3]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U25 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U24 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U23 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[0]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U22 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U21 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U20 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n110), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n109), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U19 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n109) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U18 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[0]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U17 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n110) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U16 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n108), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U15 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n107), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n106), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t[3]) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U14 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n106) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U13 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U12 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n105), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n107) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U11 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n104), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n103), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n105) );
  MUX2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U10 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .S(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n103) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U9 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U8 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U7 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114), .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n108), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n104) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U6 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n108) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U5 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U4 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U3 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n102), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n101), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U2 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n101) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U1 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out1_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n102) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U46 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132), .Z(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y[4]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U45 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U44 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U43 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U42 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U41 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U40 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x[4]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U39 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U38 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U37 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[0]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U36 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U35 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U34 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U33 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[3]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U32 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U31 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U30 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U29 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U28 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U27 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[3]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U26 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115), .B(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U25 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U24 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t[4]) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U23 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113) );
  AOI22_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U22 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U21 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[3]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U20 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U19 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110) );
  MUX2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U18 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .S(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[2]), 
        .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U17 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[0]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U16 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U15 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U14 ( 
        .A1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .A2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108) );
  OAI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U13 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .B2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U12 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[3]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U11 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U10 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z[4]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U9 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U8 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[1]), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[2]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U7 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[2]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104) );
  XNOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U6 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103) );
  NAND2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U5 ( 
        .A1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136), .A2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_hgfe2_reg4[2]), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U4 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100), .Z(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101) );
  AOI21_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U3 ( 
        .B1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[2]), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100) );
  AOI221_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U2 ( 
        .B1(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[3]), .B2(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), 
        .C1(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136), .C2(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n98), .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99) );
  INV_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U1 ( 
        .A(GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_d_GF16_inv_out2_reg[0]), 
        .ZN(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n98) );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_0_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_1_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_2_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_3_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_4_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_5_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_6_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_7_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_8_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_9_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_10_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_11_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z_reg[4]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_12_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t[1]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t_reg[1]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_13_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t[2]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t_reg[2]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_14_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t[3]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t_reg[3]), .QN() );
  DFF_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_15_ ( 
        .D(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t[4]), .CK(clk), .Q(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t_reg[4]), .QN() );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst0_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x_reg[2]), .Z(StateIn1[0]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_x_reg[4]), .Z(StateIn2[0]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y_reg[2]), .Z(StateIn1[1]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_y_reg[4]), .Z(StateIn2[1]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z_reg[2]), .Z(StateIn1[2]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_z_reg[4]), .Z(StateIn2[2]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t_reg[1]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t_reg[2]), .Z(StateIn1[3]) );
  XOR2_X1 GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U1 ( 
        .A(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t_reg[3]), .B(
        GF256Inv_o_InputAffine_Inst1_Inst_GF256_INV_Inst_Gf16_mul2_Canright2_t_reg[4]), .Z(StateIn2[3]) );
  NOR3_X1 Inst_Controller_U96 ( .A1(Inst_Controller_n173), .A2(
        Inst_Controller_n172), .A3(Inst_Controller_n171), .ZN(ShowRcon) );
  AOI21_X1 Inst_Controller_U95 ( .B1(Inst_Controller_n166), .B2(
        Inst_Controller_n35), .A(Inst_Controller_n165), .ZN(
        Inst_Controller_n113) );
  AOI22_X1 Inst_Controller_U94 ( .A1(Inst_Controller_n91), .A2(
        Inst_Controller_n165), .B1(Inst_Controller_n164), .B2(
        Inst_Controller_n116), .ZN(Inst_Controller_n112) );
  INV_X1 Inst_Controller_U93 ( .A(Inst_Controller_n163), .ZN(
        Inst_Controller_n164) );
  AOI22_X1 Inst_Controller_U92 ( .A1(Inst_Controller_n33), .A2(
        Inst_Controller_n169), .B1(Inst_Controller_n162), .B2(
        Inst_Controller_n122), .ZN(Inst_Controller_n111) );
  INV_X1 Inst_Controller_U91 ( .A(Inst_Controller_n167), .ZN(
        Inst_Controller_n162) );
  OAI21_X1 Inst_Controller_U90 ( .B1(rst), .B2(Inst_Controller_n91), .A(
        Inst_Controller_n165), .ZN(Inst_Controller_n167) );
  AOI21_X1 Inst_Controller_U89 ( .B1(Inst_Controller_n35), .B2(
        Inst_Controller_n168), .A(Inst_Controller_n166), .ZN(
        Inst_Controller_n165) );
  NAND2_X1 Inst_Controller_U88 ( .A1(Inst_Controller_n91), .A2(
        Inst_Controller_n163), .ZN(Inst_Controller_n169) );
  NOR2_X1 Inst_Controller_U87 ( .A1(Inst_Controller_n35), .A2(
        Inst_Controller_n161), .ZN(Inst_Controller_n163) );
  OAI22_X1 Inst_Controller_U86 ( .A1(Inst_Controller_n19), .A2(
        Inst_Controller_n160), .B1(Inst_Controller_n20), .B2(
        Inst_Controller_n161), .ZN(Inst_Controller_n110) );
  OAI221_X1 Inst_Controller_U85 ( .B1(Inst_Controller_n159), .B2(
        Inst_Controller_n19), .C1(Inst_Controller_n160), .C2(
        Inst_Controller_n26), .A(Inst_Controller_n168), .ZN(
        Inst_Controller_n109) );
  OAI21_X1 Inst_Controller_U84 ( .B1(Inst_Controller_n25), .B2(
        Inst_Controller_n160), .A(Inst_Controller_n158), .ZN(
        Inst_Controller_n108) );
  OAI221_X1 Inst_Controller_U83 ( .B1(Inst_Controller_n19), .B2(
        Inst_Controller_n26), .C1(Rcon_internal[7]), .C2(Rcon_internal[0]), 
        .A(Inst_Controller_n157), .ZN(Inst_Controller_n158) );
  OAI22_X1 Inst_Controller_U82 ( .A1(Inst_Controller_n24), .A2(
        Inst_Controller_n160), .B1(Inst_Controller_n25), .B2(
        Inst_Controller_n161), .ZN(Inst_Controller_n107) );
  OAI21_X1 Inst_Controller_U81 ( .B1(Inst_Controller_n23), .B2(
        Inst_Controller_n160), .A(Inst_Controller_n156), .ZN(
        Inst_Controller_n106) );
  OAI221_X1 Inst_Controller_U80 ( .B1(Inst_Controller_n19), .B2(
        Inst_Controller_n24), .C1(Rcon_internal[7]), .C2(Rcon_internal[2]), 
        .A(Inst_Controller_n157), .ZN(Inst_Controller_n156) );
  OAI21_X1 Inst_Controller_U79 ( .B1(Inst_Controller_n22), .B2(
        Inst_Controller_n160), .A(Inst_Controller_n155), .ZN(
        Inst_Controller_n105) );
  OAI221_X1 Inst_Controller_U78 ( .B1(Inst_Controller_n19), .B2(
        Inst_Controller_n23), .C1(Rcon_internal[7]), .C2(Rcon_internal[3]), 
        .A(Inst_Controller_n157), .ZN(Inst_Controller_n155) );
  INV_X1 Inst_Controller_U77 ( .A(Inst_Controller_n161), .ZN(
        Inst_Controller_n157) );
  OAI22_X1 Inst_Controller_U76 ( .A1(Inst_Controller_n22), .A2(
        Inst_Controller_n161), .B1(Inst_Controller_n21), .B2(
        Inst_Controller_n160), .ZN(Inst_Controller_n104) );
  OAI22_X1 Inst_Controller_U75 ( .A1(Inst_Controller_n21), .A2(
        Inst_Controller_n161), .B1(Inst_Controller_n20), .B2(
        Inst_Controller_n160), .ZN(Inst_Controller_n103) );
  NAND2_X1 Inst_Controller_U74 ( .A1(Inst_Controller_n168), .A2(
        Inst_Controller_n160), .ZN(Inst_Controller_n161) );
  NAND2_X1 Inst_Controller_U73 ( .A1(Inst_Controller_n178), .A2(
        Inst_Controller_n154), .ZN(key_reg_hold) );
  AOI21_X1 Inst_Controller_U72 ( .B1(Inst_Controller_n39), .B2(
        Inst_Controller_n152), .A(rst), .ZN(SboxIn_sel[0]) );
  AOI21_X1 Inst_Controller_U71 ( .B1(Inst_Controller_n151), .B2(
        Inst_Controller_n176), .A(Inst_Controller_n119), .ZN(
        Inst_Controller_n152) );
  AOI221_X1 Inst_Controller_U70 ( .B1(Inst_Controller_n37), .B2(
        Inst_Controller_n148), .C1(Inst_Controller_n119), .C2(
        Inst_Controller_n147), .A(Inst_Controller_n146), .ZN(
        Inst_Controller_N86) );
  INV_X1 Inst_Controller_U69 ( .A(Inst_Controller_n148), .ZN(
        Inst_Controller_n147) );
  OAI211_X1 Inst_Controller_U68 ( .C1(Inst_Controller_n118), .C2(
        Inst_Controller_n144), .A(Inst_Controller_n148), .B(
        Inst_Controller_n166), .ZN(Inst_Controller_n145) );
  NAND2_X1 Inst_Controller_U67 ( .A1(Inst_Controller_n118), .A2(
        Inst_Controller_n144), .ZN(Inst_Controller_n148) );
  AOI211_X1 Inst_Controller_U66 ( .C1(Inst_Controller_n6), .C2(
        Inst_Controller_n149), .A(Inst_Controller_n144), .B(
        Inst_Controller_n146), .ZN(Inst_Controller_N84) );
  NOR2_X1 Inst_Controller_U65 ( .A1(Inst_Controller_n6), .A2(
        Inst_Controller_n149), .ZN(Inst_Controller_n144) );
  NOR2_X1 Inst_Controller_U64 ( .A1(Inst_Controller_n146), .A2(
        Inst_Controller_n143), .ZN(Inst_Controller_N83) );
  AOI21_X1 Inst_Controller_U63 ( .B1(Inst_Controller_n154), .B2(
        Inst_Controller_n170), .A(Inst_Controller_n146), .ZN(
        Inst_Controller_N82) );
  INV_X1 Inst_Controller_U62 ( .A(Inst_Controller_n166), .ZN(
        Inst_Controller_n146) );
  AOI21_X1 Inst_Controller_U61 ( .B1(Inst_Controller_n142), .B2(
        Inst_Controller_n37), .A(Inst_Controller_n160), .ZN(
        Inst_Controller_n166) );
  NOR2_X1 Inst_Controller_U60 ( .A1(rst), .A2(Inst_Controller_n141), .ZN(
        Inst_Controller_n159) );
  NOR2_X1 Inst_Controller_U59 ( .A1(Inst_Controller_n151), .A2(
        Inst_Controller_n140), .ZN(Inst_Controller_n142) );
  NAND2_X1 Inst_Controller_U58 ( .A1(Inst_Controller_n139), .A2(
        Inst_Controller_n177), .ZN(Inst_Controller_n140) );
  NAND2_X1 Inst_Controller_U57 ( .A1(Inst_Controller_n94), .A2(
        Inst_Controller_PerRoundCounter_0_), .ZN(Inst_Controller_n170) );
  OAI21_X1 Inst_Controller_U56 ( .B1(Inst_Controller_PerRoundCounter_0_), .B2(
        Inst_Controller_n141), .A(Inst_Controller_n168), .ZN(
        Inst_Controller_N81) );
  AND3_X1 Inst_Controller_U55 ( .A1(Inst_Controller_n138), .A2(
        Inst_Controller_n137), .A3(Inst_Controller_n136), .ZN(
        Inst_Controller_n141) );
  NAND3_X1 Inst_Controller_U54 ( .A1(Inst_Controller_n137), .A2(
        Inst_Controller_n168), .A3(Inst_Controller_n133), .ZN(
        Inst_Controller_n134) );
  AOI221_X1 Inst_Controller_U53 ( .B1(Inst_Controller_n94), .B2(
        Inst_Controller_n132), .C1(Inst_Controller_n115), .C2(
        Inst_Controller_n171), .A(Inst_Controller_n173), .ZN(
        KeyScheduleRegisterEN) );
  NOR2_X1 Inst_Controller_U52 ( .A1(Inst_Controller_n131), .A2(
        Inst_Controller_n130), .ZN(KeyIn_sel[1]) );
  NOR2_X1 Inst_Controller_U51 ( .A1(Inst_Controller_n129), .A2(
        Inst_Controller_n130), .ZN(KeyIn_sel[0]) );
  OAI211_X1 Inst_Controller_U50 ( .C1(Inst_Controller_n128), .C2(
        Inst_Controller_n133), .A(Inst_Controller_n168), .B(
        Inst_Controller_n151), .ZN(Inst_Controller_n130) );
  NAND2_X1 Inst_Controller_U49 ( .A1(Inst_Controller_n37), .A2(
        Inst_Controller_n150), .ZN(Inst_Controller_n133) );
  NOR2_X1 Inst_Controller_U48 ( .A1(Inst_Controller_n139), .A2(
        Inst_Controller_n171), .ZN(Inst_Controller_n150) );
  NAND3_X1 Inst_Controller_U47 ( .A1(Inst_Controller_n33), .A2(
        Inst_Controller_n120), .A3(Inst_Controller_n116), .ZN(
        Inst_Controller_n128) );
  INV_X1 Inst_Controller_U46 ( .A(Inst_Controller_n131), .ZN(
        Inst_Controller_n129) );
  NOR3_X1 Inst_Controller_U45 ( .A1(Inst_Controller_n119), .A2(
        Inst_Controller_n143), .A3(Inst_Controller_n127), .ZN(
        Inst_Controller_n131) );
  OAI21_X1 Inst_Controller_U44 ( .B1(Inst_Controller_n139), .B2(
        Inst_Controller_n117), .A(Inst_Controller_n149), .ZN(
        Inst_Controller_n143) );
  NAND2_X1 Inst_Controller_U43 ( .A1(Inst_Controller_n139), .A2(
        Inst_Controller_n117), .ZN(Inst_Controller_n149) );
  NOR2_X1 Inst_Controller_U42 ( .A1(Inst_Controller_n126), .A2(
        Inst_Controller_n175), .ZN(done_internal) );
  AOI22_X1 Inst_Controller_U41 ( .A1(Inst_Controller_n39), .A2(
        Inst_Controller_n135), .B1(Inst_Controller_n177), .B2(
        Inst_Controller_n172), .ZN(Inst_Controller_n126) );
  NAND3_X1 Inst_Controller_U40 ( .A1(Inst_Controller_n6), .A2(
        Inst_Controller_n44), .A3(Inst_Controller_n172), .ZN(
        Inst_Controller_n135) );
  OAI21_X1 Inst_Controller_U39 ( .B1(Inst_Controller_n173), .B2(
        Inst_Controller_n174), .A(Inst_Controller_n124), .ZN(DoKeySbox) );
  OAI211_X1 Inst_Controller_U38 ( .C1(Inst_Controller_n123), .C2(
        Inst_Controller_n139), .A(Inst_Controller_n37), .B(
        Inst_Controller_n177), .ZN(Inst_Controller_n124) );
  NOR3_X1 Inst_Controller_U37 ( .A1(Inst_Controller_n39), .A2(
        Inst_Controller_n117), .A3(Inst_Controller_n121), .ZN(
        Inst_Controller_n177) );
  INV_X1 Inst_Controller_U36 ( .A(Inst_Controller_n172), .ZN(
        Inst_Controller_n139) );
  NAND2_X1 Inst_Controller_U35 ( .A1(Inst_Controller_n138), .A2(
        Inst_Controller_n172), .ZN(Inst_Controller_n174) );
  NOR3_X1 Inst_Controller_U34 ( .A1(Inst_Controller_n44), .A2(
        Inst_Controller_n39), .A3(Inst_Controller_n121), .ZN(
        Inst_Controller_n138) );
  NAND2_X1 Inst_Controller_U33 ( .A1(Inst_Controller_n37), .A2(
        Inst_Controller_n125), .ZN(Inst_Controller_n175) );
  AND4_X1 Inst_Controller_U32 ( .A1(Inst_Controller_n90), .A2(
        Inst_Controller_n33), .A3(Inst_Controller_n91), .A4(
        Inst_Controller_n35), .ZN(Inst_Controller_n125) );
  OR2_X1 Inst_Controller_U31 ( .A1(Inst_Controller_n127), .A2(
        Inst_Controller_n44), .ZN(Inst_Controller_n132) );
  NAND2_X1 Inst_Controller_U30 ( .A1(Inst_Controller_n39), .A2(
        Inst_Controller_n6), .ZN(Inst_Controller_n127) );
  NOR3_X1 Inst_Controller_U29 ( .A1(Inst_Controller_n173), .A2(
        Inst_Controller_n170), .A3(Inst_Controller_n171), .ZN(DoSR) );
  NAND2_X1 Inst_Controller_U28 ( .A1(Inst_Controller_n115), .A2(
        Inst_Controller_PerRoundCounter_0_), .ZN(Inst_Controller_n172) );
  NAND3_X1 Inst_Controller_U27 ( .A1(Inst_Controller_n44), .A2(
        Inst_Controller_n39), .A3(Inst_Controller_n6), .ZN(
        Inst_Controller_n171) );
  NOR2_X1 Inst_Controller_U26 ( .A1(Inst_Controller_n94), .A2(
        Inst_Controller_PerRoundCounter_0_), .ZN(Inst_Controller_n136) );
  NOR3_X1 Inst_Controller_U25 ( .A1(Inst_Controller_n173), .A2(
        Inst_Controller_n154), .A3(Inst_Controller_n171), .ZN(
        JustFirstColShift) );
  NAND4_X1 Inst_Controller_U24 ( .A1(Inst_Controller_n120), .A2(
        Inst_Controller_n116), .A3(Inst_Controller_n33), .A4(
        Inst_Controller_n35), .ZN(Inst_Controller_n151) );
  INV_X1 Inst_Controller_U23 ( .A(Inst_Controller_n151), .ZN(
        Inst_Controller_n123) );
  NOR2_X1 Inst_Controller_U22 ( .A1(Inst_Controller_n123), .A2(
        Inst_Controller_n119), .ZN(Inst_Controller_n137) );
  NAND4_X1 Inst_Controller_U21 ( .A1(Inst_Controller_n39), .A2(
        Inst_Controller_n44), .A3(Inst_Controller_n6), .A4(
        Inst_Controller_n172), .ZN(Inst_Controller_n153) );
  NOR2_X1 Inst_Controller_U20 ( .A1(Inst_Controller_n173), .A2(
        Inst_Controller_n153), .ZN(Inst_Controller_n178) );
  NAND2_X1 Inst_Controller_U19 ( .A1(Inst_Controller_n178), .A2(
        Inst_Controller_n115), .ZN(state_reg_hold) );
  INV_X1 Inst_Controller_U18 ( .A(rst), .ZN(Inst_Controller_n168) );
  INV_X1 Inst_Controller_U17 ( .A(Inst_Controller_n136), .ZN(
        Inst_Controller_n154) );
  INV_X1 Inst_Controller_U16 ( .A(Inst_Controller_n159), .ZN(
        Inst_Controller_n160) );
  INV_X1 Inst_Controller_U15 ( .A(Inst_Controller_n137), .ZN(
        Inst_Controller_n173) );
  NOR4_X1 Inst_Controller_U14 ( .A1(Inst_Controller_n125), .A2(
        Inst_Controller_n173), .A3(Inst_Controller_n118), .A4(
        Inst_Controller_n172), .ZN(Inst_Controller_n179) );
  BUF_X1 Inst_Controller_U13 ( .A(Inst_Controller_n179), .Z(DoMC) );
  NOR4_X2 Inst_Controller_U12 ( .A1(Inst_Controller_PerRoundCounter_0_), .A2(
        Inst_Controller_n115), .A3(Inst_Controller_n132), .A4(
        Inst_Controller_n175), .ZN(Corr_63_5_) );
  AOI21_X2 Inst_Controller_U11 ( .B1(Inst_Controller_n118), .B2(
        Inst_Controller_n135), .A(Inst_Controller_n134), .ZN(SboxIn_sel[1]) );
  INV_X1 Inst_Controller_U9 ( .A(Inst_Controller_n90), .ZN(
        Inst_Controller_n100) );
  AOI21_X1 Inst_Controller_U8 ( .B1(Inst_Controller_n168), .B2(
        Inst_Controller_n33), .A(Inst_Controller_n167), .ZN(
        Inst_Controller_n99) );
  NAND2_X1 Inst_Controller_U7 ( .A1(Inst_Controller_n174), .A2(
        Inst_Controller_n98), .ZN(Output_Sel) );
  NOR3_X1 Inst_Controller_U6 ( .A1(Inst_Controller_n176), .A2(
        Inst_Controller_n177), .A3(Inst_Controller_n175), .ZN(
        Inst_Controller_n98) );
  NAND3_X1 Inst_Controller_U5 ( .A1(Inst_Controller_n149), .A2(
        Inst_Controller_n6), .A3(Inst_Controller_n97), .ZN(
        Inst_Controller_n176) );
  INV_X1 Inst_Controller_U4 ( .A(Inst_Controller_n150), .ZN(
        Inst_Controller_n97) );
  OAI33_X1 Inst_Controller_U3 ( .A1(1'b0), .A2(Inst_Controller_n99), .A3(
        Inst_Controller_n100), .B1(Inst_Controller_n90), .B2(
        Inst_Controller_n33), .B3(Inst_Controller_n169), .ZN(
        Inst_Controller_n114) );
  DFF_X1 Inst_Controller_RoundCounter_reg_3_ ( .D(Inst_Controller_n114), .CK(
        clk), .Q(Inst_Controller_n90), .QN(Inst_Controller_n120) );
  DFF_X1 Inst_Controller_RoundCounter_reg_2_ ( .D(Inst_Controller_n111), .CK(
        clk), .Q(Inst_Controller_n122), .QN(Inst_Controller_n33) );
  DFF_X1 Inst_Controller_PerRoundCounter_reg_5_ ( .D(Inst_Controller_N86), 
        .CK(clk), .Q(Inst_Controller_n119), .QN(Inst_Controller_n37) );
  DFF_X1 Inst_Controller_PerRoundCounter_reg_3_ ( .D(Inst_Controller_N84), 
        .CK(clk), .Q(Inst_Controller_n121), .QN(Inst_Controller_n6) );
  DFF_X1 Inst_Controller_Rcon_Reg_reg_1_ ( .D(Inst_Controller_n108), .CK(clk), 
        .Q(Rcon_internal[1]), .QN(Inst_Controller_n25) );
  DFF_X1 Inst_Controller_Rcon_Reg_reg_3_ ( .D(Inst_Controller_n106), .CK(clk), 
        .Q(Rcon_internal[3]), .QN(Inst_Controller_n23) );
  DFF_X1 Inst_Controller_Rcon_Reg_reg_4_ ( .D(Inst_Controller_n105), .CK(clk), 
        .Q(Rcon_internal[4]), .QN(Inst_Controller_n22) );
  DFF_X1 Inst_Controller_RoundCounter_reg_1_ ( .D(Inst_Controller_n112), .CK(
        clk), .Q(Inst_Controller_n91), .QN(Inst_Controller_n116) );
  DFF_X1 Inst_Controller_PerRoundCounter_reg_1_ ( .D(Inst_Controller_N82), 
        .CK(clk), .Q(Inst_Controller_n115), .QN(Inst_Controller_n94) );
  DFF_X1 Inst_Controller_PerRoundCounter_reg_2_ ( .D(Inst_Controller_N83), 
        .CK(clk), .Q(Inst_Controller_n117), .QN(Inst_Controller_n44) );
  DFF_X1 Inst_Controller_PerRoundCounter_reg_4_ ( .D(Inst_Controller_n145), 
        .CK(clk), .Q(Inst_Controller_n39), .QN(Inst_Controller_n118) );
  DFF_X1 Inst_Controller_Rcon_Reg_reg_2_ ( .D(Inst_Controller_n107), .CK(clk), 
        .Q(Rcon_internal[2]), .QN(Inst_Controller_n24) );
  DFF_X1 Inst_Controller_Rcon_Reg_reg_7_ ( .D(Inst_Controller_n110), .CK(clk), 
        .Q(Rcon_internal[7]), .QN(Inst_Controller_n19) );
  DFF_X1 Inst_Controller_Rcon_Reg_reg_5_ ( .D(Inst_Controller_n104), .CK(clk), 
        .Q(Rcon_internal[5]), .QN(Inst_Controller_n21) );
  DFF_X1 Inst_Controller_Rcon_Reg_reg_6_ ( .D(Inst_Controller_n103), .CK(clk), 
        .Q(Rcon_internal[6]), .QN(Inst_Controller_n20) );
  DFF_X1 Inst_Controller_Rcon_Reg_reg_0_ ( .D(Inst_Controller_n109), .CK(clk), 
        .Q(Rcon_internal[0]), .QN(Inst_Controller_n26) );
  DFF_X1 Inst_Controller_PerRoundCounter_reg_0_ ( .D(Inst_Controller_N81), 
        .CK(clk), .Q(Inst_Controller_PerRoundCounter_0_), .QN() );
  DFF_X1 Inst_Controller_RoundCounter_reg_0_ ( .D(Inst_Controller_n113), .CK(
        clk), .Q(), .QN(Inst_Controller_n35) );
endmodule

