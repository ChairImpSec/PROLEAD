module circuit ( plaintext_s0, key_s0, clk, start, plaintext_s1,
        key_s1, Fresh, ciphertext_s0, done, ciphertext_s1 );
  input [127:0] plaintext_s0;
  input [127:0] key_s0;
  input [127:0] plaintext_s1;
  input [127:0] key_s1;
  input [67:0] Fresh;
  output [127:0] ciphertext_s0;
  output [127:0] ciphertext_s1;
  input clk, start;
  output done;
  wire   new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1987,
         new_AGEMA_signal_1986, new_AGEMA_signal_1990, new_AGEMA_signal_1989,
         new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1996,
         new_AGEMA_signal_1995, new_AGEMA_signal_1999, new_AGEMA_signal_1998,
         new_AGEMA_signal_2002, new_AGEMA_signal_2001, new_AGEMA_signal_2005,
         new_AGEMA_signal_2004, ctrl_N14, ctrl_n6, ctrl_seq6_SFF_0_QD,
         ctrl_seq6_SFF_1_QD, ctrl_seq6_SFF_2_QD, ctrl_seq6_SFF_3_QD,
         ctrl_seq6_SFF_4_QD, ctrl_seq4_SFF_0_QD, ctrl_seq4_SFF_1_QD,
         new_AGEMA_signal_3126, stateArray_S00reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2156, new_AGEMA_signal_3127,
         stateArray_S00reg_gff_1_SFF_1_QD, new_AGEMA_signal_2159,
         new_AGEMA_signal_3128, stateArray_S00reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2162, new_AGEMA_signal_3129,
         stateArray_S00reg_gff_1_SFF_3_QD, new_AGEMA_signal_2165,
         new_AGEMA_signal_3130, stateArray_S00reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2168, new_AGEMA_signal_3131,
         stateArray_S00reg_gff_1_SFF_5_QD, new_AGEMA_signal_2171,
         new_AGEMA_signal_3132, stateArray_S00reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2174, new_AGEMA_signal_3133,
         stateArray_S00reg_gff_1_SFF_7_QD, new_AGEMA_signal_2177,
         new_AGEMA_signal_3134, stateArray_S01reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2180, new_AGEMA_signal_3135,
         stateArray_S01reg_gff_1_SFF_1_QD, new_AGEMA_signal_2183,
         new_AGEMA_signal_3136, stateArray_S01reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2186, new_AGEMA_signal_3137,
         stateArray_S01reg_gff_1_SFF_3_QD, new_AGEMA_signal_2189,
         new_AGEMA_signal_3138, stateArray_S01reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2192, new_AGEMA_signal_3139,
         stateArray_S01reg_gff_1_SFF_5_QD, new_AGEMA_signal_2195,
         new_AGEMA_signal_3140, stateArray_S01reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2198, new_AGEMA_signal_3141,
         stateArray_S01reg_gff_1_SFF_7_QD, new_AGEMA_signal_2201,
         new_AGEMA_signal_3142, stateArray_S02reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2204, new_AGEMA_signal_3143,
         stateArray_S02reg_gff_1_SFF_1_QD, new_AGEMA_signal_2207,
         new_AGEMA_signal_3144, stateArray_S02reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2210, new_AGEMA_signal_3145,
         stateArray_S02reg_gff_1_SFF_3_QD, new_AGEMA_signal_2213,
         new_AGEMA_signal_3146, stateArray_S02reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2216, new_AGEMA_signal_3147,
         stateArray_S02reg_gff_1_SFF_5_QD, new_AGEMA_signal_2219,
         new_AGEMA_signal_3148, stateArray_S02reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2222, new_AGEMA_signal_3149,
         stateArray_S02reg_gff_1_SFF_7_QD, new_AGEMA_signal_2225,
         new_AGEMA_signal_3150, stateArray_S03reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_3046, new_AGEMA_signal_3151,
         stateArray_S03reg_gff_1_SFF_1_QD, new_AGEMA_signal_3048,
         new_AGEMA_signal_3152, stateArray_S03reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_3050, new_AGEMA_signal_3153,
         stateArray_S03reg_gff_1_SFF_3_QD, new_AGEMA_signal_3052,
         new_AGEMA_signal_3154, stateArray_S03reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_3054, new_AGEMA_signal_3155,
         stateArray_S03reg_gff_1_SFF_5_QD, new_AGEMA_signal_3056,
         new_AGEMA_signal_3156, stateArray_S03reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_3058, new_AGEMA_signal_3157,
         stateArray_S03reg_gff_1_SFF_7_QD, new_AGEMA_signal_3060,
         new_AGEMA_signal_3158, stateArray_S10reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2228, new_AGEMA_signal_3159,
         stateArray_S10reg_gff_1_SFF_1_QD, new_AGEMA_signal_2231,
         new_AGEMA_signal_3160, stateArray_S10reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2234, new_AGEMA_signal_3161,
         stateArray_S10reg_gff_1_SFF_3_QD, new_AGEMA_signal_2237,
         new_AGEMA_signal_3162, stateArray_S10reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2240, new_AGEMA_signal_3163,
         stateArray_S10reg_gff_1_SFF_5_QD, new_AGEMA_signal_2243,
         new_AGEMA_signal_3164, stateArray_S10reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2246, new_AGEMA_signal_3165,
         stateArray_S10reg_gff_1_SFF_7_QD, new_AGEMA_signal_2249,
         new_AGEMA_signal_3166, stateArray_S11reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2252, new_AGEMA_signal_3167,
         stateArray_S11reg_gff_1_SFF_1_QD, new_AGEMA_signal_2255,
         new_AGEMA_signal_3168, stateArray_S11reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2258, new_AGEMA_signal_3169,
         stateArray_S11reg_gff_1_SFF_3_QD, new_AGEMA_signal_2261,
         new_AGEMA_signal_3170, stateArray_S11reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2264, new_AGEMA_signal_3171,
         stateArray_S11reg_gff_1_SFF_5_QD, new_AGEMA_signal_2267,
         new_AGEMA_signal_3172, stateArray_S11reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2270, new_AGEMA_signal_3173,
         stateArray_S11reg_gff_1_SFF_7_QD, new_AGEMA_signal_2273,
         new_AGEMA_signal_3174, stateArray_S12reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2276, new_AGEMA_signal_3175,
         stateArray_S12reg_gff_1_SFF_1_QD, new_AGEMA_signal_2279,
         new_AGEMA_signal_3176, stateArray_S12reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2282, new_AGEMA_signal_3177,
         stateArray_S12reg_gff_1_SFF_3_QD, new_AGEMA_signal_2285,
         new_AGEMA_signal_3178, stateArray_S12reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2288, new_AGEMA_signal_3179,
         stateArray_S12reg_gff_1_SFF_5_QD, new_AGEMA_signal_2291,
         new_AGEMA_signal_3180, stateArray_S12reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2294, new_AGEMA_signal_3181,
         stateArray_S12reg_gff_1_SFF_7_QD, new_AGEMA_signal_2297,
         new_AGEMA_signal_3182, stateArray_S13reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_3062, new_AGEMA_signal_3183,
         stateArray_S13reg_gff_1_SFF_1_QD, new_AGEMA_signal_3064,
         new_AGEMA_signal_3184, stateArray_S13reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_3066, new_AGEMA_signal_3185,
         stateArray_S13reg_gff_1_SFF_3_QD, new_AGEMA_signal_3068,
         new_AGEMA_signal_3186, stateArray_S13reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_3070, new_AGEMA_signal_3187,
         stateArray_S13reg_gff_1_SFF_5_QD, new_AGEMA_signal_3072,
         new_AGEMA_signal_3188, stateArray_S13reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_3074, new_AGEMA_signal_3189,
         stateArray_S13reg_gff_1_SFF_7_QD, new_AGEMA_signal_3076,
         new_AGEMA_signal_3190, stateArray_S20reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2300, new_AGEMA_signal_3191,
         stateArray_S20reg_gff_1_SFF_1_QD, new_AGEMA_signal_2303,
         new_AGEMA_signal_3192, stateArray_S20reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2306, new_AGEMA_signal_3193,
         stateArray_S20reg_gff_1_SFF_3_QD, new_AGEMA_signal_2309,
         new_AGEMA_signal_3194, stateArray_S20reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2312, new_AGEMA_signal_3195,
         stateArray_S20reg_gff_1_SFF_5_QD, new_AGEMA_signal_2315,
         new_AGEMA_signal_3196, stateArray_S20reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2318, new_AGEMA_signal_3197,
         stateArray_S20reg_gff_1_SFF_7_QD, new_AGEMA_signal_2321,
         new_AGEMA_signal_3198, stateArray_S21reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2324, new_AGEMA_signal_3199,
         stateArray_S21reg_gff_1_SFF_1_QD, new_AGEMA_signal_2327,
         new_AGEMA_signal_3200, stateArray_S21reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2330, new_AGEMA_signal_3201,
         stateArray_S21reg_gff_1_SFF_3_QD, new_AGEMA_signal_2333,
         new_AGEMA_signal_3202, stateArray_S21reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2336, new_AGEMA_signal_3203,
         stateArray_S21reg_gff_1_SFF_5_QD, new_AGEMA_signal_2339,
         new_AGEMA_signal_3204, stateArray_S21reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2342, new_AGEMA_signal_3205,
         stateArray_S21reg_gff_1_SFF_7_QD, new_AGEMA_signal_2345,
         new_AGEMA_signal_3206, stateArray_S22reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2348, new_AGEMA_signal_3207,
         stateArray_S22reg_gff_1_SFF_1_QD, new_AGEMA_signal_2351,
         new_AGEMA_signal_3208, stateArray_S22reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2354, new_AGEMA_signal_3209,
         stateArray_S22reg_gff_1_SFF_3_QD, new_AGEMA_signal_2357,
         new_AGEMA_signal_3210, stateArray_S22reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2360, new_AGEMA_signal_3211,
         stateArray_S22reg_gff_1_SFF_5_QD, new_AGEMA_signal_2363,
         new_AGEMA_signal_3212, stateArray_S22reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2366, new_AGEMA_signal_3213,
         stateArray_S22reg_gff_1_SFF_7_QD, new_AGEMA_signal_2369,
         new_AGEMA_signal_3214, stateArray_S23reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_3078, new_AGEMA_signal_3215,
         stateArray_S23reg_gff_1_SFF_1_QD, new_AGEMA_signal_3080,
         new_AGEMA_signal_3216, stateArray_S23reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_3082, new_AGEMA_signal_3217,
         stateArray_S23reg_gff_1_SFF_3_QD, new_AGEMA_signal_3084,
         new_AGEMA_signal_3218, stateArray_S23reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_3086, new_AGEMA_signal_3219,
         stateArray_S23reg_gff_1_SFF_5_QD, new_AGEMA_signal_3088,
         new_AGEMA_signal_3220, stateArray_S23reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_3090, new_AGEMA_signal_3221,
         stateArray_S23reg_gff_1_SFF_7_QD, new_AGEMA_signal_3092,
         new_AGEMA_signal_3222, stateArray_S30reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2372, new_AGEMA_signal_3223,
         stateArray_S30reg_gff_1_SFF_1_QD, new_AGEMA_signal_2375,
         new_AGEMA_signal_3224, stateArray_S30reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2378, new_AGEMA_signal_3225,
         stateArray_S30reg_gff_1_SFF_3_QD, new_AGEMA_signal_2381,
         new_AGEMA_signal_3226, stateArray_S30reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2384, new_AGEMA_signal_3227,
         stateArray_S30reg_gff_1_SFF_5_QD, new_AGEMA_signal_2387,
         new_AGEMA_signal_3228, stateArray_S30reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2390, new_AGEMA_signal_3229,
         stateArray_S30reg_gff_1_SFF_7_QD, new_AGEMA_signal_2393,
         new_AGEMA_signal_3230, stateArray_S31reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2396, new_AGEMA_signal_3231,
         stateArray_S31reg_gff_1_SFF_1_QD, new_AGEMA_signal_2399,
         new_AGEMA_signal_3232, stateArray_S31reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2402, new_AGEMA_signal_3233,
         stateArray_S31reg_gff_1_SFF_3_QD, new_AGEMA_signal_2405,
         new_AGEMA_signal_3234, stateArray_S31reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2408, new_AGEMA_signal_3235,
         stateArray_S31reg_gff_1_SFF_5_QD, new_AGEMA_signal_2411,
         new_AGEMA_signal_3236, stateArray_S31reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2414, new_AGEMA_signal_3237,
         stateArray_S31reg_gff_1_SFF_7_QD, new_AGEMA_signal_2417,
         new_AGEMA_signal_3238, stateArray_S32reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_2420, new_AGEMA_signal_3239,
         stateArray_S32reg_gff_1_SFF_1_QD, new_AGEMA_signal_2423,
         new_AGEMA_signal_3240, stateArray_S32reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_2426, new_AGEMA_signal_3241,
         stateArray_S32reg_gff_1_SFF_3_QD, new_AGEMA_signal_2429,
         new_AGEMA_signal_3242, stateArray_S32reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_2432, new_AGEMA_signal_3243,
         stateArray_S32reg_gff_1_SFF_5_QD, new_AGEMA_signal_2435,
         new_AGEMA_signal_3244, stateArray_S32reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_2438, new_AGEMA_signal_3245,
         stateArray_S32reg_gff_1_SFF_7_QD, new_AGEMA_signal_2441,
         new_AGEMA_signal_3008, new_AGEMA_signal_2880, new_AGEMA_signal_3009,
         new_AGEMA_signal_2881, new_AGEMA_signal_3010, new_AGEMA_signal_2882,
         new_AGEMA_signal_3011, new_AGEMA_signal_2883, new_AGEMA_signal_3012,
         new_AGEMA_signal_2884, new_AGEMA_signal_3013, new_AGEMA_signal_2885,
         new_AGEMA_signal_3014, new_AGEMA_signal_2886, new_AGEMA_signal_3015,
         new_AGEMA_signal_2887, new_AGEMA_signal_3016, new_AGEMA_signal_2872,
         new_AGEMA_signal_3017, new_AGEMA_signal_2873, new_AGEMA_signal_3018,
         new_AGEMA_signal_2874, new_AGEMA_signal_3019, new_AGEMA_signal_2875,
         new_AGEMA_signal_3020, new_AGEMA_signal_2876, new_AGEMA_signal_3021,
         new_AGEMA_signal_2877, new_AGEMA_signal_3022, new_AGEMA_signal_2878,
         new_AGEMA_signal_3023, new_AGEMA_signal_2879, new_AGEMA_signal_3024,
         new_AGEMA_signal_2864, new_AGEMA_signal_3025, new_AGEMA_signal_2865,
         new_AGEMA_signal_3026, new_AGEMA_signal_2866, new_AGEMA_signal_3027,
         new_AGEMA_signal_2867, new_AGEMA_signal_3028, new_AGEMA_signal_2868,
         new_AGEMA_signal_3029, new_AGEMA_signal_2869, new_AGEMA_signal_3030,
         new_AGEMA_signal_2870, new_AGEMA_signal_3031, new_AGEMA_signal_2871,
         new_AGEMA_signal_2860, new_AGEMA_signal_2825, new_AGEMA_signal_2861,
         new_AGEMA_signal_2849, new_AGEMA_signal_2834, new_AGEMA_signal_2823,
         new_AGEMA_signal_2862, new_AGEMA_signal_2848, new_AGEMA_signal_2863,
         new_AGEMA_signal_2847, new_AGEMA_signal_2835, new_AGEMA_signal_2820,
         new_AGEMA_signal_2836, new_AGEMA_signal_2819, new_AGEMA_signal_2837,
         new_AGEMA_signal_2818, new_AGEMA_signal_2817, new_AGEMA_signal_2846,
         new_AGEMA_signal_2815, new_AGEMA_signal_2845, new_AGEMA_signal_2844,
         new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810,
         new_AGEMA_signal_2809, new_AGEMA_signal_2843, new_AGEMA_signal_2807,
         new_AGEMA_signal_2842, new_AGEMA_signal_2841, new_AGEMA_signal_2804,
         new_AGEMA_signal_2803, new_AGEMA_signal_2802, new_AGEMA_signal_2801,
         new_AGEMA_signal_2840, new_AGEMA_signal_2799, new_AGEMA_signal_2839,
         new_AGEMA_signal_2838, new_AGEMA_signal_2796, new_AGEMA_signal_2795,
         new_AGEMA_signal_2794, new_AGEMA_signal_2007, new_AGEMA_signal_2006,
         KeyArray_outS01ser_7_, new_AGEMA_signal_2009, new_AGEMA_signal_2008,
         KeyArray_outS01ser_6_, new_AGEMA_signal_2011, new_AGEMA_signal_2010,
         KeyArray_outS01ser_5_, new_AGEMA_signal_2013, new_AGEMA_signal_2012,
         KeyArray_outS01ser_4_, new_AGEMA_signal_2015, new_AGEMA_signal_2014,
         KeyArray_outS01ser_3_, new_AGEMA_signal_2017, new_AGEMA_signal_2016,
         KeyArray_outS01ser_2_, new_AGEMA_signal_2019, new_AGEMA_signal_2018,
         KeyArray_outS01ser_1_, new_AGEMA_signal_2021, new_AGEMA_signal_2020,
         KeyArray_outS01ser_0_, new_AGEMA_signal_3375,
         KeyArray_S00reg_gff_1_SFF_0_n5, new_AGEMA_signal_3267,
         KeyArray_S00reg_gff_1_SFF_0_QD, new_AGEMA_signal_2491,
         new_AGEMA_signal_3247, new_AGEMA_signal_3376,
         KeyArray_S00reg_gff_1_SFF_1_n6, new_AGEMA_signal_3268,
         KeyArray_S00reg_gff_1_SFF_1_QD, new_AGEMA_signal_2494,
         new_AGEMA_signal_3249, new_AGEMA_signal_3377,
         KeyArray_S00reg_gff_1_SFF_2_n6, new_AGEMA_signal_3269,
         KeyArray_S00reg_gff_1_SFF_2_QD, new_AGEMA_signal_2497,
         new_AGEMA_signal_3251, new_AGEMA_signal_3378,
         KeyArray_S00reg_gff_1_SFF_3_n6, new_AGEMA_signal_3270,
         KeyArray_S00reg_gff_1_SFF_3_QD, new_AGEMA_signal_2500,
         new_AGEMA_signal_3253, new_AGEMA_signal_3379,
         KeyArray_S00reg_gff_1_SFF_4_n6, new_AGEMA_signal_3271,
         KeyArray_S00reg_gff_1_SFF_4_QD, new_AGEMA_signal_2503,
         new_AGEMA_signal_3255, new_AGEMA_signal_3380,
         KeyArray_S00reg_gff_1_SFF_5_n6, new_AGEMA_signal_3272,
         KeyArray_S00reg_gff_1_SFF_5_QD, new_AGEMA_signal_2506,
         new_AGEMA_signal_3257, new_AGEMA_signal_3381,
         KeyArray_S00reg_gff_1_SFF_6_n6, new_AGEMA_signal_3273,
         KeyArray_S00reg_gff_1_SFF_6_QD, new_AGEMA_signal_2509,
         new_AGEMA_signal_3259, new_AGEMA_signal_3382,
         KeyArray_S00reg_gff_1_SFF_7_n6, new_AGEMA_signal_3274,
         KeyArray_S00reg_gff_1_SFF_7_QD, new_AGEMA_signal_2512,
         new_AGEMA_signal_3261, new_AGEMA_signal_3275,
         KeyArray_S01reg_gff_1_SFF_0_n6, new_AGEMA_signal_2888,
         KeyArray_S01reg_gff_1_SFF_0_QD, new_AGEMA_signal_2515,
         new_AGEMA_signal_2444, new_AGEMA_signal_3276,
         KeyArray_S01reg_gff_1_SFF_1_n6, new_AGEMA_signal_2889,
         KeyArray_S01reg_gff_1_SFF_1_QD, new_AGEMA_signal_2518,
         new_AGEMA_signal_2447, new_AGEMA_signal_3277,
         KeyArray_S01reg_gff_1_SFF_2_n6, new_AGEMA_signal_2890,
         KeyArray_S01reg_gff_1_SFF_2_QD, new_AGEMA_signal_2521,
         new_AGEMA_signal_2450, new_AGEMA_signal_3278,
         KeyArray_S01reg_gff_1_SFF_3_n6, new_AGEMA_signal_2891,
         KeyArray_S01reg_gff_1_SFF_3_QD, new_AGEMA_signal_2524,
         new_AGEMA_signal_2453, new_AGEMA_signal_3279,
         KeyArray_S01reg_gff_1_SFF_4_n6, new_AGEMA_signal_2892,
         KeyArray_S01reg_gff_1_SFF_4_QD, new_AGEMA_signal_2527,
         new_AGEMA_signal_2456, new_AGEMA_signal_3280,
         KeyArray_S01reg_gff_1_SFF_5_n6, new_AGEMA_signal_2893,
         KeyArray_S01reg_gff_1_SFF_5_QD, new_AGEMA_signal_2530,
         new_AGEMA_signal_2459, new_AGEMA_signal_3281,
         KeyArray_S01reg_gff_1_SFF_6_n6, new_AGEMA_signal_2894,
         KeyArray_S01reg_gff_1_SFF_6_QD, new_AGEMA_signal_2533,
         new_AGEMA_signal_2462, new_AGEMA_signal_3282,
         KeyArray_S01reg_gff_1_SFF_7_n6, new_AGEMA_signal_2895,
         KeyArray_S01reg_gff_1_SFF_7_QD, new_AGEMA_signal_2536,
         new_AGEMA_signal_2465, new_AGEMA_signal_3283,
         KeyArray_S02reg_gff_1_SFF_0_n6, new_AGEMA_signal_2896,
         KeyArray_S02reg_gff_1_SFF_0_QD, new_AGEMA_signal_2443,
         new_AGEMA_signal_2539, new_AGEMA_signal_2468, new_AGEMA_signal_3284,
         KeyArray_S02reg_gff_1_SFF_1_n6, new_AGEMA_signal_2897,
         KeyArray_S02reg_gff_1_SFF_1_QD, new_AGEMA_signal_2446,
         new_AGEMA_signal_2542, new_AGEMA_signal_2471, new_AGEMA_signal_3285,
         KeyArray_S02reg_gff_1_SFF_2_n6, new_AGEMA_signal_2898,
         KeyArray_S02reg_gff_1_SFF_2_QD, new_AGEMA_signal_2449,
         new_AGEMA_signal_2545, new_AGEMA_signal_2474, new_AGEMA_signal_3286,
         KeyArray_S02reg_gff_1_SFF_3_n6, new_AGEMA_signal_2899,
         KeyArray_S02reg_gff_1_SFF_3_QD, new_AGEMA_signal_2452,
         new_AGEMA_signal_2548, new_AGEMA_signal_2477, new_AGEMA_signal_3287,
         KeyArray_S02reg_gff_1_SFF_4_n6, new_AGEMA_signal_2900,
         KeyArray_S02reg_gff_1_SFF_4_QD, new_AGEMA_signal_2455,
         new_AGEMA_signal_2551, new_AGEMA_signal_2480, new_AGEMA_signal_3288,
         KeyArray_S02reg_gff_1_SFF_5_n6, new_AGEMA_signal_2901,
         KeyArray_S02reg_gff_1_SFF_5_QD, new_AGEMA_signal_2458,
         new_AGEMA_signal_2554, new_AGEMA_signal_2483, new_AGEMA_signal_3289,
         KeyArray_S02reg_gff_1_SFF_6_n6, new_AGEMA_signal_2902,
         KeyArray_S02reg_gff_1_SFF_6_QD, new_AGEMA_signal_2461,
         new_AGEMA_signal_2557, new_AGEMA_signal_2486, new_AGEMA_signal_3290,
         KeyArray_S02reg_gff_1_SFF_7_n6, new_AGEMA_signal_2903,
         KeyArray_S02reg_gff_1_SFF_7_QD, new_AGEMA_signal_2464,
         new_AGEMA_signal_2560, new_AGEMA_signal_2489, new_AGEMA_signal_3291,
         KeyArray_S03reg_gff_1_SFF_0_n6, new_AGEMA_signal_2904,
         KeyArray_S03reg_gff_1_SFF_0_QD, new_AGEMA_signal_2467,
         new_AGEMA_signal_2563, new_AGEMA_signal_2492, new_AGEMA_signal_3292,
         KeyArray_S03reg_gff_1_SFF_1_n6, new_AGEMA_signal_2905,
         KeyArray_S03reg_gff_1_SFF_1_QD, new_AGEMA_signal_2470,
         new_AGEMA_signal_2566, new_AGEMA_signal_2495, new_AGEMA_signal_3293,
         KeyArray_S03reg_gff_1_SFF_2_n6, new_AGEMA_signal_2906,
         KeyArray_S03reg_gff_1_SFF_2_QD, new_AGEMA_signal_2473,
         new_AGEMA_signal_2569, new_AGEMA_signal_2498, new_AGEMA_signal_3294,
         KeyArray_S03reg_gff_1_SFF_3_n6, new_AGEMA_signal_2907,
         KeyArray_S03reg_gff_1_SFF_3_QD, new_AGEMA_signal_2476,
         new_AGEMA_signal_2572, new_AGEMA_signal_2501, new_AGEMA_signal_3295,
         KeyArray_S03reg_gff_1_SFF_4_n6, new_AGEMA_signal_2908,
         KeyArray_S03reg_gff_1_SFF_4_QD, new_AGEMA_signal_2479,
         new_AGEMA_signal_2575, new_AGEMA_signal_2504, new_AGEMA_signal_3296,
         KeyArray_S03reg_gff_1_SFF_5_n5, new_AGEMA_signal_2909,
         KeyArray_S03reg_gff_1_SFF_5_QD, new_AGEMA_signal_2482,
         new_AGEMA_signal_2578, new_AGEMA_signal_2507, new_AGEMA_signal_3297,
         KeyArray_S03reg_gff_1_SFF_6_n5, new_AGEMA_signal_2910,
         KeyArray_S03reg_gff_1_SFF_6_QD, new_AGEMA_signal_2485,
         new_AGEMA_signal_2581, new_AGEMA_signal_2510, new_AGEMA_signal_3298,
         KeyArray_S03reg_gff_1_SFF_7_n5, new_AGEMA_signal_2911,
         KeyArray_S03reg_gff_1_SFF_7_QD, new_AGEMA_signal_2488,
         new_AGEMA_signal_2584, new_AGEMA_signal_2513, new_AGEMA_signal_3299,
         KeyArray_S10reg_gff_1_SFF_0_n5, new_AGEMA_signal_2912,
         KeyArray_S10reg_gff_1_SFF_0_QD, new_AGEMA_signal_2587,
         new_AGEMA_signal_2516, new_AGEMA_signal_3300,
         KeyArray_S10reg_gff_1_SFF_1_n5, new_AGEMA_signal_2913,
         KeyArray_S10reg_gff_1_SFF_1_QD, new_AGEMA_signal_2590,
         new_AGEMA_signal_2519, new_AGEMA_signal_3301,
         KeyArray_S10reg_gff_1_SFF_2_n5, new_AGEMA_signal_2914,
         KeyArray_S10reg_gff_1_SFF_2_QD, new_AGEMA_signal_2593,
         new_AGEMA_signal_2522, new_AGEMA_signal_3302,
         KeyArray_S10reg_gff_1_SFF_3_n5, new_AGEMA_signal_2915,
         KeyArray_S10reg_gff_1_SFF_3_QD, new_AGEMA_signal_2596,
         new_AGEMA_signal_2525, new_AGEMA_signal_3303,
         KeyArray_S10reg_gff_1_SFF_4_n5, new_AGEMA_signal_2916,
         KeyArray_S10reg_gff_1_SFF_4_QD, new_AGEMA_signal_2599,
         new_AGEMA_signal_2528, new_AGEMA_signal_3304,
         KeyArray_S10reg_gff_1_SFF_5_n5, new_AGEMA_signal_2917,
         KeyArray_S10reg_gff_1_SFF_5_QD, new_AGEMA_signal_2602,
         new_AGEMA_signal_2531, new_AGEMA_signal_3305,
         KeyArray_S10reg_gff_1_SFF_6_n5, new_AGEMA_signal_2918,
         KeyArray_S10reg_gff_1_SFF_6_QD, new_AGEMA_signal_2605,
         new_AGEMA_signal_2534, new_AGEMA_signal_3306,
         KeyArray_S10reg_gff_1_SFF_7_n5, new_AGEMA_signal_2919,
         KeyArray_S10reg_gff_1_SFF_7_QD, new_AGEMA_signal_2608,
         new_AGEMA_signal_2537, new_AGEMA_signal_3307,
         KeyArray_S11reg_gff_1_SFF_0_n6, new_AGEMA_signal_2920,
         KeyArray_S11reg_gff_1_SFF_0_QD, new_AGEMA_signal_2611,
         new_AGEMA_signal_2540, new_AGEMA_signal_3308,
         KeyArray_S11reg_gff_1_SFF_1_n6, new_AGEMA_signal_2921,
         KeyArray_S11reg_gff_1_SFF_1_QD, new_AGEMA_signal_2614,
         new_AGEMA_signal_2543, new_AGEMA_signal_3309,
         KeyArray_S11reg_gff_1_SFF_2_n6, new_AGEMA_signal_2922,
         KeyArray_S11reg_gff_1_SFF_2_QD, new_AGEMA_signal_2617,
         new_AGEMA_signal_2546, new_AGEMA_signal_3310,
         KeyArray_S11reg_gff_1_SFF_3_n6, new_AGEMA_signal_2923,
         KeyArray_S11reg_gff_1_SFF_3_QD, new_AGEMA_signal_2620,
         new_AGEMA_signal_2549, new_AGEMA_signal_3311,
         KeyArray_S11reg_gff_1_SFF_4_n6, new_AGEMA_signal_2924,
         KeyArray_S11reg_gff_1_SFF_4_QD, new_AGEMA_signal_2623,
         new_AGEMA_signal_2552, new_AGEMA_signal_3312,
         KeyArray_S11reg_gff_1_SFF_5_n6, new_AGEMA_signal_2925,
         KeyArray_S11reg_gff_1_SFF_5_QD, new_AGEMA_signal_2626,
         new_AGEMA_signal_2555, new_AGEMA_signal_3313,
         KeyArray_S11reg_gff_1_SFF_6_n6, new_AGEMA_signal_2926,
         KeyArray_S11reg_gff_1_SFF_6_QD, new_AGEMA_signal_2629,
         new_AGEMA_signal_2558, new_AGEMA_signal_3314,
         KeyArray_S11reg_gff_1_SFF_7_n6, new_AGEMA_signal_2927,
         KeyArray_S11reg_gff_1_SFF_7_QD, new_AGEMA_signal_2632,
         new_AGEMA_signal_2561, new_AGEMA_signal_3093,
         KeyArray_S12reg_gff_1_SFF_0_n6, new_AGEMA_signal_2928,
         KeyArray_S12reg_gff_1_SFF_0_QD, new_AGEMA_signal_2635,
         new_AGEMA_signal_2564, new_AGEMA_signal_3094,
         KeyArray_S12reg_gff_1_SFF_1_n6, new_AGEMA_signal_2929,
         KeyArray_S12reg_gff_1_SFF_1_QD, new_AGEMA_signal_2638,
         new_AGEMA_signal_2567, new_AGEMA_signal_3095,
         KeyArray_S12reg_gff_1_SFF_2_n6, new_AGEMA_signal_2930,
         KeyArray_S12reg_gff_1_SFF_2_QD, new_AGEMA_signal_2641,
         new_AGEMA_signal_2570, new_AGEMA_signal_3096,
         KeyArray_S12reg_gff_1_SFF_3_n6, new_AGEMA_signal_2931,
         KeyArray_S12reg_gff_1_SFF_3_QD, new_AGEMA_signal_2644,
         new_AGEMA_signal_2573, new_AGEMA_signal_3097,
         KeyArray_S12reg_gff_1_SFF_4_n6, new_AGEMA_signal_2932,
         KeyArray_S12reg_gff_1_SFF_4_QD, new_AGEMA_signal_2647,
         new_AGEMA_signal_2576, new_AGEMA_signal_3098,
         KeyArray_S12reg_gff_1_SFF_5_n6, new_AGEMA_signal_2933,
         KeyArray_S12reg_gff_1_SFF_5_QD, new_AGEMA_signal_2650,
         new_AGEMA_signal_2579, new_AGEMA_signal_3099,
         KeyArray_S12reg_gff_1_SFF_6_n6, new_AGEMA_signal_2934,
         KeyArray_S12reg_gff_1_SFF_6_QD, new_AGEMA_signal_2653,
         new_AGEMA_signal_2582, new_AGEMA_signal_3100,
         KeyArray_S12reg_gff_1_SFF_7_n6, new_AGEMA_signal_2935,
         KeyArray_S12reg_gff_1_SFF_7_QD, new_AGEMA_signal_2656,
         new_AGEMA_signal_2585, new_AGEMA_signal_3101,
         KeyArray_S13reg_gff_1_SFF_0_n6, new_AGEMA_signal_2936,
         KeyArray_S13reg_gff_1_SFF_0_QD, new_AGEMA_signal_2659,
         new_AGEMA_signal_2588, new_AGEMA_signal_3102,
         KeyArray_S13reg_gff_1_SFF_1_n6, new_AGEMA_signal_2937,
         KeyArray_S13reg_gff_1_SFF_1_QD, new_AGEMA_signal_2662,
         new_AGEMA_signal_2591, new_AGEMA_signal_3103,
         KeyArray_S13reg_gff_1_SFF_2_n6, new_AGEMA_signal_2938,
         KeyArray_S13reg_gff_1_SFF_2_QD, new_AGEMA_signal_2665,
         new_AGEMA_signal_2594, new_AGEMA_signal_3104,
         KeyArray_S13reg_gff_1_SFF_3_n6, new_AGEMA_signal_2939,
         KeyArray_S13reg_gff_1_SFF_3_QD, new_AGEMA_signal_2668,
         new_AGEMA_signal_2597, new_AGEMA_signal_3105,
         KeyArray_S13reg_gff_1_SFF_4_n6, new_AGEMA_signal_2940,
         KeyArray_S13reg_gff_1_SFF_4_QD, new_AGEMA_signal_2671,
         new_AGEMA_signal_2600, new_AGEMA_signal_3106,
         KeyArray_S13reg_gff_1_SFF_5_n5, new_AGEMA_signal_2941,
         KeyArray_S13reg_gff_1_SFF_5_QD, new_AGEMA_signal_2674,
         new_AGEMA_signal_2603, new_AGEMA_signal_3107,
         KeyArray_S13reg_gff_1_SFF_6_n5, new_AGEMA_signal_2942,
         KeyArray_S13reg_gff_1_SFF_6_QD, new_AGEMA_signal_2677,
         new_AGEMA_signal_2606, new_AGEMA_signal_3108,
         KeyArray_S13reg_gff_1_SFF_7_n5, new_AGEMA_signal_2943,
         KeyArray_S13reg_gff_1_SFF_7_QD, new_AGEMA_signal_2680,
         new_AGEMA_signal_2609, new_AGEMA_signal_3315,
         KeyArray_S20reg_gff_1_SFF_0_n5, new_AGEMA_signal_2944,
         KeyArray_S20reg_gff_1_SFF_0_QD, new_AGEMA_signal_2683,
         new_AGEMA_signal_2612, new_AGEMA_signal_3316,
         KeyArray_S20reg_gff_1_SFF_1_n5, new_AGEMA_signal_2945,
         KeyArray_S20reg_gff_1_SFF_1_QD, new_AGEMA_signal_2686,
         new_AGEMA_signal_2615, new_AGEMA_signal_3317,
         KeyArray_S20reg_gff_1_SFF_2_n5, new_AGEMA_signal_2946,
         KeyArray_S20reg_gff_1_SFF_2_QD, new_AGEMA_signal_2689,
         new_AGEMA_signal_2618, new_AGEMA_signal_3318,
         KeyArray_S20reg_gff_1_SFF_3_n5, new_AGEMA_signal_2947,
         KeyArray_S20reg_gff_1_SFF_3_QD, new_AGEMA_signal_2692,
         new_AGEMA_signal_2621, new_AGEMA_signal_3319,
         KeyArray_S20reg_gff_1_SFF_4_n5, new_AGEMA_signal_2948,
         KeyArray_S20reg_gff_1_SFF_4_QD, new_AGEMA_signal_2695,
         new_AGEMA_signal_2624, new_AGEMA_signal_3320,
         KeyArray_S20reg_gff_1_SFF_5_n5, new_AGEMA_signal_2949,
         KeyArray_S20reg_gff_1_SFF_5_QD, new_AGEMA_signal_2698,
         new_AGEMA_signal_2627, new_AGEMA_signal_3321,
         KeyArray_S20reg_gff_1_SFF_6_n5, new_AGEMA_signal_2950,
         KeyArray_S20reg_gff_1_SFF_6_QD, new_AGEMA_signal_2701,
         new_AGEMA_signal_2630, new_AGEMA_signal_3322,
         KeyArray_S20reg_gff_1_SFF_7_n5, new_AGEMA_signal_2951,
         KeyArray_S20reg_gff_1_SFF_7_QD, new_AGEMA_signal_2704,
         new_AGEMA_signal_2633, new_AGEMA_signal_3323,
         KeyArray_S21reg_gff_1_SFF_0_n6, new_AGEMA_signal_2952,
         KeyArray_S21reg_gff_1_SFF_0_QD, new_AGEMA_signal_2707,
         new_AGEMA_signal_2636, new_AGEMA_signal_3324,
         KeyArray_S21reg_gff_1_SFF_1_n6, new_AGEMA_signal_2953,
         KeyArray_S21reg_gff_1_SFF_1_QD, new_AGEMA_signal_2710,
         new_AGEMA_signal_2639, new_AGEMA_signal_3325,
         KeyArray_S21reg_gff_1_SFF_2_n6, new_AGEMA_signal_2954,
         KeyArray_S21reg_gff_1_SFF_2_QD, new_AGEMA_signal_2713,
         new_AGEMA_signal_2642, new_AGEMA_signal_3326,
         KeyArray_S21reg_gff_1_SFF_3_n6, new_AGEMA_signal_2955,
         KeyArray_S21reg_gff_1_SFF_3_QD, new_AGEMA_signal_2716,
         new_AGEMA_signal_2645, new_AGEMA_signal_3327,
         KeyArray_S21reg_gff_1_SFF_4_n6, new_AGEMA_signal_2956,
         KeyArray_S21reg_gff_1_SFF_4_QD, new_AGEMA_signal_2719,
         new_AGEMA_signal_2648, new_AGEMA_signal_3328,
         KeyArray_S21reg_gff_1_SFF_5_n6, new_AGEMA_signal_2957,
         KeyArray_S21reg_gff_1_SFF_5_QD, new_AGEMA_signal_2722,
         new_AGEMA_signal_2651, new_AGEMA_signal_3329,
         KeyArray_S21reg_gff_1_SFF_6_n6, new_AGEMA_signal_2958,
         KeyArray_S21reg_gff_1_SFF_6_QD, new_AGEMA_signal_2725,
         new_AGEMA_signal_2654, new_AGEMA_signal_3330,
         KeyArray_S21reg_gff_1_SFF_7_n6, new_AGEMA_signal_2959,
         KeyArray_S21reg_gff_1_SFF_7_QD, new_AGEMA_signal_2728,
         new_AGEMA_signal_2657, new_AGEMA_signal_3331,
         KeyArray_S22reg_gff_1_SFF_0_n6, new_AGEMA_signal_2960,
         KeyArray_S22reg_gff_1_SFF_0_QD, new_AGEMA_signal_2731,
         new_AGEMA_signal_2660, new_AGEMA_signal_3332,
         KeyArray_S22reg_gff_1_SFF_1_n6, new_AGEMA_signal_2961,
         KeyArray_S22reg_gff_1_SFF_1_QD, new_AGEMA_signal_2734,
         new_AGEMA_signal_2663, new_AGEMA_signal_3333,
         KeyArray_S22reg_gff_1_SFF_2_n6, new_AGEMA_signal_2962,
         KeyArray_S22reg_gff_1_SFF_2_QD, new_AGEMA_signal_2737,
         new_AGEMA_signal_2666, new_AGEMA_signal_3334,
         KeyArray_S22reg_gff_1_SFF_3_n6, new_AGEMA_signal_2963,
         KeyArray_S22reg_gff_1_SFF_3_QD, new_AGEMA_signal_2740,
         new_AGEMA_signal_2669, new_AGEMA_signal_3335,
         KeyArray_S22reg_gff_1_SFF_4_n6, new_AGEMA_signal_2964,
         KeyArray_S22reg_gff_1_SFF_4_QD, new_AGEMA_signal_2743,
         new_AGEMA_signal_2672, new_AGEMA_signal_3336,
         KeyArray_S22reg_gff_1_SFF_5_n6, new_AGEMA_signal_2965,
         KeyArray_S22reg_gff_1_SFF_5_QD, new_AGEMA_signal_2746,
         new_AGEMA_signal_2675, new_AGEMA_signal_3337,
         KeyArray_S22reg_gff_1_SFF_6_n6, new_AGEMA_signal_2966,
         KeyArray_S22reg_gff_1_SFF_6_QD, new_AGEMA_signal_2749,
         new_AGEMA_signal_2678, new_AGEMA_signal_3338,
         KeyArray_S22reg_gff_1_SFF_7_n6, new_AGEMA_signal_2967,
         KeyArray_S22reg_gff_1_SFF_7_QD, new_AGEMA_signal_2752,
         new_AGEMA_signal_2681, new_AGEMA_signal_3339,
         KeyArray_S23reg_gff_1_SFF_0_n6, new_AGEMA_signal_2968,
         KeyArray_S23reg_gff_1_SFF_0_QD, new_AGEMA_signal_2755,
         new_AGEMA_signal_2684, new_AGEMA_signal_3340,
         KeyArray_S23reg_gff_1_SFF_1_n6, new_AGEMA_signal_2969,
         KeyArray_S23reg_gff_1_SFF_1_QD, new_AGEMA_signal_2758,
         new_AGEMA_signal_2687, new_AGEMA_signal_3341,
         KeyArray_S23reg_gff_1_SFF_2_n6, new_AGEMA_signal_2970,
         KeyArray_S23reg_gff_1_SFF_2_QD, new_AGEMA_signal_2761,
         new_AGEMA_signal_2690, new_AGEMA_signal_3342,
         KeyArray_S23reg_gff_1_SFF_3_n6, new_AGEMA_signal_2971,
         KeyArray_S23reg_gff_1_SFF_3_QD, new_AGEMA_signal_2764,
         new_AGEMA_signal_2693, new_AGEMA_signal_3343,
         KeyArray_S23reg_gff_1_SFF_4_n6, new_AGEMA_signal_2972,
         KeyArray_S23reg_gff_1_SFF_4_QD, new_AGEMA_signal_2767,
         new_AGEMA_signal_2696, new_AGEMA_signal_3344,
         KeyArray_S23reg_gff_1_SFF_5_n5, new_AGEMA_signal_2973,
         KeyArray_S23reg_gff_1_SFF_5_QD, new_AGEMA_signal_2770,
         new_AGEMA_signal_2699, new_AGEMA_signal_3345,
         KeyArray_S23reg_gff_1_SFF_6_n5, new_AGEMA_signal_2974,
         KeyArray_S23reg_gff_1_SFF_6_QD, new_AGEMA_signal_2773,
         new_AGEMA_signal_2702, new_AGEMA_signal_3346,
         KeyArray_S23reg_gff_1_SFF_7_n5, new_AGEMA_signal_2975,
         KeyArray_S23reg_gff_1_SFF_7_QD, new_AGEMA_signal_2776,
         new_AGEMA_signal_2705, new_AGEMA_signal_3347,
         KeyArray_S31reg_gff_1_SFF_0_n6, new_AGEMA_signal_2976,
         KeyArray_S31reg_gff_1_SFF_0_QD, new_AGEMA_signal_2732,
         new_AGEMA_signal_3348, KeyArray_S31reg_gff_1_SFF_1_n6,
         new_AGEMA_signal_2977, KeyArray_S31reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2735, new_AGEMA_signal_3349,
         KeyArray_S31reg_gff_1_SFF_2_n6, new_AGEMA_signal_2978,
         KeyArray_S31reg_gff_1_SFF_2_QD, new_AGEMA_signal_2738,
         new_AGEMA_signal_3350, KeyArray_S31reg_gff_1_SFF_3_n6,
         new_AGEMA_signal_2979, KeyArray_S31reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2741, new_AGEMA_signal_3351,
         KeyArray_S31reg_gff_1_SFF_4_n6, new_AGEMA_signal_2980,
         KeyArray_S31reg_gff_1_SFF_4_QD, new_AGEMA_signal_2744,
         new_AGEMA_signal_3352, KeyArray_S31reg_gff_1_SFF_5_n6,
         new_AGEMA_signal_2981, KeyArray_S31reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2747, new_AGEMA_signal_3353,
         KeyArray_S31reg_gff_1_SFF_6_n6, new_AGEMA_signal_2982,
         KeyArray_S31reg_gff_1_SFF_6_QD, new_AGEMA_signal_2750,
         new_AGEMA_signal_3354, KeyArray_S31reg_gff_1_SFF_7_n6,
         new_AGEMA_signal_2983, KeyArray_S31reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2753, new_AGEMA_signal_3355,
         KeyArray_S32reg_gff_1_SFF_0_n6, new_AGEMA_signal_2984,
         KeyArray_S32reg_gff_1_SFF_0_QD, new_AGEMA_signal_2756,
         new_AGEMA_signal_3356, KeyArray_S32reg_gff_1_SFF_1_n6,
         new_AGEMA_signal_2985, KeyArray_S32reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2759, new_AGEMA_signal_3357,
         KeyArray_S32reg_gff_1_SFF_2_n6, new_AGEMA_signal_2986,
         KeyArray_S32reg_gff_1_SFF_2_QD, new_AGEMA_signal_2762,
         new_AGEMA_signal_3358, KeyArray_S32reg_gff_1_SFF_3_n6,
         new_AGEMA_signal_2987, KeyArray_S32reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2765, new_AGEMA_signal_3359,
         KeyArray_S32reg_gff_1_SFF_4_n6, new_AGEMA_signal_2988,
         KeyArray_S32reg_gff_1_SFF_4_QD, new_AGEMA_signal_2768,
         new_AGEMA_signal_3360, KeyArray_S32reg_gff_1_SFF_5_n6,
         new_AGEMA_signal_2989, KeyArray_S32reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2771, new_AGEMA_signal_3361,
         KeyArray_S32reg_gff_1_SFF_6_n5, new_AGEMA_signal_2990,
         KeyArray_S32reg_gff_1_SFF_6_QD, new_AGEMA_signal_2774,
         new_AGEMA_signal_3362, KeyArray_S32reg_gff_1_SFF_7_n5,
         new_AGEMA_signal_2991, KeyArray_S32reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2777, new_AGEMA_signal_3363,
         KeyArray_S33reg_gff_1_SFF_0_n5, new_AGEMA_signal_2992,
         KeyArray_S33reg_gff_1_SFF_0_QD, new_AGEMA_signal_2779,
         new_AGEMA_signal_3364, KeyArray_S33reg_gff_1_SFF_1_n5,
         new_AGEMA_signal_2993, KeyArray_S33reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2781, new_AGEMA_signal_3365,
         KeyArray_S33reg_gff_1_SFF_2_n5, new_AGEMA_signal_2994,
         KeyArray_S33reg_gff_1_SFF_2_QD, new_AGEMA_signal_2783,
         new_AGEMA_signal_3366, KeyArray_S33reg_gff_1_SFF_3_n5,
         new_AGEMA_signal_2995, KeyArray_S33reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2785, new_AGEMA_signal_3367,
         KeyArray_S33reg_gff_1_SFF_4_n5, new_AGEMA_signal_2996,
         KeyArray_S33reg_gff_1_SFF_4_QD, new_AGEMA_signal_2787,
         new_AGEMA_signal_3368, KeyArray_S33reg_gff_1_SFF_5_n5,
         new_AGEMA_signal_2997, KeyArray_S33reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2789, new_AGEMA_signal_3369,
         KeyArray_S33reg_gff_1_SFF_6_n5, new_AGEMA_signal_2998,
         KeyArray_S33reg_gff_1_SFF_6_QD, new_AGEMA_signal_2791,
         new_AGEMA_signal_3370, KeyArray_S33reg_gff_1_SFF_7_n5,
         new_AGEMA_signal_2999, KeyArray_S33reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2793, new_AGEMA_signal_3109, new_AGEMA_signal_3110,
         new_AGEMA_signal_3111, new_AGEMA_signal_3112, new_AGEMA_signal_3113,
         new_AGEMA_signal_3114, new_AGEMA_signal_3115, new_AGEMA_signal_3116,
         new_AGEMA_signal_2708, new_AGEMA_signal_2711, new_AGEMA_signal_2714,
         new_AGEMA_signal_2717, new_AGEMA_signal_2720, new_AGEMA_signal_2723,
         new_AGEMA_signal_2726, new_AGEMA_signal_2729, new_AGEMA_signal_2024,
         MixColumns_line0_n15, new_AGEMA_signal_2122, MixColumns_line0_n16,
         new_AGEMA_signal_2051, new_AGEMA_signal_2027, MixColumns_line0_n13,
         new_AGEMA_signal_2123, MixColumns_line0_n14, new_AGEMA_signal_2053,
         new_AGEMA_signal_2030, MixColumns_line0_n11, new_AGEMA_signal_2124,
         MixColumns_line0_n12, new_AGEMA_signal_2055, new_AGEMA_signal_2033,
         MixColumns_line0_n9, new_AGEMA_signal_2797, MixColumns_line0_n10,
         new_AGEMA_signal_2127, MixColumns_line0_S02_1, new_AGEMA_signal_2046,
         new_AGEMA_signal_2036, MixColumns_line0_n7, new_AGEMA_signal_2798,
         MixColumns_line0_n8, new_AGEMA_signal_2128, new_AGEMA_signal_2047,
         new_AGEMA_signal_2039, MixColumns_line0_n5, new_AGEMA_signal_2125,
         MixColumns_line0_n6, new_AGEMA_signal_2058, new_AGEMA_signal_2042,
         MixColumns_line0_n3, new_AGEMA_signal_2800, MixColumns_line0_n4,
         new_AGEMA_signal_2129, new_AGEMA_signal_2048, new_AGEMA_signal_2045,
         MixColumns_line0_n1, new_AGEMA_signal_2126, MixColumns_line0_n2,
         new_AGEMA_signal_2060, MixColumns_line0_timesTHREE_input2_1,
         new_AGEMA_signal_2062, new_AGEMA_signal_2063, new_AGEMA_signal_2064,
         new_AGEMA_signal_2065, MixColumns_line1_n15, new_AGEMA_signal_2130,
         MixColumns_line1_n16, new_AGEMA_signal_2076, new_AGEMA_signal_2066,
         MixColumns_line1_n13, new_AGEMA_signal_2131, MixColumns_line1_n14,
         new_AGEMA_signal_2077, new_AGEMA_signal_2067, MixColumns_line1_n11,
         new_AGEMA_signal_2132, MixColumns_line1_n12, new_AGEMA_signal_2078,
         new_AGEMA_signal_2068, MixColumns_line1_n9, new_AGEMA_signal_2805,
         MixColumns_line1_n10, new_AGEMA_signal_2135, new_AGEMA_signal_2073,
         MixColumns_line1_S02_4_, new_AGEMA_signal_2069, MixColumns_line1_n7,
         new_AGEMA_signal_2806, MixColumns_line1_n8, new_AGEMA_signal_2136,
         new_AGEMA_signal_2074, MixColumns_line1_S02_3_, new_AGEMA_signal_2070,
         MixColumns_line1_n5, new_AGEMA_signal_2133, MixColumns_line1_n6,
         new_AGEMA_signal_2079, new_AGEMA_signal_2071, MixColumns_line1_n3,
         new_AGEMA_signal_2808, MixColumns_line1_n4, new_AGEMA_signal_2137,
         new_AGEMA_signal_2075, MixColumns_line1_S02_1_, new_AGEMA_signal_2072,
         MixColumns_line1_n1, new_AGEMA_signal_2134, MixColumns_line1_n2,
         new_AGEMA_signal_2080, MixColumns_line1_timesTHREE_input2_1,
         new_AGEMA_signal_2081, new_AGEMA_signal_2082, new_AGEMA_signal_2083,
         new_AGEMA_signal_2084, MixColumns_line2_n15, new_AGEMA_signal_2138,
         MixColumns_line2_n16, new_AGEMA_signal_2095, new_AGEMA_signal_2085,
         MixColumns_line2_n13, new_AGEMA_signal_2139, MixColumns_line2_n14,
         new_AGEMA_signal_2096, new_AGEMA_signal_2086, MixColumns_line2_n11,
         new_AGEMA_signal_2140, MixColumns_line2_n12, new_AGEMA_signal_2097,
         new_AGEMA_signal_2087, MixColumns_line2_n9, new_AGEMA_signal_2813,
         MixColumns_line2_n10, new_AGEMA_signal_2143, new_AGEMA_signal_2092,
         MixColumns_line2_S02_4_, new_AGEMA_signal_2088, MixColumns_line2_n7,
         new_AGEMA_signal_2814, MixColumns_line2_n8, new_AGEMA_signal_2144,
         new_AGEMA_signal_2093, MixColumns_line2_S02_3_, new_AGEMA_signal_2089,
         MixColumns_line2_n5, new_AGEMA_signal_2141, MixColumns_line2_n6,
         new_AGEMA_signal_2098, new_AGEMA_signal_2090, MixColumns_line2_n3,
         new_AGEMA_signal_2816, MixColumns_line2_n4, new_AGEMA_signal_2145,
         new_AGEMA_signal_2094, MixColumns_line2_S02_1_, new_AGEMA_signal_2091,
         MixColumns_line2_n1, new_AGEMA_signal_2142, MixColumns_line2_n2,
         new_AGEMA_signal_2099, MixColumns_line2_timesTHREE_input2_1,
         new_AGEMA_signal_2100, new_AGEMA_signal_2101, new_AGEMA_signal_2102,
         new_AGEMA_signal_2103, MixColumns_line3_n15, new_AGEMA_signal_2146,
         MixColumns_line3_n16, new_AGEMA_signal_2114, new_AGEMA_signal_2104,
         MixColumns_line3_n13, new_AGEMA_signal_2147, MixColumns_line3_n14,
         new_AGEMA_signal_2115, new_AGEMA_signal_2105, MixColumns_line3_n11,
         new_AGEMA_signal_2148, MixColumns_line3_n12, new_AGEMA_signal_2116,
         new_AGEMA_signal_2106, MixColumns_line3_n9, new_AGEMA_signal_2821,
         MixColumns_line3_n10, new_AGEMA_signal_2151, new_AGEMA_signal_2111,
         MixColumns_line3_S02_4_, new_AGEMA_signal_2107, MixColumns_line3_n7,
         new_AGEMA_signal_2822, MixColumns_line3_n8, new_AGEMA_signal_2152,
         new_AGEMA_signal_2112, MixColumns_line3_S02_3_, new_AGEMA_signal_2108,
         MixColumns_line3_n5, new_AGEMA_signal_2149, MixColumns_line3_n6,
         new_AGEMA_signal_2117, new_AGEMA_signal_2109, MixColumns_line3_n3,
         new_AGEMA_signal_2824, MixColumns_line3_n4, new_AGEMA_signal_2153,
         new_AGEMA_signal_2113, MixColumns_line3_S02_1_, new_AGEMA_signal_2110,
         MixColumns_line3_n1, new_AGEMA_signal_2150, MixColumns_line3_n2,
         new_AGEMA_signal_2118, new_AGEMA_signal_2119,
         MixColumns_line3_timesTHREE_input2_4_, new_AGEMA_signal_2120,
         MixColumns_line3_timesTHREE_input2_3_, new_AGEMA_signal_2121,
         MixColumns_line3_timesTHREE_input2_1_, calcRCon_n51, calcRCon_n50,
         calcRCon_n49, calcRCon_n48, calcRCon_n47, calcRCon_n46, calcRCon_n45,
         calcRCon_n44, new_AGEMA_signal_2826, new_AGEMA_signal_2827,
         new_AGEMA_signal_2828, new_AGEMA_signal_2829, new_AGEMA_signal_2830,
         new_AGEMA_signal_2831, new_AGEMA_signal_2832, new_AGEMA_signal_2833,
         new_AGEMA_signal_2850, Inst_bSbox_T1, new_AGEMA_signal_2851,
         Inst_bSbox_T2, new_AGEMA_signal_2852, Inst_bSbox_T3,
         new_AGEMA_signal_2853, Inst_bSbox_T4, new_AGEMA_signal_2854,
         Inst_bSbox_T5, new_AGEMA_signal_3000, Inst_bSbox_T6,
         new_AGEMA_signal_2855, Inst_bSbox_T7, new_AGEMA_signal_3032,
         Inst_bSbox_T8, new_AGEMA_signal_3001, Inst_bSbox_T9,
         new_AGEMA_signal_3033, Inst_bSbox_T10, new_AGEMA_signal_2856,
         Inst_bSbox_T11, new_AGEMA_signal_2857, Inst_bSbox_T12,
         new_AGEMA_signal_3002, Inst_bSbox_T13, new_AGEMA_signal_3034,
         Inst_bSbox_T14, new_AGEMA_signal_3003, Inst_bSbox_T15,
         new_AGEMA_signal_3004, Inst_bSbox_T16, new_AGEMA_signal_3035,
         Inst_bSbox_T17, new_AGEMA_signal_2858, Inst_bSbox_T18,
         new_AGEMA_signal_3005, Inst_bSbox_T19, new_AGEMA_signal_3036,
         Inst_bSbox_T20, new_AGEMA_signal_2859, Inst_bSbox_T21,
         new_AGEMA_signal_3006, Inst_bSbox_T22, new_AGEMA_signal_3037,
         Inst_bSbox_T23, new_AGEMA_signal_3117, Inst_bSbox_T24,
         new_AGEMA_signal_3118, Inst_bSbox_T25, new_AGEMA_signal_3038,
         Inst_bSbox_T26, new_AGEMA_signal_3007, Inst_bSbox_T27,
         new_AGEMA_signal_3039, Inst_bSbox_M1, new_AGEMA_signal_3119,
         Inst_bSbox_M2, new_AGEMA_signal_3120, Inst_bSbox_M3,
         new_AGEMA_signal_3603, new_AGEMA_signal_3602, new_AGEMA_signal_3040,
         Inst_bSbox_M4, new_AGEMA_signal_3121, Inst_bSbox_M5,
         new_AGEMA_signal_3041, Inst_bSbox_M6, new_AGEMA_signal_3042,
         Inst_bSbox_M7, new_AGEMA_signal_3122, Inst_bSbox_M8,
         new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3123,
         Inst_bSbox_M9, new_AGEMA_signal_3262, Inst_bSbox_M10,
         new_AGEMA_signal_3043, Inst_bSbox_M11, new_AGEMA_signal_3044,
         Inst_bSbox_M12, new_AGEMA_signal_3124, Inst_bSbox_M13,
         new_AGEMA_signal_3125, Inst_bSbox_M14, new_AGEMA_signal_3263,
         Inst_bSbox_M15, new_AGEMA_signal_3264, Inst_bSbox_M16,
         new_AGEMA_signal_3265, Inst_bSbox_M17, new_AGEMA_signal_3607,
         new_AGEMA_signal_3606, new_AGEMA_signal_3266, Inst_bSbox_M18,
         new_AGEMA_signal_3371, Inst_bSbox_M19, new_AGEMA_signal_3372,
         Inst_bSbox_M20, new_AGEMA_signal_3373, Inst_bSbox_M21,
         new_AGEMA_signal_3374, Inst_bSbox_M22, new_AGEMA_signal_3383,
         Inst_bSbox_M23, new_AGEMA_signal_3609, new_AGEMA_signal_3608,
         new_AGEMA_signal_3387, Inst_bSbox_M24, new_AGEMA_signal_3385,
         Inst_bSbox_M27, new_AGEMA_signal_3626, new_AGEMA_signal_3630,
         new_AGEMA_signal_3634, new_AGEMA_signal_3638, new_AGEMA_signal_3642,
         new_AGEMA_signal_3646, new_AGEMA_signal_3650, new_AGEMA_signal_3654,
         new_AGEMA_signal_3658, new_AGEMA_signal_3662, new_AGEMA_signal_3666,
         new_AGEMA_signal_3670, new_AGEMA_signal_3674, new_AGEMA_signal_3678,
         new_AGEMA_signal_3682, new_AGEMA_signal_3686, new_AGEMA_signal_3690,
         new_AGEMA_signal_3694, new_AGEMA_signal_3698, new_AGEMA_signal_3702,
         new_AGEMA_signal_3706, new_AGEMA_signal_3710, new_AGEMA_signal_3714,
         new_AGEMA_signal_3718, new_AGEMA_signal_3722, new_AGEMA_signal_3726,
         new_AGEMA_signal_3730, new_AGEMA_signal_3734, new_AGEMA_signal_3738,
         new_AGEMA_signal_3742, new_AGEMA_signal_3746, new_AGEMA_signal_3750,
         new_AGEMA_signal_3754, new_AGEMA_signal_3758, new_AGEMA_signal_3762,
         new_AGEMA_signal_3766, new_AGEMA_signal_3770, new_AGEMA_signal_3774,
         new_AGEMA_signal_3778, new_AGEMA_signal_3782, new_AGEMA_signal_3786,
         new_AGEMA_signal_3790, new_AGEMA_signal_3794, new_AGEMA_signal_3798,
         new_AGEMA_signal_3802, new_AGEMA_signal_3806, new_AGEMA_signal_3810,
         new_AGEMA_signal_3814, new_AGEMA_signal_3818, new_AGEMA_signal_3822,
         new_AGEMA_signal_3826, new_AGEMA_signal_3830, new_AGEMA_signal_3834,
         new_AGEMA_signal_3838, new_AGEMA_signal_3842, new_AGEMA_signal_3846,
         new_AGEMA_signal_3850, new_AGEMA_signal_3854, new_AGEMA_signal_3858,
         new_AGEMA_signal_3862, new_AGEMA_signal_3866, new_AGEMA_signal_3870,
         new_AGEMA_signal_3874, new_AGEMA_signal_3878, new_AGEMA_signal_3882,
         new_AGEMA_signal_3886, new_AGEMA_signal_3890, new_AGEMA_signal_3894,
         new_AGEMA_signal_3898, new_AGEMA_signal_3902, new_AGEMA_signal_3906,
         new_AGEMA_signal_3910, new_AGEMA_signal_3914, new_AGEMA_signal_3918,
         new_AGEMA_signal_3922, new_AGEMA_signal_3926, new_AGEMA_signal_3930,
         new_AGEMA_signal_3934, new_AGEMA_signal_3938, new_AGEMA_signal_3942,
         new_AGEMA_signal_3946, new_AGEMA_signal_3950, new_AGEMA_signal_3954,
         new_AGEMA_signal_3958, new_AGEMA_signal_3962, new_AGEMA_signal_3966,
         new_AGEMA_signal_3970, new_AGEMA_signal_3974, new_AGEMA_signal_3978,
         new_AGEMA_signal_3982, new_AGEMA_signal_3986, new_AGEMA_signal_3990,
         new_AGEMA_signal_3994, new_AGEMA_signal_3998, new_AGEMA_signal_4002,
         new_AGEMA_signal_4006, new_AGEMA_signal_4010, new_AGEMA_signal_4014,
         new_AGEMA_signal_4018, new_AGEMA_signal_4022, new_AGEMA_signal_4026,
         new_AGEMA_signal_4030, new_AGEMA_signal_4034, new_AGEMA_signal_4038,
         new_AGEMA_signal_4042, new_AGEMA_signal_4046, new_AGEMA_signal_4050,
         new_AGEMA_signal_4054, new_AGEMA_signal_4058, new_AGEMA_signal_4062,
         new_AGEMA_signal_4066, new_AGEMA_signal_4070, new_AGEMA_signal_4074,
         new_AGEMA_signal_4078, new_AGEMA_signal_4082, new_AGEMA_signal_4086,
         new_AGEMA_signal_4090, new_AGEMA_signal_4094, new_AGEMA_signal_4098,
         new_AGEMA_signal_4102, new_AGEMA_signal_4106, new_AGEMA_signal_4110,
         new_AGEMA_signal_4114, new_AGEMA_signal_4118, new_AGEMA_signal_4122,
         new_AGEMA_signal_4126, new_AGEMA_signal_4130, new_AGEMA_signal_4133,
         new_AGEMA_signal_4136, new_AGEMA_signal_4139, new_AGEMA_signal_4142,
         new_AGEMA_signal_4145, new_AGEMA_signal_4148, new_AGEMA_signal_4151,
         new_AGEMA_signal_4154, new_AGEMA_signal_4157, new_AGEMA_signal_4160,
         new_AGEMA_signal_4163, new_AGEMA_signal_4166, new_AGEMA_signal_4169,
         new_AGEMA_signal_4172, new_AGEMA_signal_4175, new_AGEMA_signal_4178,
         new_AGEMA_signal_4181, new_AGEMA_signal_4184, new_AGEMA_signal_4187,
         new_AGEMA_signal_4190, new_AGEMA_signal_4193, new_AGEMA_signal_4196,
         new_AGEMA_signal_4199, new_AGEMA_signal_4202, new_AGEMA_signal_4205,
         new_AGEMA_signal_4208, new_AGEMA_signal_4211, new_AGEMA_signal_4214,
         new_AGEMA_signal_4217, new_AGEMA_signal_4220, new_AGEMA_signal_4223,
         new_AGEMA_signal_4226, new_AGEMA_signal_4229, new_AGEMA_signal_4232,
         new_AGEMA_signal_4235, new_AGEMA_signal_4238, new_AGEMA_signal_4242,
         new_AGEMA_signal_4246, new_AGEMA_signal_4250, new_AGEMA_signal_4254,
         new_AGEMA_signal_4258, new_AGEMA_signal_4262, new_AGEMA_signal_4266,
         new_AGEMA_signal_4270, new_AGEMA_signal_4274, new_AGEMA_signal_4278,
         new_AGEMA_signal_4282, new_AGEMA_signal_4286, new_AGEMA_signal_4290,
         new_AGEMA_signal_4294, new_AGEMA_signal_4298, new_AGEMA_signal_4302,
         new_AGEMA_signal_4306, new_AGEMA_signal_4310, new_AGEMA_signal_4314,
         new_AGEMA_signal_4318, new_AGEMA_signal_4322, new_AGEMA_signal_4326,
         new_AGEMA_signal_4330, new_AGEMA_signal_4334, new_AGEMA_signal_4338,
         new_AGEMA_signal_4342, new_AGEMA_signal_4346, new_AGEMA_signal_4350,
         new_AGEMA_signal_4354, new_AGEMA_signal_4358, new_AGEMA_signal_4362,
         new_AGEMA_signal_4366, new_AGEMA_signal_4370, new_AGEMA_signal_4374,
         new_AGEMA_signal_4378, new_AGEMA_signal_4382, new_AGEMA_signal_4386,
         new_AGEMA_signal_4390, new_AGEMA_signal_4394, new_AGEMA_signal_4398,
         new_AGEMA_signal_4402, new_AGEMA_signal_4406, new_AGEMA_signal_4410,
         new_AGEMA_signal_4414, new_AGEMA_signal_4418, new_AGEMA_signal_4422,
         new_AGEMA_signal_4426, new_AGEMA_signal_4430, new_AGEMA_signal_4434,
         new_AGEMA_signal_4438, new_AGEMA_signal_4442, new_AGEMA_signal_4446,
         new_AGEMA_signal_4450, new_AGEMA_signal_4454, new_AGEMA_signal_4458,
         new_AGEMA_signal_4462, new_AGEMA_signal_4466, new_AGEMA_signal_4470,
         new_AGEMA_signal_4474, new_AGEMA_signal_4478, new_AGEMA_signal_4482,
         new_AGEMA_signal_4486, new_AGEMA_signal_4490, new_AGEMA_signal_4494,
         new_AGEMA_signal_4498, new_AGEMA_signal_4502, new_AGEMA_signal_4506,
         new_AGEMA_signal_4510, new_AGEMA_signal_4514, new_AGEMA_signal_4518,
         new_AGEMA_signal_4522, new_AGEMA_signal_4526, new_AGEMA_signal_4530,
         new_AGEMA_signal_4534, new_AGEMA_signal_4538, new_AGEMA_signal_4542,
         new_AGEMA_signal_4546, new_AGEMA_signal_4550, new_AGEMA_signal_4554,
         new_AGEMA_signal_4558, new_AGEMA_signal_4562, new_AGEMA_signal_4566,
         new_AGEMA_signal_4570, new_AGEMA_signal_4574, new_AGEMA_signal_4578,
         new_AGEMA_signal_4582, new_AGEMA_signal_4586, new_AGEMA_signal_4590,
         new_AGEMA_signal_4594, new_AGEMA_signal_4598, new_AGEMA_signal_4602,
         new_AGEMA_signal_4606, new_AGEMA_signal_4610, new_AGEMA_signal_4614,
         new_AGEMA_signal_4618, new_AGEMA_signal_4622, new_AGEMA_signal_4626,
         new_AGEMA_signal_4630, new_AGEMA_signal_4634, new_AGEMA_signal_4638,
         new_AGEMA_signal_4642, new_AGEMA_signal_4646, new_AGEMA_signal_4650,
         new_AGEMA_signal_4654, new_AGEMA_signal_4658, new_AGEMA_signal_4662,
         new_AGEMA_signal_4666, new_AGEMA_signal_4670, new_AGEMA_signal_4674,
         new_AGEMA_signal_4678, new_AGEMA_signal_4682, new_AGEMA_signal_4686,
         new_AGEMA_signal_4690, new_AGEMA_signal_4694, new_AGEMA_signal_4698,
         new_AGEMA_signal_4702, new_AGEMA_signal_4706, new_AGEMA_signal_4710,
         new_AGEMA_signal_4714, new_AGEMA_signal_4718, new_AGEMA_signal_4722,
         new_AGEMA_signal_4726, new_AGEMA_signal_4730, new_AGEMA_signal_4734,
         new_AGEMA_signal_4738, new_AGEMA_signal_4742, new_AGEMA_signal_4746,
         new_AGEMA_signal_4750, new_AGEMA_signal_4754, new_AGEMA_signal_4758,
         new_AGEMA_signal_4762, new_AGEMA_signal_4766, new_AGEMA_signal_4770,
         new_AGEMA_signal_4774, new_AGEMA_signal_4778, new_AGEMA_signal_4782,
         new_AGEMA_signal_4786, new_AGEMA_signal_4790, new_AGEMA_signal_4794,
         new_AGEMA_signal_4798, new_AGEMA_signal_4802, new_AGEMA_signal_4806,
         new_AGEMA_signal_4810, new_AGEMA_signal_4814, new_AGEMA_signal_4818,
         new_AGEMA_signal_4822, new_AGEMA_signal_4826, new_AGEMA_signal_4830,
         new_AGEMA_signal_4834, new_AGEMA_signal_4838, new_AGEMA_signal_4842,
         new_AGEMA_signal_4846, new_AGEMA_signal_4850, new_AGEMA_signal_4854,
         new_AGEMA_signal_4858, new_AGEMA_signal_4862, new_AGEMA_signal_4866,
         new_AGEMA_signal_4870, new_AGEMA_signal_4874, new_AGEMA_signal_4878,
         new_AGEMA_signal_4882, new_AGEMA_signal_4886, new_AGEMA_signal_4890,
         new_AGEMA_signal_4894, new_AGEMA_signal_4898, new_AGEMA_signal_4902,
         new_AGEMA_signal_4906, new_AGEMA_signal_4910, new_AGEMA_signal_4914,
         new_AGEMA_signal_4918, new_AGEMA_signal_4922, new_AGEMA_signal_4926,
         new_AGEMA_signal_4930, new_AGEMA_signal_4934, new_AGEMA_signal_4938,
         new_AGEMA_signal_4942, new_AGEMA_signal_4946, new_AGEMA_signal_4950,
         new_AGEMA_signal_4954, new_AGEMA_signal_4958, new_AGEMA_signal_4962,
         new_AGEMA_signal_4966, new_AGEMA_signal_4970, new_AGEMA_signal_4974,
         new_AGEMA_signal_4978, new_AGEMA_signal_4982, new_AGEMA_signal_4986,
         new_AGEMA_signal_4990, new_AGEMA_signal_4994, new_AGEMA_signal_4998,
         new_AGEMA_signal_5002, new_AGEMA_signal_5006, new_AGEMA_signal_5010,
         new_AGEMA_signal_5014, new_AGEMA_signal_5018, new_AGEMA_signal_5022,
         new_AGEMA_signal_5026, new_AGEMA_signal_5030, new_AGEMA_signal_5034,
         new_AGEMA_signal_5038, new_AGEMA_signal_5042, new_AGEMA_signal_5046,
         new_AGEMA_signal_5050, new_AGEMA_signal_5054, new_AGEMA_signal_5058,
         new_AGEMA_signal_5062, new_AGEMA_signal_5066, new_AGEMA_signal_5070,
         new_AGEMA_signal_5074, new_AGEMA_signal_5078, new_AGEMA_signal_5082,
         new_AGEMA_signal_5086, new_AGEMA_signal_5090, new_AGEMA_signal_5094,
         new_AGEMA_signal_5098, new_AGEMA_signal_5102, new_AGEMA_signal_5106,
         new_AGEMA_signal_5110, new_AGEMA_signal_5114, new_AGEMA_signal_5118,
         new_AGEMA_signal_5122, new_AGEMA_signal_5126, new_AGEMA_signal_5130,
         new_AGEMA_signal_5134, new_AGEMA_signal_5138, new_AGEMA_signal_5142,
         new_AGEMA_signal_5146, new_AGEMA_signal_5150, new_AGEMA_signal_5154,
         new_AGEMA_signal_5158, new_AGEMA_signal_5162, new_AGEMA_signal_5166,
         new_AGEMA_signal_5170, new_AGEMA_signal_5174, new_AGEMA_signal_5178,
         new_AGEMA_signal_5182, new_AGEMA_signal_5186, new_AGEMA_signal_5190,
         new_AGEMA_signal_5194, new_AGEMA_signal_5198, new_AGEMA_signal_5202,
         new_AGEMA_signal_5206, new_AGEMA_signal_5210, new_AGEMA_signal_5214,
         new_AGEMA_signal_5218, new_AGEMA_signal_5222, new_AGEMA_signal_5226,
         new_AGEMA_signal_5230, new_AGEMA_signal_5234, new_AGEMA_signal_5238,
         new_AGEMA_signal_5242, new_AGEMA_signal_5246, new_AGEMA_signal_5250,
         new_AGEMA_signal_5254, new_AGEMA_signal_5258, new_AGEMA_signal_5262,
         new_AGEMA_signal_5266, new_AGEMA_signal_5270, new_AGEMA_signal_5274,
         new_AGEMA_signal_5278, new_AGEMA_signal_5282, new_AGEMA_signal_5286,
         new_AGEMA_signal_5290, new_AGEMA_signal_5294, new_AGEMA_signal_5298,
         new_AGEMA_signal_5302, new_AGEMA_signal_5306, new_AGEMA_signal_5310,
         new_AGEMA_signal_5314, new_AGEMA_signal_5318, new_AGEMA_signal_5322,
         new_AGEMA_signal_5326, new_AGEMA_signal_5330, new_AGEMA_signal_5334,
         new_AGEMA_signal_5338, new_AGEMA_signal_5342, new_AGEMA_signal_5346,
         new_AGEMA_signal_5350, new_AGEMA_signal_5354, new_AGEMA_signal_5358,
         new_AGEMA_signal_5362, new_AGEMA_signal_5366, new_AGEMA_signal_5370,
         new_AGEMA_signal_5374, new_AGEMA_signal_5378, new_AGEMA_signal_5382,
         new_AGEMA_signal_5386, new_AGEMA_signal_5390, new_AGEMA_signal_5394,
         new_AGEMA_signal_5398, new_AGEMA_signal_5402, new_AGEMA_signal_5406,
         new_AGEMA_signal_5410, new_AGEMA_signal_5414, new_AGEMA_signal_5418,
         new_AGEMA_signal_5422, new_AGEMA_signal_5426, new_AGEMA_signal_5430,
         new_AGEMA_signal_5434, new_AGEMA_signal_5438, new_AGEMA_signal_5442,
         new_AGEMA_signal_5446, new_AGEMA_signal_5450, new_AGEMA_signal_5454,
         new_AGEMA_signal_5458, new_AGEMA_signal_5462, new_AGEMA_signal_5466,
         new_AGEMA_signal_5470, new_AGEMA_signal_5474, new_AGEMA_signal_5478,
         new_AGEMA_signal_5482, new_AGEMA_signal_5486, new_AGEMA_signal_5490,
         new_AGEMA_signal_5494, new_AGEMA_signal_5498, new_AGEMA_signal_5502,
         new_AGEMA_signal_5506, new_AGEMA_signal_5510, new_AGEMA_signal_5514,
         new_AGEMA_signal_5518, new_AGEMA_signal_5522, new_AGEMA_signal_5526,
         new_AGEMA_signal_5530, new_AGEMA_signal_5534, new_AGEMA_signal_5538,
         new_AGEMA_signal_5542, new_AGEMA_signal_5546, new_AGEMA_signal_5550,
         new_AGEMA_signal_5554, new_AGEMA_signal_5558, new_AGEMA_signal_5562,
         new_AGEMA_signal_5566, new_AGEMA_signal_5570, new_AGEMA_signal_5574,
         new_AGEMA_signal_5578, new_AGEMA_signal_5582, new_AGEMA_signal_5586,
         new_AGEMA_signal_5590, new_AGEMA_signal_5594, new_AGEMA_signal_5598,
         new_AGEMA_signal_5602, new_AGEMA_signal_5606, new_AGEMA_signal_5610,
         new_AGEMA_signal_5614, new_AGEMA_signal_5618, new_AGEMA_signal_5622,
         new_AGEMA_signal_5626, new_AGEMA_signal_5630, new_AGEMA_signal_5634,
         new_AGEMA_signal_5638, new_AGEMA_signal_5642, new_AGEMA_signal_5646,
         new_AGEMA_signal_5650, new_AGEMA_signal_5654, new_AGEMA_signal_5658,
         new_AGEMA_signal_5662, new_AGEMA_signal_5666, new_AGEMA_signal_5670,
         new_AGEMA_signal_5674, new_AGEMA_signal_5678, new_AGEMA_signal_5682,
         new_AGEMA_signal_5686, new_AGEMA_signal_5690, new_AGEMA_signal_5694,
         new_AGEMA_signal_5698, new_AGEMA_signal_5702, new_AGEMA_signal_5706,
         new_AGEMA_signal_5710, new_AGEMA_signal_5714, new_AGEMA_signal_5718,
         new_AGEMA_signal_5722, new_AGEMA_signal_5726, new_AGEMA_signal_5730,
         new_AGEMA_signal_5734, new_AGEMA_signal_5738, new_AGEMA_signal_5742,
         new_AGEMA_signal_5746, new_AGEMA_signal_5750, new_AGEMA_signal_5754,
         new_AGEMA_signal_5758, new_AGEMA_signal_5762, new_AGEMA_signal_5766,
         new_AGEMA_signal_5770, new_AGEMA_signal_5774, new_AGEMA_signal_5778,
         new_AGEMA_signal_5782, new_AGEMA_signal_5786, new_AGEMA_signal_5790,
         new_AGEMA_signal_5794, new_AGEMA_signal_5798, new_AGEMA_signal_5802,
         new_AGEMA_signal_5806, new_AGEMA_signal_5810, new_AGEMA_signal_5814,
         new_AGEMA_signal_5818, new_AGEMA_signal_5822, new_AGEMA_signal_5826,
         new_AGEMA_signal_5830, new_AGEMA_signal_5834, new_AGEMA_signal_5838,
         new_AGEMA_signal_5842, new_AGEMA_signal_5846, new_AGEMA_signal_5850,
         new_AGEMA_signal_5854, new_AGEMA_signal_5858, new_AGEMA_signal_5862,
         new_AGEMA_signal_5866, new_AGEMA_signal_5870, new_AGEMA_signal_5874,
         new_AGEMA_signal_5878, new_AGEMA_signal_5882, new_AGEMA_signal_5886,
         new_AGEMA_signal_5890, new_AGEMA_signal_5894, new_AGEMA_signal_5898,
         new_AGEMA_signal_5902, new_AGEMA_signal_5906, new_AGEMA_signal_5910,
         new_AGEMA_signal_5914, new_AGEMA_signal_5918, new_AGEMA_signal_5922,
         new_AGEMA_signal_5926, new_AGEMA_signal_5930, new_AGEMA_signal_5934,
         new_AGEMA_signal_5938, new_AGEMA_signal_5942, new_AGEMA_signal_5946,
         new_AGEMA_signal_5950, new_AGEMA_signal_5954, new_AGEMA_signal_5958,
         new_AGEMA_signal_5962, new_AGEMA_signal_5966, new_AGEMA_signal_5970,
         new_AGEMA_signal_5974, new_AGEMA_signal_5978, new_AGEMA_signal_5982,
         new_AGEMA_signal_5986, new_AGEMA_signal_5990, new_AGEMA_signal_5994,
         new_AGEMA_signal_5998, new_AGEMA_signal_6002, new_AGEMA_signal_6006,
         new_AGEMA_signal_6010, new_AGEMA_signal_6014, new_AGEMA_signal_6018,
         new_AGEMA_signal_6022, new_AGEMA_signal_6026, new_AGEMA_signal_6030,
         new_AGEMA_signal_6034, new_AGEMA_signal_6038, new_AGEMA_signal_6042,
         new_AGEMA_signal_6046, new_AGEMA_signal_6050, new_AGEMA_signal_6054,
         new_AGEMA_signal_6058, new_AGEMA_signal_6062, new_AGEMA_signal_6066,
         new_AGEMA_signal_6070, new_AGEMA_signal_6074, new_AGEMA_signal_6078,
         new_AGEMA_signal_6082, new_AGEMA_signal_6086, new_AGEMA_signal_6090,
         new_AGEMA_signal_6094, new_AGEMA_signal_6098, new_AGEMA_signal_6102,
         new_AGEMA_signal_6106, new_AGEMA_signal_6110, new_AGEMA_signal_6114,
         new_AGEMA_signal_6118, new_AGEMA_signal_6122, new_AGEMA_signal_6126,
         new_AGEMA_signal_6130, new_AGEMA_signal_6134, new_AGEMA_signal_6138,
         new_AGEMA_signal_6142, new_AGEMA_signal_6146, new_AGEMA_signal_6150,
         new_AGEMA_signal_6154, new_AGEMA_signal_6158, new_AGEMA_signal_6162,
         new_AGEMA_signal_6166, new_AGEMA_signal_6170, new_AGEMA_signal_6174,
         new_AGEMA_signal_6178, new_AGEMA_signal_6182, new_AGEMA_signal_6186,
         new_AGEMA_signal_6190, new_AGEMA_signal_6194, new_AGEMA_signal_6198,
         new_AGEMA_signal_6202, new_AGEMA_signal_6206, new_AGEMA_signal_6210,
         new_AGEMA_signal_6214, new_AGEMA_signal_6218, new_AGEMA_signal_6222,
         new_AGEMA_signal_6226, new_AGEMA_signal_3384, Inst_bSbox_M25,
         new_AGEMA_signal_3388, Inst_bSbox_M26, new_AGEMA_signal_3611,
         new_AGEMA_signal_3610, new_AGEMA_signal_3389, Inst_bSbox_M28,
         new_AGEMA_signal_3613, new_AGEMA_signal_3612, new_AGEMA_signal_3390,
         Inst_bSbox_M31, new_AGEMA_signal_3391, Inst_bSbox_M33,
         new_AGEMA_signal_3615, new_AGEMA_signal_3614, new_AGEMA_signal_3386,
         Inst_bSbox_M34, new_AGEMA_signal_3396, Inst_bSbox_M36,
         new_AGEMA_signal_3617, new_AGEMA_signal_3616, new_AGEMA_signal_3627,
         new_AGEMA_signal_3631, new_AGEMA_signal_3635, new_AGEMA_signal_3639,
         new_AGEMA_signal_3643, new_AGEMA_signal_3647, new_AGEMA_signal_3651,
         new_AGEMA_signal_3655, new_AGEMA_signal_3659, new_AGEMA_signal_3663,
         new_AGEMA_signal_3667, new_AGEMA_signal_3671, new_AGEMA_signal_3675,
         new_AGEMA_signal_3679, new_AGEMA_signal_3683, new_AGEMA_signal_3687,
         new_AGEMA_signal_3691, new_AGEMA_signal_3695, new_AGEMA_signal_3699,
         new_AGEMA_signal_3703, new_AGEMA_signal_3707, new_AGEMA_signal_3711,
         new_AGEMA_signal_3715, new_AGEMA_signal_3719, new_AGEMA_signal_3723,
         new_AGEMA_signal_3727, new_AGEMA_signal_3731, new_AGEMA_signal_3735,
         new_AGEMA_signal_3739, new_AGEMA_signal_3743, new_AGEMA_signal_3747,
         new_AGEMA_signal_3751, new_AGEMA_signal_3755, new_AGEMA_signal_3759,
         new_AGEMA_signal_3763, new_AGEMA_signal_3767, new_AGEMA_signal_3771,
         new_AGEMA_signal_3775, new_AGEMA_signal_3779, new_AGEMA_signal_3783,
         new_AGEMA_signal_3787, new_AGEMA_signal_3791, new_AGEMA_signal_3795,
         new_AGEMA_signal_3799, new_AGEMA_signal_3803, new_AGEMA_signal_3807,
         new_AGEMA_signal_3811, new_AGEMA_signal_3815, new_AGEMA_signal_3819,
         new_AGEMA_signal_3823, new_AGEMA_signal_3827, new_AGEMA_signal_3831,
         new_AGEMA_signal_3835, new_AGEMA_signal_3839, new_AGEMA_signal_3843,
         new_AGEMA_signal_3847, new_AGEMA_signal_3851, new_AGEMA_signal_3855,
         new_AGEMA_signal_3859, new_AGEMA_signal_3863, new_AGEMA_signal_3867,
         new_AGEMA_signal_3871, new_AGEMA_signal_3875, new_AGEMA_signal_3879,
         new_AGEMA_signal_3883, new_AGEMA_signal_3887, new_AGEMA_signal_3891,
         new_AGEMA_signal_3895, new_AGEMA_signal_3899, new_AGEMA_signal_3903,
         new_AGEMA_signal_3907, new_AGEMA_signal_3911, new_AGEMA_signal_3915,
         new_AGEMA_signal_3919, new_AGEMA_signal_3923, new_AGEMA_signal_3927,
         new_AGEMA_signal_3931, new_AGEMA_signal_3935, new_AGEMA_signal_3939,
         new_AGEMA_signal_3943, new_AGEMA_signal_3947, new_AGEMA_signal_3951,
         new_AGEMA_signal_3955, new_AGEMA_signal_3959, new_AGEMA_signal_3963,
         new_AGEMA_signal_3967, new_AGEMA_signal_3971, new_AGEMA_signal_3975,
         new_AGEMA_signal_3979, new_AGEMA_signal_3983, new_AGEMA_signal_3987,
         new_AGEMA_signal_3991, new_AGEMA_signal_3995, new_AGEMA_signal_3999,
         new_AGEMA_signal_4003, new_AGEMA_signal_4007, new_AGEMA_signal_4011,
         new_AGEMA_signal_4015, new_AGEMA_signal_4019, new_AGEMA_signal_4023,
         new_AGEMA_signal_4027, new_AGEMA_signal_4031, new_AGEMA_signal_4035,
         new_AGEMA_signal_4039, new_AGEMA_signal_4043, new_AGEMA_signal_4047,
         new_AGEMA_signal_4051, new_AGEMA_signal_4055, new_AGEMA_signal_4059,
         new_AGEMA_signal_4063, new_AGEMA_signal_4067, new_AGEMA_signal_4071,
         new_AGEMA_signal_4075, new_AGEMA_signal_4079, new_AGEMA_signal_4083,
         new_AGEMA_signal_4087, new_AGEMA_signal_4091, new_AGEMA_signal_4095,
         new_AGEMA_signal_4099, new_AGEMA_signal_4103, new_AGEMA_signal_4107,
         new_AGEMA_signal_4111, new_AGEMA_signal_4115, new_AGEMA_signal_4119,
         new_AGEMA_signal_4123, new_AGEMA_signal_4127, new_AGEMA_signal_4131,
         new_AGEMA_signal_4134, new_AGEMA_signal_4137, new_AGEMA_signal_4140,
         new_AGEMA_signal_4143, new_AGEMA_signal_4146, new_AGEMA_signal_4149,
         new_AGEMA_signal_4152, new_AGEMA_signal_4155, new_AGEMA_signal_4158,
         new_AGEMA_signal_4161, new_AGEMA_signal_4164, new_AGEMA_signal_4167,
         new_AGEMA_signal_4170, new_AGEMA_signal_4173, new_AGEMA_signal_4176,
         new_AGEMA_signal_4179, new_AGEMA_signal_4182, new_AGEMA_signal_4185,
         new_AGEMA_signal_4188, new_AGEMA_signal_4191, new_AGEMA_signal_4194,
         new_AGEMA_signal_4197, new_AGEMA_signal_4200, new_AGEMA_signal_4203,
         new_AGEMA_signal_4206, new_AGEMA_signal_4209, new_AGEMA_signal_4212,
         new_AGEMA_signal_4215, new_AGEMA_signal_4218, new_AGEMA_signal_4221,
         new_AGEMA_signal_4224, new_AGEMA_signal_4227, new_AGEMA_signal_4230,
         new_AGEMA_signal_4233, new_AGEMA_signal_4236, new_AGEMA_signal_4239,
         new_AGEMA_signal_4243, new_AGEMA_signal_4247, new_AGEMA_signal_4251,
         new_AGEMA_signal_4255, new_AGEMA_signal_4259, new_AGEMA_signal_4263,
         new_AGEMA_signal_4267, new_AGEMA_signal_4271, new_AGEMA_signal_4275,
         new_AGEMA_signal_4279, new_AGEMA_signal_4283, new_AGEMA_signal_4287,
         new_AGEMA_signal_4291, new_AGEMA_signal_4295, new_AGEMA_signal_4299,
         new_AGEMA_signal_4303, new_AGEMA_signal_4307, new_AGEMA_signal_4311,
         new_AGEMA_signal_4315, new_AGEMA_signal_4319, new_AGEMA_signal_4323,
         new_AGEMA_signal_4327, new_AGEMA_signal_4331, new_AGEMA_signal_4335,
         new_AGEMA_signal_4339, new_AGEMA_signal_4343, new_AGEMA_signal_4347,
         new_AGEMA_signal_4351, new_AGEMA_signal_4355, new_AGEMA_signal_4359,
         new_AGEMA_signal_4363, new_AGEMA_signal_4367, new_AGEMA_signal_4371,
         new_AGEMA_signal_4375, new_AGEMA_signal_4379, new_AGEMA_signal_4383,
         new_AGEMA_signal_4387, new_AGEMA_signal_4391, new_AGEMA_signal_4395,
         new_AGEMA_signal_4399, new_AGEMA_signal_4403, new_AGEMA_signal_4407,
         new_AGEMA_signal_4411, new_AGEMA_signal_4415, new_AGEMA_signal_4419,
         new_AGEMA_signal_4423, new_AGEMA_signal_4427, new_AGEMA_signal_4431,
         new_AGEMA_signal_4435, new_AGEMA_signal_4439, new_AGEMA_signal_4443,
         new_AGEMA_signal_4447, new_AGEMA_signal_4451, new_AGEMA_signal_4455,
         new_AGEMA_signal_4459, new_AGEMA_signal_4463, new_AGEMA_signal_4467,
         new_AGEMA_signal_4471, new_AGEMA_signal_4475, new_AGEMA_signal_4479,
         new_AGEMA_signal_4483, new_AGEMA_signal_4487, new_AGEMA_signal_4491,
         new_AGEMA_signal_4495, new_AGEMA_signal_4499, new_AGEMA_signal_4503,
         new_AGEMA_signal_4507, new_AGEMA_signal_4511, new_AGEMA_signal_4515,
         new_AGEMA_signal_4519, new_AGEMA_signal_4523, new_AGEMA_signal_4527,
         new_AGEMA_signal_4531, new_AGEMA_signal_4535, new_AGEMA_signal_4539,
         new_AGEMA_signal_4543, new_AGEMA_signal_4547, new_AGEMA_signal_4551,
         new_AGEMA_signal_4555, new_AGEMA_signal_4559, new_AGEMA_signal_4563,
         new_AGEMA_signal_4567, new_AGEMA_signal_4571, new_AGEMA_signal_4575,
         new_AGEMA_signal_4579, new_AGEMA_signal_4583, new_AGEMA_signal_4587,
         new_AGEMA_signal_4591, new_AGEMA_signal_4595, new_AGEMA_signal_4599,
         new_AGEMA_signal_4603, new_AGEMA_signal_4607, new_AGEMA_signal_4611,
         new_AGEMA_signal_4615, new_AGEMA_signal_4619, new_AGEMA_signal_4623,
         new_AGEMA_signal_4627, new_AGEMA_signal_4631, new_AGEMA_signal_4635,
         new_AGEMA_signal_4639, new_AGEMA_signal_4643, new_AGEMA_signal_4647,
         new_AGEMA_signal_4651, new_AGEMA_signal_4655, new_AGEMA_signal_4659,
         new_AGEMA_signal_4663, new_AGEMA_signal_4667, new_AGEMA_signal_4671,
         new_AGEMA_signal_4675, new_AGEMA_signal_4679, new_AGEMA_signal_4683,
         new_AGEMA_signal_4687, new_AGEMA_signal_4691, new_AGEMA_signal_4695,
         new_AGEMA_signal_4699, new_AGEMA_signal_4703, new_AGEMA_signal_4707,
         new_AGEMA_signal_4711, new_AGEMA_signal_4715, new_AGEMA_signal_4719,
         new_AGEMA_signal_4723, new_AGEMA_signal_4727, new_AGEMA_signal_4731,
         new_AGEMA_signal_4735, new_AGEMA_signal_4739, new_AGEMA_signal_4743,
         new_AGEMA_signal_4747, new_AGEMA_signal_4751, new_AGEMA_signal_4755,
         new_AGEMA_signal_4759, new_AGEMA_signal_4763, new_AGEMA_signal_4767,
         new_AGEMA_signal_4771, new_AGEMA_signal_4775, new_AGEMA_signal_4779,
         new_AGEMA_signal_4783, new_AGEMA_signal_4787, new_AGEMA_signal_4791,
         new_AGEMA_signal_4795, new_AGEMA_signal_4799, new_AGEMA_signal_4803,
         new_AGEMA_signal_4807, new_AGEMA_signal_4811, new_AGEMA_signal_4815,
         new_AGEMA_signal_4819, new_AGEMA_signal_4823, new_AGEMA_signal_4827,
         new_AGEMA_signal_4831, new_AGEMA_signal_4835, new_AGEMA_signal_4839,
         new_AGEMA_signal_4843, new_AGEMA_signal_4847, new_AGEMA_signal_4851,
         new_AGEMA_signal_4855, new_AGEMA_signal_4859, new_AGEMA_signal_4863,
         new_AGEMA_signal_4867, new_AGEMA_signal_4871, new_AGEMA_signal_4875,
         new_AGEMA_signal_4879, new_AGEMA_signal_4883, new_AGEMA_signal_4887,
         new_AGEMA_signal_4891, new_AGEMA_signal_4895, new_AGEMA_signal_4899,
         new_AGEMA_signal_4903, new_AGEMA_signal_4907, new_AGEMA_signal_4911,
         new_AGEMA_signal_4915, new_AGEMA_signal_4919, new_AGEMA_signal_4923,
         new_AGEMA_signal_4927, new_AGEMA_signal_4931, new_AGEMA_signal_4935,
         new_AGEMA_signal_4939, new_AGEMA_signal_4943, new_AGEMA_signal_4947,
         new_AGEMA_signal_4951, new_AGEMA_signal_4955, new_AGEMA_signal_4959,
         new_AGEMA_signal_4963, new_AGEMA_signal_4967, new_AGEMA_signal_4971,
         new_AGEMA_signal_4975, new_AGEMA_signal_4979, new_AGEMA_signal_4983,
         new_AGEMA_signal_4987, new_AGEMA_signal_4991, new_AGEMA_signal_4995,
         new_AGEMA_signal_4999, new_AGEMA_signal_5003, new_AGEMA_signal_5007,
         new_AGEMA_signal_5011, new_AGEMA_signal_5015, new_AGEMA_signal_5019,
         new_AGEMA_signal_5023, new_AGEMA_signal_5027, new_AGEMA_signal_5031,
         new_AGEMA_signal_5035, new_AGEMA_signal_5039, new_AGEMA_signal_5043,
         new_AGEMA_signal_5047, new_AGEMA_signal_5051, new_AGEMA_signal_5055,
         new_AGEMA_signal_5059, new_AGEMA_signal_5063, new_AGEMA_signal_5067,
         new_AGEMA_signal_5071, new_AGEMA_signal_5075, new_AGEMA_signal_5079,
         new_AGEMA_signal_5083, new_AGEMA_signal_5087, new_AGEMA_signal_5091,
         new_AGEMA_signal_5095, new_AGEMA_signal_5099, new_AGEMA_signal_5103,
         new_AGEMA_signal_5107, new_AGEMA_signal_5111, new_AGEMA_signal_5115,
         new_AGEMA_signal_5119, new_AGEMA_signal_5123, new_AGEMA_signal_5127,
         new_AGEMA_signal_5131, new_AGEMA_signal_5135, new_AGEMA_signal_5139,
         new_AGEMA_signal_5143, new_AGEMA_signal_5147, new_AGEMA_signal_5151,
         new_AGEMA_signal_5155, new_AGEMA_signal_5159, new_AGEMA_signal_5163,
         new_AGEMA_signal_5167, new_AGEMA_signal_5171, new_AGEMA_signal_5175,
         new_AGEMA_signal_5179, new_AGEMA_signal_5183, new_AGEMA_signal_5187,
         new_AGEMA_signal_5191, new_AGEMA_signal_5195, new_AGEMA_signal_5199,
         new_AGEMA_signal_5203, new_AGEMA_signal_5207, new_AGEMA_signal_5211,
         new_AGEMA_signal_5215, new_AGEMA_signal_5219, new_AGEMA_signal_5223,
         new_AGEMA_signal_5227, new_AGEMA_signal_5231, new_AGEMA_signal_5235,
         new_AGEMA_signal_5239, new_AGEMA_signal_5243, new_AGEMA_signal_5247,
         new_AGEMA_signal_5251, new_AGEMA_signal_5255, new_AGEMA_signal_5259,
         new_AGEMA_signal_5263, new_AGEMA_signal_5267, new_AGEMA_signal_5271,
         new_AGEMA_signal_5275, new_AGEMA_signal_5279, new_AGEMA_signal_5283,
         new_AGEMA_signal_5287, new_AGEMA_signal_5291, new_AGEMA_signal_5295,
         new_AGEMA_signal_5299, new_AGEMA_signal_5303, new_AGEMA_signal_5307,
         new_AGEMA_signal_5311, new_AGEMA_signal_5315, new_AGEMA_signal_5319,
         new_AGEMA_signal_5323, new_AGEMA_signal_5327, new_AGEMA_signal_5331,
         new_AGEMA_signal_5335, new_AGEMA_signal_5339, new_AGEMA_signal_5343,
         new_AGEMA_signal_5347, new_AGEMA_signal_5351, new_AGEMA_signal_5355,
         new_AGEMA_signal_5359, new_AGEMA_signal_5363, new_AGEMA_signal_5367,
         new_AGEMA_signal_5371, new_AGEMA_signal_5375, new_AGEMA_signal_5379,
         new_AGEMA_signal_5383, new_AGEMA_signal_5387, new_AGEMA_signal_5391,
         new_AGEMA_signal_5395, new_AGEMA_signal_5399, new_AGEMA_signal_5403,
         new_AGEMA_signal_5407, new_AGEMA_signal_5411, new_AGEMA_signal_5415,
         new_AGEMA_signal_5419, new_AGEMA_signal_5423, new_AGEMA_signal_5427,
         new_AGEMA_signal_5431, new_AGEMA_signal_5435, new_AGEMA_signal_5439,
         new_AGEMA_signal_5443, new_AGEMA_signal_5447, new_AGEMA_signal_5451,
         new_AGEMA_signal_5455, new_AGEMA_signal_5459, new_AGEMA_signal_5463,
         new_AGEMA_signal_5467, new_AGEMA_signal_5471, new_AGEMA_signal_5475,
         new_AGEMA_signal_5479, new_AGEMA_signal_5483, new_AGEMA_signal_5487,
         new_AGEMA_signal_5491, new_AGEMA_signal_5495, new_AGEMA_signal_5499,
         new_AGEMA_signal_5503, new_AGEMA_signal_5507, new_AGEMA_signal_5511,
         new_AGEMA_signal_5515, new_AGEMA_signal_5519, new_AGEMA_signal_5523,
         new_AGEMA_signal_5527, new_AGEMA_signal_5531, new_AGEMA_signal_5535,
         new_AGEMA_signal_5539, new_AGEMA_signal_5543, new_AGEMA_signal_5547,
         new_AGEMA_signal_5551, new_AGEMA_signal_5555, new_AGEMA_signal_5559,
         new_AGEMA_signal_5563, new_AGEMA_signal_5567, new_AGEMA_signal_5571,
         new_AGEMA_signal_5575, new_AGEMA_signal_5579, new_AGEMA_signal_5583,
         new_AGEMA_signal_5587, new_AGEMA_signal_5591, new_AGEMA_signal_5595,
         new_AGEMA_signal_5599, new_AGEMA_signal_5603, new_AGEMA_signal_5607,
         new_AGEMA_signal_5611, new_AGEMA_signal_5615, new_AGEMA_signal_5619,
         new_AGEMA_signal_5623, new_AGEMA_signal_5627, new_AGEMA_signal_5631,
         new_AGEMA_signal_5635, new_AGEMA_signal_5639, new_AGEMA_signal_5643,
         new_AGEMA_signal_5647, new_AGEMA_signal_5651, new_AGEMA_signal_5655,
         new_AGEMA_signal_5659, new_AGEMA_signal_5663, new_AGEMA_signal_5667,
         new_AGEMA_signal_5671, new_AGEMA_signal_5675, new_AGEMA_signal_5679,
         new_AGEMA_signal_5683, new_AGEMA_signal_5687, new_AGEMA_signal_5691,
         new_AGEMA_signal_5695, new_AGEMA_signal_5699, new_AGEMA_signal_5703,
         new_AGEMA_signal_5707, new_AGEMA_signal_5711, new_AGEMA_signal_5715,
         new_AGEMA_signal_5719, new_AGEMA_signal_5723, new_AGEMA_signal_5727,
         new_AGEMA_signal_5731, new_AGEMA_signal_5735, new_AGEMA_signal_5739,
         new_AGEMA_signal_5743, new_AGEMA_signal_5747, new_AGEMA_signal_5751,
         new_AGEMA_signal_5755, new_AGEMA_signal_5759, new_AGEMA_signal_5763,
         new_AGEMA_signal_5767, new_AGEMA_signal_5771, new_AGEMA_signal_5775,
         new_AGEMA_signal_5779, new_AGEMA_signal_5783, new_AGEMA_signal_5787,
         new_AGEMA_signal_5791, new_AGEMA_signal_5795, new_AGEMA_signal_5799,
         new_AGEMA_signal_5803, new_AGEMA_signal_5807, new_AGEMA_signal_5811,
         new_AGEMA_signal_5815, new_AGEMA_signal_5819, new_AGEMA_signal_5823,
         new_AGEMA_signal_5827, new_AGEMA_signal_5831, new_AGEMA_signal_5835,
         new_AGEMA_signal_5839, new_AGEMA_signal_5843, new_AGEMA_signal_5847,
         new_AGEMA_signal_5851, new_AGEMA_signal_5855, new_AGEMA_signal_5859,
         new_AGEMA_signal_5863, new_AGEMA_signal_5867, new_AGEMA_signal_5871,
         new_AGEMA_signal_5875, new_AGEMA_signal_5879, new_AGEMA_signal_5883,
         new_AGEMA_signal_5887, new_AGEMA_signal_5891, new_AGEMA_signal_5895,
         new_AGEMA_signal_5899, new_AGEMA_signal_5903, new_AGEMA_signal_5907,
         new_AGEMA_signal_5911, new_AGEMA_signal_5915, new_AGEMA_signal_5919,
         new_AGEMA_signal_5923, new_AGEMA_signal_5927, new_AGEMA_signal_5931,
         new_AGEMA_signal_5935, new_AGEMA_signal_5939, new_AGEMA_signal_5943,
         new_AGEMA_signal_5947, new_AGEMA_signal_5951, new_AGEMA_signal_5955,
         new_AGEMA_signal_5959, new_AGEMA_signal_5963, new_AGEMA_signal_5967,
         new_AGEMA_signal_5971, new_AGEMA_signal_5975, new_AGEMA_signal_5979,
         new_AGEMA_signal_5983, new_AGEMA_signal_5987, new_AGEMA_signal_5991,
         new_AGEMA_signal_5995, new_AGEMA_signal_5999, new_AGEMA_signal_6003,
         new_AGEMA_signal_6007, new_AGEMA_signal_6011, new_AGEMA_signal_6015,
         new_AGEMA_signal_6019, new_AGEMA_signal_6023, new_AGEMA_signal_6027,
         new_AGEMA_signal_6031, new_AGEMA_signal_6035, new_AGEMA_signal_6039,
         new_AGEMA_signal_6043, new_AGEMA_signal_6047, new_AGEMA_signal_6051,
         new_AGEMA_signal_6055, new_AGEMA_signal_6059, new_AGEMA_signal_6063,
         new_AGEMA_signal_6067, new_AGEMA_signal_6071, new_AGEMA_signal_6075,
         new_AGEMA_signal_6079, new_AGEMA_signal_6083, new_AGEMA_signal_6087,
         new_AGEMA_signal_6091, new_AGEMA_signal_6095, new_AGEMA_signal_6099,
         new_AGEMA_signal_6103, new_AGEMA_signal_6107, new_AGEMA_signal_6111,
         new_AGEMA_signal_6115, new_AGEMA_signal_6119, new_AGEMA_signal_6123,
         new_AGEMA_signal_6127, new_AGEMA_signal_6131, new_AGEMA_signal_6135,
         new_AGEMA_signal_6139, new_AGEMA_signal_6143, new_AGEMA_signal_6147,
         new_AGEMA_signal_6151, new_AGEMA_signal_6155, new_AGEMA_signal_6159,
         new_AGEMA_signal_6163, new_AGEMA_signal_6167, new_AGEMA_signal_6171,
         new_AGEMA_signal_6175, new_AGEMA_signal_6179, new_AGEMA_signal_6183,
         new_AGEMA_signal_6187, new_AGEMA_signal_6191, new_AGEMA_signal_6195,
         new_AGEMA_signal_6199, new_AGEMA_signal_6203, new_AGEMA_signal_6207,
         new_AGEMA_signal_6211, new_AGEMA_signal_6215, new_AGEMA_signal_6219,
         new_AGEMA_signal_6223, new_AGEMA_signal_6227, new_AGEMA_signal_3392,
         Inst_bSbox_M29, new_AGEMA_signal_3393, Inst_bSbox_M30,
         new_AGEMA_signal_3394, Inst_bSbox_M32, new_AGEMA_signal_3395,
         Inst_bSbox_M35, new_AGEMA_signal_3397, Inst_bSbox_M37,
         new_AGEMA_signal_3619, new_AGEMA_signal_3618, new_AGEMA_signal_3398,
         Inst_bSbox_M38, new_AGEMA_signal_3621, new_AGEMA_signal_3620,
         new_AGEMA_signal_3399, Inst_bSbox_M39, new_AGEMA_signal_3623,
         new_AGEMA_signal_3622, new_AGEMA_signal_3400, Inst_bSbox_M40,
         new_AGEMA_signal_3625, new_AGEMA_signal_3624, new_AGEMA_signal_3401,
         Inst_bSbox_M41, new_AGEMA_signal_3402, Inst_bSbox_M42,
         new_AGEMA_signal_3403, Inst_bSbox_M43, new_AGEMA_signal_3404,
         Inst_bSbox_M44, new_AGEMA_signal_3413, Inst_bSbox_M45,
         new_AGEMA_signal_3628, new_AGEMA_signal_3632, new_AGEMA_signal_3636,
         new_AGEMA_signal_3640, new_AGEMA_signal_3644, new_AGEMA_signal_3648,
         new_AGEMA_signal_3652, new_AGEMA_signal_3656, new_AGEMA_signal_3660,
         new_AGEMA_signal_3664, new_AGEMA_signal_3668, new_AGEMA_signal_3672,
         new_AGEMA_signal_3676, new_AGEMA_signal_3680, new_AGEMA_signal_3684,
         new_AGEMA_signal_3688, new_AGEMA_signal_3692, new_AGEMA_signal_3696,
         new_AGEMA_signal_3700, new_AGEMA_signal_3704, new_AGEMA_signal_3708,
         new_AGEMA_signal_3712, new_AGEMA_signal_3716, new_AGEMA_signal_3720,
         new_AGEMA_signal_3724, new_AGEMA_signal_3728, new_AGEMA_signal_3732,
         new_AGEMA_signal_3736, new_AGEMA_signal_3740, new_AGEMA_signal_3744,
         new_AGEMA_signal_3748, new_AGEMA_signal_3752, new_AGEMA_signal_3756,
         new_AGEMA_signal_3760, new_AGEMA_signal_3764, new_AGEMA_signal_3768,
         new_AGEMA_signal_3772, new_AGEMA_signal_3776, new_AGEMA_signal_3780,
         new_AGEMA_signal_3784, new_AGEMA_signal_3788, new_AGEMA_signal_3792,
         new_AGEMA_signal_3796, new_AGEMA_signal_3800, new_AGEMA_signal_3804,
         new_AGEMA_signal_3808, new_AGEMA_signal_3812, new_AGEMA_signal_3816,
         new_AGEMA_signal_3820, new_AGEMA_signal_3824, new_AGEMA_signal_3828,
         new_AGEMA_signal_3832, new_AGEMA_signal_3836, new_AGEMA_signal_3840,
         new_AGEMA_signal_3844, new_AGEMA_signal_3848, new_AGEMA_signal_3852,
         new_AGEMA_signal_3856, new_AGEMA_signal_3860, new_AGEMA_signal_3864,
         new_AGEMA_signal_3868, new_AGEMA_signal_3872, new_AGEMA_signal_3876,
         new_AGEMA_signal_3880, new_AGEMA_signal_3884, new_AGEMA_signal_3888,
         new_AGEMA_signal_3892, new_AGEMA_signal_3896, new_AGEMA_signal_3900,
         new_AGEMA_signal_3904, new_AGEMA_signal_3908, new_AGEMA_signal_3912,
         new_AGEMA_signal_3916, new_AGEMA_signal_3920, new_AGEMA_signal_3924,
         new_AGEMA_signal_3928, new_AGEMA_signal_3932, new_AGEMA_signal_3936,
         new_AGEMA_signal_3940, new_AGEMA_signal_3944, new_AGEMA_signal_3948,
         new_AGEMA_signal_3952, new_AGEMA_signal_3956, new_AGEMA_signal_3960,
         new_AGEMA_signal_3964, new_AGEMA_signal_3968, new_AGEMA_signal_3972,
         new_AGEMA_signal_3976, new_AGEMA_signal_3980, new_AGEMA_signal_3984,
         new_AGEMA_signal_3988, new_AGEMA_signal_3992, new_AGEMA_signal_3996,
         new_AGEMA_signal_4000, new_AGEMA_signal_4004, new_AGEMA_signal_4008,
         new_AGEMA_signal_4012, new_AGEMA_signal_4016, new_AGEMA_signal_4020,
         new_AGEMA_signal_4024, new_AGEMA_signal_4028, new_AGEMA_signal_4032,
         new_AGEMA_signal_4036, new_AGEMA_signal_4040, new_AGEMA_signal_4044,
         new_AGEMA_signal_4048, new_AGEMA_signal_4052, new_AGEMA_signal_4056,
         new_AGEMA_signal_4060, new_AGEMA_signal_4064, new_AGEMA_signal_4068,
         new_AGEMA_signal_4072, new_AGEMA_signal_4076, new_AGEMA_signal_4080,
         new_AGEMA_signal_4084, new_AGEMA_signal_4088, new_AGEMA_signal_4092,
         new_AGEMA_signal_4096, new_AGEMA_signal_4100, new_AGEMA_signal_4104,
         new_AGEMA_signal_4108, new_AGEMA_signal_4112, new_AGEMA_signal_4116,
         new_AGEMA_signal_4120, new_AGEMA_signal_4124, new_AGEMA_signal_4128,
         new_AGEMA_signal_4132, new_AGEMA_signal_4135, new_AGEMA_signal_4138,
         new_AGEMA_signal_4141, new_AGEMA_signal_4144, new_AGEMA_signal_4147,
         new_AGEMA_signal_4150, new_AGEMA_signal_4153, new_AGEMA_signal_4156,
         new_AGEMA_signal_4159, new_AGEMA_signal_4162, new_AGEMA_signal_4165,
         new_AGEMA_signal_4168, new_AGEMA_signal_4171, new_AGEMA_signal_4174,
         new_AGEMA_signal_4177, new_AGEMA_signal_4180, new_AGEMA_signal_4183,
         new_AGEMA_signal_4186, new_AGEMA_signal_4189, new_AGEMA_signal_4192,
         new_AGEMA_signal_4195, new_AGEMA_signal_4198, new_AGEMA_signal_4201,
         new_AGEMA_signal_4204, new_AGEMA_signal_4207, new_AGEMA_signal_4210,
         new_AGEMA_signal_4213, new_AGEMA_signal_4216, new_AGEMA_signal_4219,
         new_AGEMA_signal_4222, new_AGEMA_signal_4225, new_AGEMA_signal_4228,
         new_AGEMA_signal_4231, new_AGEMA_signal_4234, new_AGEMA_signal_4237,
         new_AGEMA_signal_4240, new_AGEMA_signal_4244, new_AGEMA_signal_4248,
         new_AGEMA_signal_4252, new_AGEMA_signal_4256, new_AGEMA_signal_4260,
         new_AGEMA_signal_4264, new_AGEMA_signal_4268, new_AGEMA_signal_4272,
         new_AGEMA_signal_4276, new_AGEMA_signal_4280, new_AGEMA_signal_4284,
         new_AGEMA_signal_4288, new_AGEMA_signal_4292, new_AGEMA_signal_4296,
         new_AGEMA_signal_4300, new_AGEMA_signal_4304, new_AGEMA_signal_4308,
         new_AGEMA_signal_4312, new_AGEMA_signal_4316, new_AGEMA_signal_4320,
         new_AGEMA_signal_4324, new_AGEMA_signal_4328, new_AGEMA_signal_4332,
         new_AGEMA_signal_4336, new_AGEMA_signal_4340, new_AGEMA_signal_4344,
         new_AGEMA_signal_4348, new_AGEMA_signal_4352, new_AGEMA_signal_4356,
         new_AGEMA_signal_4360, new_AGEMA_signal_4364, new_AGEMA_signal_4368,
         new_AGEMA_signal_4372, new_AGEMA_signal_4376, new_AGEMA_signal_4380,
         new_AGEMA_signal_4384, new_AGEMA_signal_4388, new_AGEMA_signal_4392,
         new_AGEMA_signal_4396, new_AGEMA_signal_4400, new_AGEMA_signal_4404,
         new_AGEMA_signal_4408, new_AGEMA_signal_4412, new_AGEMA_signal_4416,
         new_AGEMA_signal_4420, new_AGEMA_signal_4424, new_AGEMA_signal_4428,
         new_AGEMA_signal_4432, new_AGEMA_signal_4436, new_AGEMA_signal_4440,
         new_AGEMA_signal_4444, new_AGEMA_signal_4448, new_AGEMA_signal_4452,
         new_AGEMA_signal_4456, new_AGEMA_signal_4460, new_AGEMA_signal_4464,
         new_AGEMA_signal_4468, new_AGEMA_signal_4472, new_AGEMA_signal_4476,
         new_AGEMA_signal_4480, new_AGEMA_signal_4484, new_AGEMA_signal_4488,
         new_AGEMA_signal_4492, new_AGEMA_signal_4496, new_AGEMA_signal_4500,
         new_AGEMA_signal_4504, new_AGEMA_signal_4508, new_AGEMA_signal_4512,
         new_AGEMA_signal_4516, new_AGEMA_signal_4520, new_AGEMA_signal_4524,
         new_AGEMA_signal_4528, new_AGEMA_signal_4532, new_AGEMA_signal_4536,
         new_AGEMA_signal_4540, new_AGEMA_signal_4544, new_AGEMA_signal_4548,
         new_AGEMA_signal_4552, new_AGEMA_signal_4556, new_AGEMA_signal_4560,
         new_AGEMA_signal_4564, new_AGEMA_signal_4568, new_AGEMA_signal_4572,
         new_AGEMA_signal_4576, new_AGEMA_signal_4580, new_AGEMA_signal_4584,
         new_AGEMA_signal_4588, new_AGEMA_signal_4592, new_AGEMA_signal_4596,
         new_AGEMA_signal_4600, new_AGEMA_signal_4604, new_AGEMA_signal_4608,
         new_AGEMA_signal_4612, new_AGEMA_signal_4616, new_AGEMA_signal_4620,
         new_AGEMA_signal_4624, new_AGEMA_signal_4628, new_AGEMA_signal_4632,
         new_AGEMA_signal_4636, new_AGEMA_signal_4640, new_AGEMA_signal_4644,
         new_AGEMA_signal_4648, new_AGEMA_signal_4652, new_AGEMA_signal_4656,
         new_AGEMA_signal_4660, new_AGEMA_signal_4664, new_AGEMA_signal_4668,
         new_AGEMA_signal_4672, new_AGEMA_signal_4676, new_AGEMA_signal_4680,
         new_AGEMA_signal_4684, new_AGEMA_signal_4688, new_AGEMA_signal_4692,
         new_AGEMA_signal_4696, new_AGEMA_signal_4700, new_AGEMA_signal_4704,
         new_AGEMA_signal_4708, new_AGEMA_signal_4712, new_AGEMA_signal_4716,
         new_AGEMA_signal_4720, new_AGEMA_signal_4724, new_AGEMA_signal_4728,
         new_AGEMA_signal_4732, new_AGEMA_signal_4736, new_AGEMA_signal_4740,
         new_AGEMA_signal_4744, new_AGEMA_signal_4748, new_AGEMA_signal_4752,
         new_AGEMA_signal_4756, new_AGEMA_signal_4760, new_AGEMA_signal_4764,
         new_AGEMA_signal_4768, new_AGEMA_signal_4772, new_AGEMA_signal_4776,
         new_AGEMA_signal_4780, new_AGEMA_signal_4784, new_AGEMA_signal_4788,
         new_AGEMA_signal_4792, new_AGEMA_signal_4796, new_AGEMA_signal_4800,
         new_AGEMA_signal_4804, new_AGEMA_signal_4808, new_AGEMA_signal_4812,
         new_AGEMA_signal_4816, new_AGEMA_signal_4820, new_AGEMA_signal_4824,
         new_AGEMA_signal_4828, new_AGEMA_signal_4832, new_AGEMA_signal_4836,
         new_AGEMA_signal_4840, new_AGEMA_signal_4844, new_AGEMA_signal_4848,
         new_AGEMA_signal_4852, new_AGEMA_signal_4856, new_AGEMA_signal_4860,
         new_AGEMA_signal_4864, new_AGEMA_signal_4868, new_AGEMA_signal_4872,
         new_AGEMA_signal_4876, new_AGEMA_signal_4880, new_AGEMA_signal_4884,
         new_AGEMA_signal_4888, new_AGEMA_signal_4892, new_AGEMA_signal_4896,
         new_AGEMA_signal_4900, new_AGEMA_signal_4904, new_AGEMA_signal_4908,
         new_AGEMA_signal_4912, new_AGEMA_signal_4916, new_AGEMA_signal_4920,
         new_AGEMA_signal_4924, new_AGEMA_signal_4928, new_AGEMA_signal_4932,
         new_AGEMA_signal_4936, new_AGEMA_signal_4940, new_AGEMA_signal_4944,
         new_AGEMA_signal_4948, new_AGEMA_signal_4952, new_AGEMA_signal_4956,
         new_AGEMA_signal_4960, new_AGEMA_signal_4964, new_AGEMA_signal_4968,
         new_AGEMA_signal_4972, new_AGEMA_signal_4976, new_AGEMA_signal_4980,
         new_AGEMA_signal_4984, new_AGEMA_signal_4988, new_AGEMA_signal_4992,
         new_AGEMA_signal_4996, new_AGEMA_signal_5000, new_AGEMA_signal_5004,
         new_AGEMA_signal_5008, new_AGEMA_signal_5012, new_AGEMA_signal_5016,
         new_AGEMA_signal_5020, new_AGEMA_signal_5024, new_AGEMA_signal_5028,
         new_AGEMA_signal_5032, new_AGEMA_signal_5036, new_AGEMA_signal_5040,
         new_AGEMA_signal_5044, new_AGEMA_signal_5048, new_AGEMA_signal_5052,
         new_AGEMA_signal_5056, new_AGEMA_signal_5060, new_AGEMA_signal_5064,
         new_AGEMA_signal_5068, new_AGEMA_signal_5072, new_AGEMA_signal_5076,
         new_AGEMA_signal_5080, new_AGEMA_signal_5084, new_AGEMA_signal_5088,
         new_AGEMA_signal_5092, new_AGEMA_signal_5096, new_AGEMA_signal_5100,
         new_AGEMA_signal_5104, new_AGEMA_signal_5108, new_AGEMA_signal_5112,
         new_AGEMA_signal_5116, new_AGEMA_signal_5120, new_AGEMA_signal_5124,
         new_AGEMA_signal_5128, new_AGEMA_signal_5132, new_AGEMA_signal_5136,
         new_AGEMA_signal_5140, new_AGEMA_signal_5144, new_AGEMA_signal_5148,
         new_AGEMA_signal_5152, new_AGEMA_signal_5156, new_AGEMA_signal_5160,
         new_AGEMA_signal_5164, new_AGEMA_signal_5168, new_AGEMA_signal_5172,
         new_AGEMA_signal_5176, new_AGEMA_signal_5180, new_AGEMA_signal_5184,
         new_AGEMA_signal_5188, new_AGEMA_signal_5192, new_AGEMA_signal_5196,
         new_AGEMA_signal_5200, new_AGEMA_signal_5204, new_AGEMA_signal_5208,
         new_AGEMA_signal_5212, new_AGEMA_signal_5216, new_AGEMA_signal_5220,
         new_AGEMA_signal_5224, new_AGEMA_signal_5228, new_AGEMA_signal_5232,
         new_AGEMA_signal_5236, new_AGEMA_signal_5240, new_AGEMA_signal_5244,
         new_AGEMA_signal_5248, new_AGEMA_signal_5252, new_AGEMA_signal_5256,
         new_AGEMA_signal_5260, new_AGEMA_signal_5264, new_AGEMA_signal_5268,
         new_AGEMA_signal_5272, new_AGEMA_signal_5276, new_AGEMA_signal_5280,
         new_AGEMA_signal_5284, new_AGEMA_signal_5288, new_AGEMA_signal_5292,
         new_AGEMA_signal_5296, new_AGEMA_signal_5300, new_AGEMA_signal_5304,
         new_AGEMA_signal_5308, new_AGEMA_signal_5312, new_AGEMA_signal_5316,
         new_AGEMA_signal_5320, new_AGEMA_signal_5324, new_AGEMA_signal_5328,
         new_AGEMA_signal_5332, new_AGEMA_signal_5336, new_AGEMA_signal_5340,
         new_AGEMA_signal_5344, new_AGEMA_signal_5348, new_AGEMA_signal_5352,
         new_AGEMA_signal_5356, new_AGEMA_signal_5360, new_AGEMA_signal_5364,
         new_AGEMA_signal_5368, new_AGEMA_signal_5372, new_AGEMA_signal_5376,
         new_AGEMA_signal_5380, new_AGEMA_signal_5384, new_AGEMA_signal_5388,
         new_AGEMA_signal_5392, new_AGEMA_signal_5396, new_AGEMA_signal_5400,
         new_AGEMA_signal_5404, new_AGEMA_signal_5408, new_AGEMA_signal_5412,
         new_AGEMA_signal_5416, new_AGEMA_signal_5420, new_AGEMA_signal_5424,
         new_AGEMA_signal_5428, new_AGEMA_signal_5432, new_AGEMA_signal_5436,
         new_AGEMA_signal_5440, new_AGEMA_signal_5444, new_AGEMA_signal_5448,
         new_AGEMA_signal_5452, new_AGEMA_signal_5456, new_AGEMA_signal_5460,
         new_AGEMA_signal_5464, new_AGEMA_signal_5468, new_AGEMA_signal_5472,
         new_AGEMA_signal_5476, new_AGEMA_signal_5480, new_AGEMA_signal_5484,
         new_AGEMA_signal_5488, new_AGEMA_signal_5492, new_AGEMA_signal_5496,
         new_AGEMA_signal_5500, new_AGEMA_signal_5504, new_AGEMA_signal_5508,
         new_AGEMA_signal_5512, new_AGEMA_signal_5516, new_AGEMA_signal_5520,
         new_AGEMA_signal_5524, new_AGEMA_signal_5528, new_AGEMA_signal_5532,
         new_AGEMA_signal_5536, new_AGEMA_signal_5540, new_AGEMA_signal_5544,
         new_AGEMA_signal_5548, new_AGEMA_signal_5552, new_AGEMA_signal_5556,
         new_AGEMA_signal_5560, new_AGEMA_signal_5564, new_AGEMA_signal_5568,
         new_AGEMA_signal_5572, new_AGEMA_signal_5576, new_AGEMA_signal_5580,
         new_AGEMA_signal_5584, new_AGEMA_signal_5588, new_AGEMA_signal_5592,
         new_AGEMA_signal_5596, new_AGEMA_signal_5600, new_AGEMA_signal_5604,
         new_AGEMA_signal_5608, new_AGEMA_signal_5612, new_AGEMA_signal_5616,
         new_AGEMA_signal_5620, new_AGEMA_signal_5624, new_AGEMA_signal_5628,
         new_AGEMA_signal_5632, new_AGEMA_signal_5636, new_AGEMA_signal_5640,
         new_AGEMA_signal_5644, new_AGEMA_signal_5648, new_AGEMA_signal_5652,
         new_AGEMA_signal_5656, new_AGEMA_signal_5660, new_AGEMA_signal_5664,
         new_AGEMA_signal_5668, new_AGEMA_signal_5672, new_AGEMA_signal_5676,
         new_AGEMA_signal_5680, new_AGEMA_signal_5684, new_AGEMA_signal_5688,
         new_AGEMA_signal_5692, new_AGEMA_signal_5696, new_AGEMA_signal_5700,
         new_AGEMA_signal_5704, new_AGEMA_signal_5708, new_AGEMA_signal_5712,
         new_AGEMA_signal_5716, new_AGEMA_signal_5720, new_AGEMA_signal_5724,
         new_AGEMA_signal_5728, new_AGEMA_signal_5732, new_AGEMA_signal_5736,
         new_AGEMA_signal_5740, new_AGEMA_signal_5744, new_AGEMA_signal_5748,
         new_AGEMA_signal_5752, new_AGEMA_signal_5756, new_AGEMA_signal_5760,
         new_AGEMA_signal_5764, new_AGEMA_signal_5768, new_AGEMA_signal_5772,
         new_AGEMA_signal_5776, new_AGEMA_signal_5780, new_AGEMA_signal_5784,
         new_AGEMA_signal_5788, new_AGEMA_signal_5792, new_AGEMA_signal_5796,
         new_AGEMA_signal_5800, new_AGEMA_signal_5804, new_AGEMA_signal_5808,
         new_AGEMA_signal_5812, new_AGEMA_signal_5816, new_AGEMA_signal_5820,
         new_AGEMA_signal_5824, new_AGEMA_signal_5828, new_AGEMA_signal_5832,
         new_AGEMA_signal_5836, new_AGEMA_signal_5840, new_AGEMA_signal_5844,
         new_AGEMA_signal_5848, new_AGEMA_signal_5852, new_AGEMA_signal_5856,
         new_AGEMA_signal_5860, new_AGEMA_signal_5864, new_AGEMA_signal_5868,
         new_AGEMA_signal_5872, new_AGEMA_signal_5876, new_AGEMA_signal_5880,
         new_AGEMA_signal_5884, new_AGEMA_signal_5888, new_AGEMA_signal_5892,
         new_AGEMA_signal_5896, new_AGEMA_signal_5900, new_AGEMA_signal_5904,
         new_AGEMA_signal_5908, new_AGEMA_signal_5912, new_AGEMA_signal_5916,
         new_AGEMA_signal_5920, new_AGEMA_signal_5924, new_AGEMA_signal_5928,
         new_AGEMA_signal_5932, new_AGEMA_signal_5936, new_AGEMA_signal_5940,
         new_AGEMA_signal_5944, new_AGEMA_signal_5948, new_AGEMA_signal_5952,
         new_AGEMA_signal_5956, new_AGEMA_signal_5960, new_AGEMA_signal_5964,
         new_AGEMA_signal_5968, new_AGEMA_signal_5972, new_AGEMA_signal_5976,
         new_AGEMA_signal_5980, new_AGEMA_signal_5984, new_AGEMA_signal_5988,
         new_AGEMA_signal_5992, new_AGEMA_signal_5996, new_AGEMA_signal_6000,
         new_AGEMA_signal_6004, new_AGEMA_signal_6008, new_AGEMA_signal_6012,
         new_AGEMA_signal_6016, new_AGEMA_signal_6020, new_AGEMA_signal_6024,
         new_AGEMA_signal_6028, new_AGEMA_signal_6032, new_AGEMA_signal_6036,
         new_AGEMA_signal_6040, new_AGEMA_signal_6044, new_AGEMA_signal_6048,
         new_AGEMA_signal_6052, new_AGEMA_signal_6056, new_AGEMA_signal_6060,
         new_AGEMA_signal_6064, new_AGEMA_signal_6068, new_AGEMA_signal_6072,
         new_AGEMA_signal_6076, new_AGEMA_signal_6080, new_AGEMA_signal_6084,
         new_AGEMA_signal_6088, new_AGEMA_signal_6092, new_AGEMA_signal_6096,
         new_AGEMA_signal_6100, new_AGEMA_signal_6104, new_AGEMA_signal_6108,
         new_AGEMA_signal_6112, new_AGEMA_signal_6116, new_AGEMA_signal_6120,
         new_AGEMA_signal_6124, new_AGEMA_signal_6128, new_AGEMA_signal_6132,
         new_AGEMA_signal_6136, new_AGEMA_signal_6140, new_AGEMA_signal_6144,
         new_AGEMA_signal_6148, new_AGEMA_signal_6152, new_AGEMA_signal_6156,
         new_AGEMA_signal_6160, new_AGEMA_signal_6164, new_AGEMA_signal_6168,
         new_AGEMA_signal_6172, new_AGEMA_signal_6176, new_AGEMA_signal_6180,
         new_AGEMA_signal_6184, new_AGEMA_signal_6188, new_AGEMA_signal_6192,
         new_AGEMA_signal_6196, new_AGEMA_signal_6200, new_AGEMA_signal_6204,
         new_AGEMA_signal_6208, new_AGEMA_signal_6212, new_AGEMA_signal_6216,
         new_AGEMA_signal_6220, new_AGEMA_signal_6224, new_AGEMA_signal_6228,
         new_AGEMA_signal_3629, new_AGEMA_signal_3455, new_AGEMA_signal_3637,
         new_AGEMA_signal_3633, new_AGEMA_signal_3464, new_AGEMA_signal_3645,
         new_AGEMA_signal_3641, new_AGEMA_signal_3465, new_AGEMA_signal_3653,
         new_AGEMA_signal_3649, new_AGEMA_signal_3466, new_AGEMA_signal_3661,
         new_AGEMA_signal_3657, new_AGEMA_signal_3467, new_AGEMA_signal_3669,
         new_AGEMA_signal_3665, new_AGEMA_signal_3468, new_AGEMA_signal_3677,
         new_AGEMA_signal_3673, new_AGEMA_signal_3469, new_AGEMA_signal_3685,
         new_AGEMA_signal_3681, new_AGEMA_signal_3470, new_AGEMA_signal_3693,
         new_AGEMA_signal_3689, new_AGEMA_signal_3697, new_AGEMA_signal_3497,
         stateArray_S33reg_gff_1_SFF_0_QD, new_AGEMA_signal_3705,
         new_AGEMA_signal_3701, new_AGEMA_signal_3488, new_AGEMA_signal_3520,
         stateArray_S33reg_gff_1_SFF_1_QD, new_AGEMA_signal_3713,
         new_AGEMA_signal_3709, new_AGEMA_signal_3499, new_AGEMA_signal_3521,
         stateArray_S33reg_gff_1_SFF_2_QD, new_AGEMA_signal_3721,
         new_AGEMA_signal_3717, new_AGEMA_signal_3501, new_AGEMA_signal_3522,
         stateArray_S33reg_gff_1_SFF_3_QD, new_AGEMA_signal_3729,
         new_AGEMA_signal_3725, new_AGEMA_signal_3503, new_AGEMA_signal_3523,
         stateArray_S33reg_gff_1_SFF_4_QD, new_AGEMA_signal_3737,
         new_AGEMA_signal_3733, new_AGEMA_signal_3505, new_AGEMA_signal_3524,
         stateArray_S33reg_gff_1_SFF_5_QD, new_AGEMA_signal_3745,
         new_AGEMA_signal_3741, new_AGEMA_signal_3507, new_AGEMA_signal_3525,
         stateArray_S33reg_gff_1_SFF_6_QD, new_AGEMA_signal_3753,
         new_AGEMA_signal_3749, new_AGEMA_signal_3509, new_AGEMA_signal_3526,
         stateArray_S33reg_gff_1_SFF_7_QD, new_AGEMA_signal_3761,
         new_AGEMA_signal_3757, new_AGEMA_signal_3511, new_AGEMA_signal_3765,
         new_AGEMA_signal_3471, new_AGEMA_signal_3773, new_AGEMA_signal_3769,
         new_AGEMA_signal_3480, new_AGEMA_signal_3781, new_AGEMA_signal_3777,
         new_AGEMA_signal_3481, new_AGEMA_signal_3789, new_AGEMA_signal_3785,
         new_AGEMA_signal_3482, new_AGEMA_signal_3797, new_AGEMA_signal_3793,
         new_AGEMA_signal_3483, new_AGEMA_signal_3805, new_AGEMA_signal_3801,
         new_AGEMA_signal_3484, new_AGEMA_signal_3813, new_AGEMA_signal_3809,
         new_AGEMA_signal_3485, new_AGEMA_signal_3821, new_AGEMA_signal_3817,
         new_AGEMA_signal_3486, new_AGEMA_signal_3829, new_AGEMA_signal_3825,
         new_AGEMA_signal_3833, new_AGEMA_signal_3841, new_AGEMA_signal_3837,
         new_AGEMA_signal_3849, new_AGEMA_signal_3845, new_AGEMA_signal_3857,
         new_AGEMA_signal_3853, new_AGEMA_signal_3865, new_AGEMA_signal_3861,
         new_AGEMA_signal_3873, new_AGEMA_signal_3869, new_AGEMA_signal_3881,
         new_AGEMA_signal_3877, new_AGEMA_signal_3889, new_AGEMA_signal_3885,
         new_AGEMA_signal_3897, new_AGEMA_signal_3893, new_AGEMA_signal_3489,
         new_AGEMA_signal_3905, new_AGEMA_signal_3901, new_AGEMA_signal_3472,
         KeyArray_n55, new_AGEMA_signal_3909, new_AGEMA_signal_3490,
         new_AGEMA_signal_3917, new_AGEMA_signal_3913, new_AGEMA_signal_3473,
         KeyArray_n54, new_AGEMA_signal_3921, new_AGEMA_signal_3491,
         new_AGEMA_signal_3929, new_AGEMA_signal_3925, new_AGEMA_signal_3474,
         KeyArray_n53, new_AGEMA_signal_3933, new_AGEMA_signal_3492,
         new_AGEMA_signal_3941, new_AGEMA_signal_3937, new_AGEMA_signal_3475,
         KeyArray_n52, new_AGEMA_signal_3945, new_AGEMA_signal_3493,
         new_AGEMA_signal_3953, new_AGEMA_signal_3949, new_AGEMA_signal_3476,
         KeyArray_n51, new_AGEMA_signal_3957, new_AGEMA_signal_3494,
         new_AGEMA_signal_3965, new_AGEMA_signal_3961, new_AGEMA_signal_3477,
         KeyArray_n50, new_AGEMA_signal_3969, new_AGEMA_signal_3495,
         new_AGEMA_signal_3977, new_AGEMA_signal_3973, new_AGEMA_signal_3478,
         KeyArray_n49, new_AGEMA_signal_3981, new_AGEMA_signal_3479,
         new_AGEMA_signal_3989, new_AGEMA_signal_3985, new_AGEMA_signal_3456,
         KeyArray_n48, new_AGEMA_signal_3993, new_AGEMA_signal_3997,
         new_AGEMA_signal_3512, KeyArray_S30reg_gff_1_SFF_0_n5,
         new_AGEMA_signal_3496, KeyArray_S30reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_4005, new_AGEMA_signal_4001, new_AGEMA_signal_4009,
         new_AGEMA_signal_4017, new_AGEMA_signal_4013, new_AGEMA_signal_3527,
         KeyArray_S30reg_gff_1_SFF_1_n5, new_AGEMA_signal_3513,
         KeyArray_S30reg_gff_1_SFF_1_QD, new_AGEMA_signal_4025,
         new_AGEMA_signal_4021, new_AGEMA_signal_4033, new_AGEMA_signal_4029,
         new_AGEMA_signal_3528, KeyArray_S30reg_gff_1_SFF_2_n5,
         new_AGEMA_signal_3514, KeyArray_S30reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_4041, new_AGEMA_signal_4037, new_AGEMA_signal_4049,
         new_AGEMA_signal_4045, new_AGEMA_signal_3529,
         KeyArray_S30reg_gff_1_SFF_3_n5, new_AGEMA_signal_3515,
         KeyArray_S30reg_gff_1_SFF_3_QD, new_AGEMA_signal_4057,
         new_AGEMA_signal_4053, new_AGEMA_signal_4065, new_AGEMA_signal_4061,
         new_AGEMA_signal_3530, KeyArray_S30reg_gff_1_SFF_4_n5,
         new_AGEMA_signal_3516, KeyArray_S30reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_4073, new_AGEMA_signal_4069, new_AGEMA_signal_4081,
         new_AGEMA_signal_4077, new_AGEMA_signal_3531,
         KeyArray_S30reg_gff_1_SFF_5_n5, new_AGEMA_signal_3517,
         KeyArray_S30reg_gff_1_SFF_5_QD, new_AGEMA_signal_4089,
         new_AGEMA_signal_4085, new_AGEMA_signal_4097, new_AGEMA_signal_4093,
         new_AGEMA_signal_3532, KeyArray_S30reg_gff_1_SFF_6_n5,
         new_AGEMA_signal_3518, KeyArray_S30reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_4105, new_AGEMA_signal_4101, new_AGEMA_signal_4113,
         new_AGEMA_signal_4109, new_AGEMA_signal_3533,
         KeyArray_S30reg_gff_1_SFF_7_n5, new_AGEMA_signal_3519,
         KeyArray_S30reg_gff_1_SFF_7_QD, new_AGEMA_signal_4121,
         new_AGEMA_signal_4117, new_AGEMA_signal_4129, new_AGEMA_signal_4125,
         new_AGEMA_signal_3414, Inst_bSbox_M46, new_AGEMA_signal_3405,
         Inst_bSbox_M47, new_AGEMA_signal_3406, Inst_bSbox_M48,
         new_AGEMA_signal_3415, Inst_bSbox_M49, new_AGEMA_signal_3407,
         Inst_bSbox_M50, new_AGEMA_signal_3408, Inst_bSbox_M51,
         new_AGEMA_signal_3416, Inst_bSbox_M52, new_AGEMA_signal_3425,
         Inst_bSbox_M53, new_AGEMA_signal_3417, Inst_bSbox_M54,
         new_AGEMA_signal_3418, Inst_bSbox_M55, new_AGEMA_signal_3409,
         Inst_bSbox_M56, new_AGEMA_signal_3410, Inst_bSbox_M57,
         new_AGEMA_signal_3419, Inst_bSbox_M58, new_AGEMA_signal_3411,
         Inst_bSbox_M59, new_AGEMA_signal_3412, Inst_bSbox_M60,
         new_AGEMA_signal_3420, Inst_bSbox_M61, new_AGEMA_signal_3426,
         Inst_bSbox_M62, new_AGEMA_signal_3421, Inst_bSbox_M63,
         new_AGEMA_signal_3435, Inst_bSbox_L0, new_AGEMA_signal_3422,
         Inst_bSbox_L1, new_AGEMA_signal_3427, Inst_bSbox_L2,
         new_AGEMA_signal_3428, Inst_bSbox_L3, new_AGEMA_signal_3429,
         Inst_bSbox_L4, new_AGEMA_signal_3430, Inst_bSbox_L5,
         new_AGEMA_signal_3436, Inst_bSbox_L6, new_AGEMA_signal_3437,
         Inst_bSbox_L7, new_AGEMA_signal_3423, Inst_bSbox_L8,
         new_AGEMA_signal_3438, Inst_bSbox_L9, new_AGEMA_signal_3439,
         Inst_bSbox_L10, new_AGEMA_signal_3440, Inst_bSbox_L11,
         new_AGEMA_signal_3424, Inst_bSbox_L12, new_AGEMA_signal_3444,
         Inst_bSbox_L13, new_AGEMA_signal_3431, Inst_bSbox_L14,
         new_AGEMA_signal_3432, Inst_bSbox_L15, new_AGEMA_signal_3445,
         Inst_bSbox_L16, new_AGEMA_signal_3433, Inst_bSbox_L17,
         new_AGEMA_signal_3434, Inst_bSbox_L18, new_AGEMA_signal_3441,
         Inst_bSbox_L19, new_AGEMA_signal_3446, Inst_bSbox_L20,
         new_AGEMA_signal_3447, Inst_bSbox_L21, new_AGEMA_signal_3442,
         Inst_bSbox_L22, new_AGEMA_signal_3443, Inst_bSbox_L23,
         new_AGEMA_signal_3448, Inst_bSbox_L24, new_AGEMA_signal_3449,
         Inst_bSbox_L25, new_AGEMA_signal_3450, Inst_bSbox_L26,
         new_AGEMA_signal_3451, Inst_bSbox_L27, new_AGEMA_signal_3452,
         Inst_bSbox_L28, new_AGEMA_signal_3453, Inst_bSbox_L29,
         new_AGEMA_signal_4241, new_AGEMA_signal_4245, new_AGEMA_signal_4249,
         new_AGEMA_signal_4253, new_AGEMA_signal_4257, new_AGEMA_signal_4261,
         new_AGEMA_signal_4265, new_AGEMA_signal_4269, new_AGEMA_signal_4273,
         new_AGEMA_signal_4277, new_AGEMA_signal_4281, new_AGEMA_signal_4285,
         new_AGEMA_signal_4289, new_AGEMA_signal_4293, new_AGEMA_signal_4297,
         new_AGEMA_signal_4301, new_AGEMA_signal_4305, new_AGEMA_signal_4309,
         new_AGEMA_signal_4313, new_AGEMA_signal_4317, new_AGEMA_signal_4321,
         new_AGEMA_signal_4325, new_AGEMA_signal_4329, new_AGEMA_signal_4333,
         new_AGEMA_signal_4337, new_AGEMA_signal_4341, new_AGEMA_signal_4345,
         new_AGEMA_signal_4349, new_AGEMA_signal_4353, new_AGEMA_signal_4357,
         new_AGEMA_signal_4361, new_AGEMA_signal_4365, new_AGEMA_signal_4369,
         new_AGEMA_signal_4373, new_AGEMA_signal_4377, new_AGEMA_signal_4381,
         new_AGEMA_signal_4385, new_AGEMA_signal_4389, new_AGEMA_signal_4393,
         new_AGEMA_signal_4397, new_AGEMA_signal_4401, new_AGEMA_signal_4405,
         new_AGEMA_signal_4409, new_AGEMA_signal_4413, new_AGEMA_signal_4417,
         new_AGEMA_signal_4421, new_AGEMA_signal_4425, new_AGEMA_signal_4429,
         new_AGEMA_signal_4433, new_AGEMA_signal_4437, new_AGEMA_signal_4441,
         new_AGEMA_signal_4445, new_AGEMA_signal_4449, new_AGEMA_signal_4453,
         new_AGEMA_signal_4457, new_AGEMA_signal_4461, new_AGEMA_signal_4465,
         new_AGEMA_signal_4469, new_AGEMA_signal_4473, new_AGEMA_signal_4477,
         new_AGEMA_signal_4481, new_AGEMA_signal_4485, new_AGEMA_signal_4489,
         new_AGEMA_signal_4493, new_AGEMA_signal_4497, new_AGEMA_signal_4501,
         new_AGEMA_signal_4505, new_AGEMA_signal_4509, new_AGEMA_signal_4513,
         new_AGEMA_signal_4517, new_AGEMA_signal_4521, new_AGEMA_signal_4525,
         new_AGEMA_signal_4529, new_AGEMA_signal_4533, new_AGEMA_signal_4537,
         new_AGEMA_signal_4541, new_AGEMA_signal_4545, new_AGEMA_signal_4549,
         new_AGEMA_signal_4553, new_AGEMA_signal_4557, new_AGEMA_signal_4561,
         new_AGEMA_signal_4565, new_AGEMA_signal_4569, new_AGEMA_signal_4573,
         new_AGEMA_signal_4577, new_AGEMA_signal_4581, new_AGEMA_signal_4585,
         new_AGEMA_signal_4589, new_AGEMA_signal_4593, new_AGEMA_signal_4597,
         new_AGEMA_signal_4601, new_AGEMA_signal_4605, new_AGEMA_signal_4609,
         new_AGEMA_signal_4613, new_AGEMA_signal_4617, new_AGEMA_signal_4621,
         new_AGEMA_signal_4625, new_AGEMA_signal_4629, new_AGEMA_signal_4633,
         new_AGEMA_signal_4637, new_AGEMA_signal_4641, new_AGEMA_signal_4645,
         new_AGEMA_signal_4649, new_AGEMA_signal_4653, new_AGEMA_signal_4657,
         new_AGEMA_signal_4661, new_AGEMA_signal_4665, new_AGEMA_signal_4669,
         new_AGEMA_signal_4673, new_AGEMA_signal_4677, new_AGEMA_signal_4681,
         new_AGEMA_signal_4685, new_AGEMA_signal_4689, new_AGEMA_signal_4693,
         new_AGEMA_signal_4697, new_AGEMA_signal_4701, new_AGEMA_signal_4705,
         new_AGEMA_signal_4709, new_AGEMA_signal_4713, new_AGEMA_signal_4717,
         new_AGEMA_signal_4721, new_AGEMA_signal_4725, new_AGEMA_signal_4729,
         new_AGEMA_signal_4733, new_AGEMA_signal_4737, new_AGEMA_signal_4741,
         new_AGEMA_signal_4745, new_AGEMA_signal_4749, new_AGEMA_signal_4753,
         new_AGEMA_signal_4757, new_AGEMA_signal_4761, new_AGEMA_signal_4765,
         new_AGEMA_signal_4769, new_AGEMA_signal_4773, new_AGEMA_signal_4777,
         new_AGEMA_signal_4781, new_AGEMA_signal_4785, new_AGEMA_signal_4789,
         new_AGEMA_signal_4793, new_AGEMA_signal_4797, new_AGEMA_signal_4801,
         new_AGEMA_signal_4805, new_AGEMA_signal_4809, new_AGEMA_signal_4813,
         new_AGEMA_signal_4817, new_AGEMA_signal_4821, new_AGEMA_signal_4825,
         new_AGEMA_signal_4829, new_AGEMA_signal_4833, new_AGEMA_signal_4837,
         new_AGEMA_signal_4841, new_AGEMA_signal_4845, new_AGEMA_signal_4849,
         new_AGEMA_signal_4853, new_AGEMA_signal_4857, new_AGEMA_signal_4861,
         new_AGEMA_signal_4865, new_AGEMA_signal_4869, new_AGEMA_signal_4873,
         new_AGEMA_signal_4877, new_AGEMA_signal_4881, new_AGEMA_signal_4885,
         new_AGEMA_signal_4889, new_AGEMA_signal_4893, new_AGEMA_signal_4897,
         new_AGEMA_signal_4901, new_AGEMA_signal_4905, new_AGEMA_signal_4909,
         new_AGEMA_signal_4913, new_AGEMA_signal_4917, new_AGEMA_signal_4921,
         new_AGEMA_signal_4925, new_AGEMA_signal_4929, new_AGEMA_signal_4933,
         new_AGEMA_signal_4937, new_AGEMA_signal_4941, new_AGEMA_signal_4945,
         new_AGEMA_signal_4949, new_AGEMA_signal_4953, new_AGEMA_signal_4957,
         new_AGEMA_signal_4961, new_AGEMA_signal_4965, new_AGEMA_signal_4969,
         new_AGEMA_signal_4973, new_AGEMA_signal_4977, new_AGEMA_signal_4981,
         new_AGEMA_signal_4985, new_AGEMA_signal_4989, new_AGEMA_signal_4993,
         new_AGEMA_signal_4997, new_AGEMA_signal_5001, new_AGEMA_signal_5005,
         new_AGEMA_signal_5009, new_AGEMA_signal_5013, new_AGEMA_signal_5017,
         new_AGEMA_signal_5021, new_AGEMA_signal_5025, new_AGEMA_signal_5029,
         new_AGEMA_signal_5033, new_AGEMA_signal_5037, new_AGEMA_signal_5041,
         new_AGEMA_signal_5045, new_AGEMA_signal_5049, new_AGEMA_signal_5053,
         new_AGEMA_signal_5057, new_AGEMA_signal_5061, new_AGEMA_signal_5065,
         new_AGEMA_signal_5069, new_AGEMA_signal_5073, new_AGEMA_signal_5077,
         new_AGEMA_signal_5081, new_AGEMA_signal_5085, new_AGEMA_signal_5089,
         new_AGEMA_signal_5093, new_AGEMA_signal_5097, new_AGEMA_signal_5101,
         new_AGEMA_signal_5105, new_AGEMA_signal_5109, new_AGEMA_signal_5113,
         new_AGEMA_signal_5117, new_AGEMA_signal_5121, new_AGEMA_signal_5125,
         new_AGEMA_signal_5129, new_AGEMA_signal_5133, new_AGEMA_signal_5137,
         new_AGEMA_signal_5141, new_AGEMA_signal_5145, new_AGEMA_signal_5149,
         new_AGEMA_signal_5153, new_AGEMA_signal_5157, new_AGEMA_signal_5161,
         new_AGEMA_signal_5165, new_AGEMA_signal_5169, new_AGEMA_signal_5173,
         new_AGEMA_signal_5177, new_AGEMA_signal_5181, new_AGEMA_signal_5185,
         new_AGEMA_signal_5189, new_AGEMA_signal_5193, new_AGEMA_signal_5197,
         new_AGEMA_signal_5201, new_AGEMA_signal_5205, new_AGEMA_signal_5209,
         new_AGEMA_signal_5213, new_AGEMA_signal_5217, new_AGEMA_signal_5221,
         new_AGEMA_signal_5225, new_AGEMA_signal_5229, new_AGEMA_signal_5233,
         new_AGEMA_signal_5237, new_AGEMA_signal_5241, new_AGEMA_signal_5245,
         new_AGEMA_signal_5249, new_AGEMA_signal_5253, new_AGEMA_signal_5257,
         new_AGEMA_signal_5261, new_AGEMA_signal_5265, new_AGEMA_signal_5269,
         new_AGEMA_signal_5273, new_AGEMA_signal_5277, new_AGEMA_signal_5281,
         new_AGEMA_signal_5285, new_AGEMA_signal_5289, new_AGEMA_signal_5293,
         new_AGEMA_signal_5297, new_AGEMA_signal_5301, new_AGEMA_signal_5305,
         new_AGEMA_signal_5309, new_AGEMA_signal_5313, new_AGEMA_signal_5317,
         new_AGEMA_signal_5321, new_AGEMA_signal_5325, new_AGEMA_signal_5329,
         new_AGEMA_signal_5333, new_AGEMA_signal_5337, new_AGEMA_signal_5341,
         new_AGEMA_signal_5345, new_AGEMA_signal_5349, new_AGEMA_signal_5353,
         new_AGEMA_signal_5357, new_AGEMA_signal_5361, new_AGEMA_signal_5365,
         new_AGEMA_signal_5369, new_AGEMA_signal_5373, new_AGEMA_signal_5377,
         new_AGEMA_signal_5381, new_AGEMA_signal_5385, new_AGEMA_signal_5389,
         new_AGEMA_signal_5393, new_AGEMA_signal_5397, new_AGEMA_signal_5401,
         new_AGEMA_signal_5405, new_AGEMA_signal_5409, new_AGEMA_signal_5413,
         new_AGEMA_signal_5417, new_AGEMA_signal_5421, new_AGEMA_signal_5425,
         new_AGEMA_signal_5429, new_AGEMA_signal_5433, new_AGEMA_signal_5437,
         new_AGEMA_signal_5441, new_AGEMA_signal_5445, new_AGEMA_signal_5449,
         new_AGEMA_signal_5453, new_AGEMA_signal_5457, new_AGEMA_signal_5461,
         new_AGEMA_signal_5465, new_AGEMA_signal_5469, new_AGEMA_signal_5473,
         new_AGEMA_signal_5477, new_AGEMA_signal_5481, new_AGEMA_signal_5485,
         new_AGEMA_signal_5489, new_AGEMA_signal_5493, new_AGEMA_signal_5497,
         new_AGEMA_signal_5501, new_AGEMA_signal_5505, new_AGEMA_signal_5509,
         new_AGEMA_signal_5513, new_AGEMA_signal_5517, new_AGEMA_signal_5521,
         new_AGEMA_signal_5525, new_AGEMA_signal_5529, new_AGEMA_signal_5533,
         new_AGEMA_signal_5537, new_AGEMA_signal_5541, new_AGEMA_signal_5545,
         new_AGEMA_signal_5549, new_AGEMA_signal_5553, new_AGEMA_signal_5557,
         new_AGEMA_signal_5561, new_AGEMA_signal_5565, new_AGEMA_signal_5569,
         new_AGEMA_signal_5573, new_AGEMA_signal_5577, new_AGEMA_signal_5581,
         new_AGEMA_signal_5585, new_AGEMA_signal_5589, new_AGEMA_signal_5593,
         new_AGEMA_signal_5597, new_AGEMA_signal_5601, new_AGEMA_signal_5605,
         new_AGEMA_signal_5609, new_AGEMA_signal_5613, new_AGEMA_signal_5617,
         new_AGEMA_signal_5621, new_AGEMA_signal_5625, new_AGEMA_signal_5629,
         new_AGEMA_signal_5633, new_AGEMA_signal_5637, new_AGEMA_signal_5641,
         new_AGEMA_signal_5645, new_AGEMA_signal_5649, new_AGEMA_signal_5653,
         new_AGEMA_signal_5657, new_AGEMA_signal_5661, new_AGEMA_signal_5665,
         new_AGEMA_signal_5669, new_AGEMA_signal_5673, new_AGEMA_signal_5677,
         new_AGEMA_signal_5681, new_AGEMA_signal_5685, new_AGEMA_signal_5689,
         new_AGEMA_signal_5693, new_AGEMA_signal_5697, new_AGEMA_signal_5701,
         new_AGEMA_signal_5705, new_AGEMA_signal_5709, new_AGEMA_signal_5713,
         new_AGEMA_signal_5717, new_AGEMA_signal_5721, new_AGEMA_signal_5725,
         new_AGEMA_signal_5729, new_AGEMA_signal_5733, new_AGEMA_signal_5737,
         new_AGEMA_signal_5741, new_AGEMA_signal_5745, new_AGEMA_signal_5749,
         new_AGEMA_signal_5753, new_AGEMA_signal_5757, new_AGEMA_signal_5761,
         new_AGEMA_signal_5765, new_AGEMA_signal_5769, new_AGEMA_signal_5773,
         new_AGEMA_signal_5777, new_AGEMA_signal_5781, new_AGEMA_signal_5785,
         new_AGEMA_signal_5789, new_AGEMA_signal_5793, new_AGEMA_signal_5797,
         new_AGEMA_signal_5801, new_AGEMA_signal_5805, new_AGEMA_signal_5809,
         new_AGEMA_signal_5813, new_AGEMA_signal_5817, new_AGEMA_signal_5821,
         new_AGEMA_signal_5825, new_AGEMA_signal_5829, new_AGEMA_signal_5833,
         new_AGEMA_signal_5837, new_AGEMA_signal_5841, new_AGEMA_signal_5845,
         new_AGEMA_signal_5849, new_AGEMA_signal_5853, new_AGEMA_signal_5857,
         new_AGEMA_signal_5861, new_AGEMA_signal_5865, new_AGEMA_signal_5869,
         new_AGEMA_signal_5873, new_AGEMA_signal_5877, new_AGEMA_signal_5881,
         new_AGEMA_signal_5885, new_AGEMA_signal_5889, new_AGEMA_signal_5893,
         new_AGEMA_signal_5897, new_AGEMA_signal_5901, new_AGEMA_signal_5905,
         new_AGEMA_signal_5909, new_AGEMA_signal_5913, new_AGEMA_signal_5917,
         new_AGEMA_signal_5921, new_AGEMA_signal_5925, new_AGEMA_signal_5929,
         new_AGEMA_signal_5933, new_AGEMA_signal_5937, new_AGEMA_signal_5941,
         new_AGEMA_signal_5945, new_AGEMA_signal_5949, new_AGEMA_signal_5953,
         new_AGEMA_signal_5957, new_AGEMA_signal_5961, new_AGEMA_signal_5965,
         new_AGEMA_signal_5969, new_AGEMA_signal_5973, new_AGEMA_signal_5977,
         new_AGEMA_signal_5981, new_AGEMA_signal_5985, new_AGEMA_signal_5989,
         new_AGEMA_signal_5993, new_AGEMA_signal_5997, new_AGEMA_signal_6001,
         new_AGEMA_signal_6005, new_AGEMA_signal_6009, new_AGEMA_signal_6013,
         new_AGEMA_signal_6017, new_AGEMA_signal_6021, new_AGEMA_signal_6025,
         new_AGEMA_signal_6029, new_AGEMA_signal_6033, new_AGEMA_signal_6037,
         new_AGEMA_signal_6041, new_AGEMA_signal_6045, new_AGEMA_signal_6049,
         new_AGEMA_signal_6053, new_AGEMA_signal_6057, new_AGEMA_signal_6061,
         new_AGEMA_signal_6065, new_AGEMA_signal_6069, new_AGEMA_signal_6073,
         new_AGEMA_signal_6077, new_AGEMA_signal_6081, new_AGEMA_signal_6085,
         new_AGEMA_signal_6089, new_AGEMA_signal_6093, new_AGEMA_signal_6097,
         new_AGEMA_signal_6101, new_AGEMA_signal_6105, new_AGEMA_signal_6109,
         new_AGEMA_signal_6113, new_AGEMA_signal_6117, new_AGEMA_signal_6121,
         new_AGEMA_signal_6125, new_AGEMA_signal_6129, new_AGEMA_signal_6133,
         new_AGEMA_signal_6137, new_AGEMA_signal_6141, new_AGEMA_signal_6145,
         new_AGEMA_signal_6149, new_AGEMA_signal_6153, new_AGEMA_signal_6157,
         new_AGEMA_signal_6161, new_AGEMA_signal_6165, new_AGEMA_signal_6169,
         new_AGEMA_signal_6173, new_AGEMA_signal_6177, new_AGEMA_signal_6181,
         new_AGEMA_signal_6185, new_AGEMA_signal_6189, new_AGEMA_signal_6193,
         new_AGEMA_signal_6197, new_AGEMA_signal_6201, new_AGEMA_signal_6205,
         new_AGEMA_signal_6209, new_AGEMA_signal_6213, new_AGEMA_signal_6217,
         new_AGEMA_signal_6221, new_AGEMA_signal_6225, new_AGEMA_signal_6229,
         n14, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n55, n56, n57,
         n58, n59, n66, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n4,
         stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n3,
         stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n2,
         stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_0_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_0_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_0_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_0_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_0_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_0_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_1_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_1_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_1_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_1_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_1_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_1_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_2_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_2_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_2_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_2_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_2_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_2_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_3_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_3_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_3_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_3_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_3_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_3_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_4_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_4_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_4_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_4_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_4_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_4_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_5_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_5_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_5_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_5_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_5_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_5_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_6_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_6_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_6_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_6_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_6_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_6_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_7_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_7_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_7_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_7_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_7_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_7_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_8_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_8_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_8_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_8_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_8_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_8_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_9_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_9_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_9_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_9_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_9_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_9_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_10_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_10_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_10_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_10_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_10_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_10_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_11_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_11_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_11_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_11_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_11_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_11_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_12_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_12_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_12_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_12_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_12_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_12_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_13_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_13_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_13_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_13_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_13_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_13_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_14_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_14_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_14_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_14_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_14_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_14_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_15_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_15_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_15_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_15_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_15_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_15_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_16_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_16_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_16_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_16_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_16_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_16_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_17_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_17_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_17_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_17_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_17_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_17_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_18_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_18_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_18_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_18_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_18_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_18_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_19_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_19_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_19_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_19_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_19_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_19_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_20_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_20_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_20_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_20_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_20_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_20_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_21_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_21_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_21_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_21_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_21_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_21_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_22_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_22_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_22_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_22_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_22_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_22_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_23_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_23_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_23_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_23_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_23_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_23_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_24_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_24_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_24_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_24_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_24_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_24_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_25_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_25_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_25_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_25_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_25_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_25_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_26_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_26_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_26_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_26_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_26_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_26_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_27_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_27_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_27_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_27_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_27_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_27_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_28_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_28_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_28_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_28_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_28_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_28_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_29_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_29_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_29_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_29_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_29_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_29_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_30_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_30_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_30_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_30_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_30_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_30_U1_Ins_1_n6,
         MUX_StateInMC_mux_inst_31_U1_Ins_0_n8,
         MUX_StateInMC_mux_inst_31_U1_Ins_0_n7,
         MUX_StateInMC_mux_inst_31_U1_Ins_0_n6,
         MUX_StateInMC_mux_inst_31_U1_Ins_1_n8,
         MUX_StateInMC_mux_inst_31_U1_Ins_1_n7,
         MUX_StateInMC_mux_inst_31_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n8,
         KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n7,
         KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n6,
         KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n8,
         KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n7,
         KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n6,
         KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n8,
         KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n7,
         KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n6,
         KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n8,
         KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n7,
         KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n6,
         KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n8,
         KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n7,
         KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n6,
         KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n8,
         KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n7,
         KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n6,
         KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n8,
         KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n7,
         KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n6,
         KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n8,
         KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n7,
         KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n6,
         KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n8,
         KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n7,
         KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n6,
         KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n8,
         KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n7,
         KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n6,
         KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n8,
         KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n7,
         KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n6,
         KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n8,
         KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n7,
         KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n6,
         KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n8,
         KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n7,
         KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n6,
         KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n8,
         KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n7,
         KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n6,
         KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n8,
         KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n7,
         KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n6,
         KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n8,
         KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n7,
         KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n6,
         MUX_SboxIn_mux_inst_0_U1_Ins_0_n8, MUX_SboxIn_mux_inst_0_U1_Ins_0_n7,
         MUX_SboxIn_mux_inst_0_U1_Ins_0_n6, MUX_SboxIn_mux_inst_0_U1_Ins_1_n8,
         MUX_SboxIn_mux_inst_0_U1_Ins_1_n7, MUX_SboxIn_mux_inst_0_U1_Ins_1_n6,
         MUX_SboxIn_mux_inst_1_U1_Ins_0_n8, MUX_SboxIn_mux_inst_1_U1_Ins_0_n7,
         MUX_SboxIn_mux_inst_1_U1_Ins_0_n6, MUX_SboxIn_mux_inst_1_U1_Ins_1_n8,
         MUX_SboxIn_mux_inst_1_U1_Ins_1_n7, MUX_SboxIn_mux_inst_1_U1_Ins_1_n6,
         MUX_SboxIn_mux_inst_2_U1_Ins_0_n8, MUX_SboxIn_mux_inst_2_U1_Ins_0_n7,
         MUX_SboxIn_mux_inst_2_U1_Ins_0_n6, MUX_SboxIn_mux_inst_2_U1_Ins_1_n8,
         MUX_SboxIn_mux_inst_2_U1_Ins_1_n7, MUX_SboxIn_mux_inst_2_U1_Ins_1_n6,
         MUX_SboxIn_mux_inst_3_U1_Ins_0_n8, MUX_SboxIn_mux_inst_3_U1_Ins_0_n7,
         MUX_SboxIn_mux_inst_3_U1_Ins_0_n6, MUX_SboxIn_mux_inst_3_U1_Ins_1_n8,
         MUX_SboxIn_mux_inst_3_U1_Ins_1_n7, MUX_SboxIn_mux_inst_3_U1_Ins_1_n6,
         MUX_SboxIn_mux_inst_4_U1_Ins_0_n8, MUX_SboxIn_mux_inst_4_U1_Ins_0_n7,
         MUX_SboxIn_mux_inst_4_U1_Ins_0_n6, MUX_SboxIn_mux_inst_4_U1_Ins_1_n8,
         MUX_SboxIn_mux_inst_4_U1_Ins_1_n7, MUX_SboxIn_mux_inst_4_U1_Ins_1_n6,
         MUX_SboxIn_mux_inst_5_U1_Ins_0_n8, MUX_SboxIn_mux_inst_5_U1_Ins_0_n7,
         MUX_SboxIn_mux_inst_5_U1_Ins_0_n6, MUX_SboxIn_mux_inst_5_U1_Ins_1_n8,
         MUX_SboxIn_mux_inst_5_U1_Ins_1_n7, MUX_SboxIn_mux_inst_5_U1_Ins_1_n6,
         MUX_SboxIn_mux_inst_6_U1_Ins_0_n8, MUX_SboxIn_mux_inst_6_U1_Ins_0_n7,
         MUX_SboxIn_mux_inst_6_U1_Ins_0_n6, MUX_SboxIn_mux_inst_6_U1_Ins_1_n8,
         MUX_SboxIn_mux_inst_6_U1_Ins_1_n7, MUX_SboxIn_mux_inst_6_U1_Ins_1_n6,
         MUX_SboxIn_mux_inst_7_U1_Ins_0_n8, MUX_SboxIn_mux_inst_7_U1_Ins_0_n7,
         MUX_SboxIn_mux_inst_7_U1_Ins_0_n6, MUX_SboxIn_mux_inst_7_U1_Ins_1_n8,
         MUX_SboxIn_mux_inst_7_U1_Ins_1_n7, MUX_SboxIn_mux_inst_7_U1_Ins_1_n6,
         Inst_bSbox_AND_M1_U1_n7, Inst_bSbox_AND_M1_U1_n6,
         Inst_bSbox_AND_M1_U1_n5, Inst_bSbox_AND_M1_U1_n4,
         Inst_bSbox_AND_M1_U1_n3, Inst_bSbox_AND_M1_U1_n2,
         Inst_bSbox_AND_M1_U1_n1, Inst_bSbox_AND_M1_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M1_U1_p_0_out_1__0_, Inst_bSbox_AND_M1_U1_s_out_0__1_,
         Inst_bSbox_AND_M1_U1_s_out_1__0_, Inst_bSbox_AND_M1_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M1_U1_p_0_in_1__0_, Inst_bSbox_AND_M1_U1_s_in_0__1_,
         Inst_bSbox_AND_M1_U1_s_in_1__0_, Inst_bSbox_AND_M2_U1_n23,
         Inst_bSbox_AND_M2_U1_n22, Inst_bSbox_AND_M2_U1_n21,
         Inst_bSbox_AND_M2_U1_n20, Inst_bSbox_AND_M2_U1_n19,
         Inst_bSbox_AND_M2_U1_n18, Inst_bSbox_AND_M2_U1_n17,
         Inst_bSbox_AND_M2_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M2_U1_p_0_out_1__0_, Inst_bSbox_AND_M2_U1_s_out_0__1_,
         Inst_bSbox_AND_M2_U1_s_out_1__0_, Inst_bSbox_AND_M2_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M2_U1_p_0_in_1__0_, Inst_bSbox_AND_M2_U1_s_in_0__1_,
         Inst_bSbox_AND_M2_U1_s_in_1__0_, Inst_bSbox_AND_M4_U1_n23,
         Inst_bSbox_AND_M4_U1_n22, Inst_bSbox_AND_M4_U1_n21,
         Inst_bSbox_AND_M4_U1_n20, Inst_bSbox_AND_M4_U1_n19,
         Inst_bSbox_AND_M4_U1_n18, Inst_bSbox_AND_M4_U1_n17,
         Inst_bSbox_AND_M4_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M4_U1_p_0_out_1__0_, Inst_bSbox_AND_M4_U1_s_out_0__1_,
         Inst_bSbox_AND_M4_U1_s_out_1__0_, Inst_bSbox_AND_M4_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M4_U1_p_0_in_1__0_, Inst_bSbox_AND_M4_U1_s_in_0__1_,
         Inst_bSbox_AND_M4_U1_s_in_1__0_, Inst_bSbox_AND_M6_U1_n23,
         Inst_bSbox_AND_M6_U1_n22, Inst_bSbox_AND_M6_U1_n21,
         Inst_bSbox_AND_M6_U1_n20, Inst_bSbox_AND_M6_U1_n19,
         Inst_bSbox_AND_M6_U1_n18, Inst_bSbox_AND_M6_U1_n17,
         Inst_bSbox_AND_M6_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M6_U1_p_0_out_1__0_, Inst_bSbox_AND_M6_U1_s_out_0__1_,
         Inst_bSbox_AND_M6_U1_s_out_1__0_, Inst_bSbox_AND_M6_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M6_U1_p_0_in_1__0_, Inst_bSbox_AND_M6_U1_s_in_0__1_,
         Inst_bSbox_AND_M6_U1_s_in_1__0_, Inst_bSbox_AND_M7_U1_n23,
         Inst_bSbox_AND_M7_U1_n22, Inst_bSbox_AND_M7_U1_n21,
         Inst_bSbox_AND_M7_U1_n20, Inst_bSbox_AND_M7_U1_n19,
         Inst_bSbox_AND_M7_U1_n18, Inst_bSbox_AND_M7_U1_n17,
         Inst_bSbox_AND_M7_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M7_U1_p_0_out_1__0_, Inst_bSbox_AND_M7_U1_s_out_0__1_,
         Inst_bSbox_AND_M7_U1_s_out_1__0_, Inst_bSbox_AND_M7_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M7_U1_p_0_in_1__0_, Inst_bSbox_AND_M7_U1_s_in_0__1_,
         Inst_bSbox_AND_M7_U1_s_in_1__0_, Inst_bSbox_AND_M9_U1_n23,
         Inst_bSbox_AND_M9_U1_n22, Inst_bSbox_AND_M9_U1_n21,
         Inst_bSbox_AND_M9_U1_n20, Inst_bSbox_AND_M9_U1_n19,
         Inst_bSbox_AND_M9_U1_n18, Inst_bSbox_AND_M9_U1_n17,
         Inst_bSbox_AND_M9_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M9_U1_p_0_out_1__0_, Inst_bSbox_AND_M9_U1_s_out_0__1_,
         Inst_bSbox_AND_M9_U1_s_out_1__0_, Inst_bSbox_AND_M9_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M9_U1_p_0_in_1__0_, Inst_bSbox_AND_M9_U1_s_in_0__1_,
         Inst_bSbox_AND_M9_U1_s_in_1__0_, Inst_bSbox_AND_M11_U1_n23,
         Inst_bSbox_AND_M11_U1_n22, Inst_bSbox_AND_M11_U1_n21,
         Inst_bSbox_AND_M11_U1_n20, Inst_bSbox_AND_M11_U1_n19,
         Inst_bSbox_AND_M11_U1_n18, Inst_bSbox_AND_M11_U1_n17,
         Inst_bSbox_AND_M11_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M11_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M11_U1_s_out_0__1_, Inst_bSbox_AND_M11_U1_s_out_1__0_,
         Inst_bSbox_AND_M11_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M11_U1_p_0_in_1__0_, Inst_bSbox_AND_M11_U1_s_in_0__1_,
         Inst_bSbox_AND_M11_U1_s_in_1__0_, Inst_bSbox_AND_M12_U1_n23,
         Inst_bSbox_AND_M12_U1_n22, Inst_bSbox_AND_M12_U1_n21,
         Inst_bSbox_AND_M12_U1_n20, Inst_bSbox_AND_M12_U1_n19,
         Inst_bSbox_AND_M12_U1_n18, Inst_bSbox_AND_M12_U1_n17,
         Inst_bSbox_AND_M12_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M12_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M12_U1_s_out_0__1_, Inst_bSbox_AND_M12_U1_s_out_1__0_,
         Inst_bSbox_AND_M12_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M12_U1_p_0_in_1__0_, Inst_bSbox_AND_M12_U1_s_in_0__1_,
         Inst_bSbox_AND_M12_U1_s_in_1__0_, Inst_bSbox_AND_M14_U1_n23,
         Inst_bSbox_AND_M14_U1_n22, Inst_bSbox_AND_M14_U1_n21,
         Inst_bSbox_AND_M14_U1_n20, Inst_bSbox_AND_M14_U1_n19,
         Inst_bSbox_AND_M14_U1_n18, Inst_bSbox_AND_M14_U1_n17,
         Inst_bSbox_AND_M14_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M14_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M14_U1_s_out_0__1_, Inst_bSbox_AND_M14_U1_s_out_1__0_,
         Inst_bSbox_AND_M14_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M14_U1_p_0_in_1__0_, Inst_bSbox_AND_M14_U1_s_in_0__1_,
         Inst_bSbox_AND_M14_U1_s_in_1__0_, Inst_bSbox_AND_M25_U1_n23,
         Inst_bSbox_AND_M25_U1_n22, Inst_bSbox_AND_M25_U1_n21,
         Inst_bSbox_AND_M25_U1_n20, Inst_bSbox_AND_M25_U1_n19,
         Inst_bSbox_AND_M25_U1_n18, Inst_bSbox_AND_M25_U1_n17,
         Inst_bSbox_AND_M25_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M25_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M25_U1_s_out_0__1_, Inst_bSbox_AND_M25_U1_s_out_1__0_,
         Inst_bSbox_AND_M25_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M25_U1_p_0_in_1__0_, Inst_bSbox_AND_M25_U1_s_in_0__1_,
         Inst_bSbox_AND_M25_U1_s_in_1__0_, Inst_bSbox_AND_M31_U1_n23,
         Inst_bSbox_AND_M31_U1_n22, Inst_bSbox_AND_M31_U1_n21,
         Inst_bSbox_AND_M31_U1_n20, Inst_bSbox_AND_M31_U1_n19,
         Inst_bSbox_AND_M31_U1_n18, Inst_bSbox_AND_M31_U1_n17,
         Inst_bSbox_AND_M31_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M31_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M31_U1_s_out_0__1_, Inst_bSbox_AND_M31_U1_s_out_1__0_,
         Inst_bSbox_AND_M31_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M31_U1_p_0_in_1__0_, Inst_bSbox_AND_M31_U1_s_in_0__1_,
         Inst_bSbox_AND_M31_U1_s_in_1__0_, Inst_bSbox_AND_M34_U1_n23,
         Inst_bSbox_AND_M34_U1_n22, Inst_bSbox_AND_M34_U1_n21,
         Inst_bSbox_AND_M34_U1_n20, Inst_bSbox_AND_M34_U1_n19,
         Inst_bSbox_AND_M34_U1_n18, Inst_bSbox_AND_M34_U1_n17,
         Inst_bSbox_AND_M34_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M34_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M34_U1_s_out_0__1_, Inst_bSbox_AND_M34_U1_s_out_1__0_,
         Inst_bSbox_AND_M34_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M34_U1_p_0_in_1__0_, Inst_bSbox_AND_M34_U1_s_in_0__1_,
         Inst_bSbox_AND_M34_U1_s_in_1__0_, Inst_bSbox_AND_M29_U1_n23,
         Inst_bSbox_AND_M29_U1_n22, Inst_bSbox_AND_M29_U1_n21,
         Inst_bSbox_AND_M29_U1_n20, Inst_bSbox_AND_M29_U1_n19,
         Inst_bSbox_AND_M29_U1_n18, Inst_bSbox_AND_M29_U1_n17,
         Inst_bSbox_AND_M29_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M29_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M29_U1_s_out_0__1_, Inst_bSbox_AND_M29_U1_s_out_1__0_,
         Inst_bSbox_AND_M29_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M29_U1_p_0_in_1__0_, Inst_bSbox_AND_M29_U1_s_in_0__1_,
         Inst_bSbox_AND_M29_U1_s_in_1__0_, Inst_bSbox_AND_M30_U1_n23,
         Inst_bSbox_AND_M30_U1_n22, Inst_bSbox_AND_M30_U1_n21,
         Inst_bSbox_AND_M30_U1_n20, Inst_bSbox_AND_M30_U1_n19,
         Inst_bSbox_AND_M30_U1_n18, Inst_bSbox_AND_M30_U1_n17,
         Inst_bSbox_AND_M30_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M30_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M30_U1_s_out_0__1_, Inst_bSbox_AND_M30_U1_s_out_1__0_,
         Inst_bSbox_AND_M30_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M30_U1_p_0_in_1__0_, Inst_bSbox_AND_M30_U1_s_in_0__1_,
         Inst_bSbox_AND_M30_U1_s_in_1__0_, Inst_bSbox_AND_M32_U1_n23,
         Inst_bSbox_AND_M32_U1_n22, Inst_bSbox_AND_M32_U1_n21,
         Inst_bSbox_AND_M32_U1_n20, Inst_bSbox_AND_M32_U1_n19,
         Inst_bSbox_AND_M32_U1_n18, Inst_bSbox_AND_M32_U1_n17,
         Inst_bSbox_AND_M32_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M32_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M32_U1_s_out_0__1_, Inst_bSbox_AND_M32_U1_s_out_1__0_,
         Inst_bSbox_AND_M32_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M32_U1_p_0_in_1__0_, Inst_bSbox_AND_M32_U1_s_in_0__1_,
         Inst_bSbox_AND_M32_U1_s_in_1__0_, Inst_bSbox_AND_M35_U1_n23,
         Inst_bSbox_AND_M35_U1_n22, Inst_bSbox_AND_M35_U1_n21,
         Inst_bSbox_AND_M35_U1_n20, Inst_bSbox_AND_M35_U1_n19,
         Inst_bSbox_AND_M35_U1_n18, Inst_bSbox_AND_M35_U1_n17,
         Inst_bSbox_AND_M35_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M35_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M35_U1_s_out_0__1_, Inst_bSbox_AND_M35_U1_s_out_1__0_,
         Inst_bSbox_AND_M35_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M35_U1_p_0_in_1__0_, Inst_bSbox_AND_M35_U1_s_in_0__1_,
         Inst_bSbox_AND_M35_U1_s_in_1__0_, MUX_StateIn_mux_inst_0_U1_Ins_0_n8,
         MUX_StateIn_mux_inst_0_U1_Ins_0_n7,
         MUX_StateIn_mux_inst_0_U1_Ins_0_n6,
         MUX_StateIn_mux_inst_0_U1_Ins_1_n8,
         MUX_StateIn_mux_inst_0_U1_Ins_1_n7,
         MUX_StateIn_mux_inst_0_U1_Ins_1_n6,
         MUX_StateIn_mux_inst_1_U1_Ins_0_n8,
         MUX_StateIn_mux_inst_1_U1_Ins_0_n7,
         MUX_StateIn_mux_inst_1_U1_Ins_0_n6,
         MUX_StateIn_mux_inst_1_U1_Ins_1_n8,
         MUX_StateIn_mux_inst_1_U1_Ins_1_n7,
         MUX_StateIn_mux_inst_1_U1_Ins_1_n6,
         MUX_StateIn_mux_inst_2_U1_Ins_0_n8,
         MUX_StateIn_mux_inst_2_U1_Ins_0_n7,
         MUX_StateIn_mux_inst_2_U1_Ins_0_n6,
         MUX_StateIn_mux_inst_2_U1_Ins_1_n8,
         MUX_StateIn_mux_inst_2_U1_Ins_1_n7,
         MUX_StateIn_mux_inst_2_U1_Ins_1_n6,
         MUX_StateIn_mux_inst_3_U1_Ins_0_n8,
         MUX_StateIn_mux_inst_3_U1_Ins_0_n7,
         MUX_StateIn_mux_inst_3_U1_Ins_0_n6,
         MUX_StateIn_mux_inst_3_U1_Ins_1_n8,
         MUX_StateIn_mux_inst_3_U1_Ins_1_n7,
         MUX_StateIn_mux_inst_3_U1_Ins_1_n6,
         MUX_StateIn_mux_inst_4_U1_Ins_0_n8,
         MUX_StateIn_mux_inst_4_U1_Ins_0_n7,
         MUX_StateIn_mux_inst_4_U1_Ins_0_n6,
         MUX_StateIn_mux_inst_4_U1_Ins_1_n8,
         MUX_StateIn_mux_inst_4_U1_Ins_1_n7,
         MUX_StateIn_mux_inst_4_U1_Ins_1_n6,
         MUX_StateIn_mux_inst_5_U1_Ins_0_n8,
         MUX_StateIn_mux_inst_5_U1_Ins_0_n7,
         MUX_StateIn_mux_inst_5_U1_Ins_0_n6,
         MUX_StateIn_mux_inst_5_U1_Ins_1_n8,
         MUX_StateIn_mux_inst_5_U1_Ins_1_n7,
         MUX_StateIn_mux_inst_5_U1_Ins_1_n6,
         MUX_StateIn_mux_inst_6_U1_Ins_0_n8,
         MUX_StateIn_mux_inst_6_U1_Ins_0_n7,
         MUX_StateIn_mux_inst_6_U1_Ins_0_n6,
         MUX_StateIn_mux_inst_6_U1_Ins_1_n8,
         MUX_StateIn_mux_inst_6_U1_Ins_1_n7,
         MUX_StateIn_mux_inst_6_U1_Ins_1_n6,
         MUX_StateIn_mux_inst_7_U1_Ins_0_n8,
         MUX_StateIn_mux_inst_7_U1_Ins_0_n7,
         MUX_StateIn_mux_inst_7_U1_Ins_0_n6,
         MUX_StateIn_mux_inst_7_U1_Ins_1_n8,
         MUX_StateIn_mux_inst_7_U1_Ins_1_n7,
         MUX_StateIn_mux_inst_7_U1_Ins_1_n6,
         stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_n6,
         stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n8,
         stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n7,
         stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n6,
         stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n8,
         stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n7,
         stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n6,
         stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n8,
         stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n7,
         stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n6,
         stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n8,
         stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n7,
         stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n6,
         stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n8,
         stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n7,
         stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n6,
         stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n8,
         stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n7,
         stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n6,
         stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n8,
         stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n7,
         stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n6,
         stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n8,
         stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n7,
         stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n6,
         stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n8,
         stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n7,
         stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n6,
         stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n8,
         stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n7,
         stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n6,
         stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n8,
         stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n7,
         stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n6,
         stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n8,
         stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n7,
         stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n6,
         stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n8,
         stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n7,
         stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n6,
         stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n8,
         stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n7,
         stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n6,
         stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n8,
         stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n7,
         stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n6,
         stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n8,
         stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n7,
         stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_n6,
         KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8,
         KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7,
         KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6,
         KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8,
         KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7,
         KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6,
         Inst_bSbox_AND_M46_U1_n23, Inst_bSbox_AND_M46_U1_n22,
         Inst_bSbox_AND_M46_U1_n21, Inst_bSbox_AND_M46_U1_n20,
         Inst_bSbox_AND_M46_U1_n19, Inst_bSbox_AND_M46_U1_n18,
         Inst_bSbox_AND_M46_U1_n17, Inst_bSbox_AND_M46_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M46_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M46_U1_s_out_0__1_, Inst_bSbox_AND_M46_U1_s_out_1__0_,
         Inst_bSbox_AND_M46_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M46_U1_p_0_in_1__0_, Inst_bSbox_AND_M46_U1_s_in_0__1_,
         Inst_bSbox_AND_M46_U1_s_in_1__0_, Inst_bSbox_AND_M47_U1_n23,
         Inst_bSbox_AND_M47_U1_n22, Inst_bSbox_AND_M47_U1_n21,
         Inst_bSbox_AND_M47_U1_n20, Inst_bSbox_AND_M47_U1_n19,
         Inst_bSbox_AND_M47_U1_n18, Inst_bSbox_AND_M47_U1_n17,
         Inst_bSbox_AND_M47_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M47_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M47_U1_s_out_0__1_, Inst_bSbox_AND_M47_U1_s_out_1__0_,
         Inst_bSbox_AND_M47_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M47_U1_p_0_in_1__0_, Inst_bSbox_AND_M47_U1_s_in_0__1_,
         Inst_bSbox_AND_M47_U1_s_in_1__0_, Inst_bSbox_AND_M48_U1_n23,
         Inst_bSbox_AND_M48_U1_n22, Inst_bSbox_AND_M48_U1_n21,
         Inst_bSbox_AND_M48_U1_n20, Inst_bSbox_AND_M48_U1_n19,
         Inst_bSbox_AND_M48_U1_n18, Inst_bSbox_AND_M48_U1_n17,
         Inst_bSbox_AND_M48_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M48_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M48_U1_s_out_0__1_, Inst_bSbox_AND_M48_U1_s_out_1__0_,
         Inst_bSbox_AND_M48_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M48_U1_p_0_in_1__0_, Inst_bSbox_AND_M48_U1_s_in_0__1_,
         Inst_bSbox_AND_M48_U1_s_in_1__0_, Inst_bSbox_AND_M49_U1_n23,
         Inst_bSbox_AND_M49_U1_n22, Inst_bSbox_AND_M49_U1_n21,
         Inst_bSbox_AND_M49_U1_n20, Inst_bSbox_AND_M49_U1_n19,
         Inst_bSbox_AND_M49_U1_n18, Inst_bSbox_AND_M49_U1_n17,
         Inst_bSbox_AND_M49_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M49_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M49_U1_s_out_0__1_, Inst_bSbox_AND_M49_U1_s_out_1__0_,
         Inst_bSbox_AND_M49_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M49_U1_p_0_in_1__0_, Inst_bSbox_AND_M49_U1_s_in_0__1_,
         Inst_bSbox_AND_M49_U1_s_in_1__0_, Inst_bSbox_AND_M50_U1_n23,
         Inst_bSbox_AND_M50_U1_n22, Inst_bSbox_AND_M50_U1_n21,
         Inst_bSbox_AND_M50_U1_n20, Inst_bSbox_AND_M50_U1_n19,
         Inst_bSbox_AND_M50_U1_n18, Inst_bSbox_AND_M50_U1_n17,
         Inst_bSbox_AND_M50_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M50_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M50_U1_s_out_0__1_, Inst_bSbox_AND_M50_U1_s_out_1__0_,
         Inst_bSbox_AND_M50_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M50_U1_p_0_in_1__0_, Inst_bSbox_AND_M50_U1_s_in_0__1_,
         Inst_bSbox_AND_M50_U1_s_in_1__0_, Inst_bSbox_AND_M51_U1_n23,
         Inst_bSbox_AND_M51_U1_n22, Inst_bSbox_AND_M51_U1_n21,
         Inst_bSbox_AND_M51_U1_n20, Inst_bSbox_AND_M51_U1_n19,
         Inst_bSbox_AND_M51_U1_n18, Inst_bSbox_AND_M51_U1_n17,
         Inst_bSbox_AND_M51_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M51_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M51_U1_s_out_0__1_, Inst_bSbox_AND_M51_U1_s_out_1__0_,
         Inst_bSbox_AND_M51_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M51_U1_p_0_in_1__0_, Inst_bSbox_AND_M51_U1_s_in_0__1_,
         Inst_bSbox_AND_M51_U1_s_in_1__0_, Inst_bSbox_AND_M52_U1_n23,
         Inst_bSbox_AND_M52_U1_n22, Inst_bSbox_AND_M52_U1_n21,
         Inst_bSbox_AND_M52_U1_n20, Inst_bSbox_AND_M52_U1_n19,
         Inst_bSbox_AND_M52_U1_n18, Inst_bSbox_AND_M52_U1_n17,
         Inst_bSbox_AND_M52_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M52_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M52_U1_s_out_0__1_, Inst_bSbox_AND_M52_U1_s_out_1__0_,
         Inst_bSbox_AND_M52_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M52_U1_p_0_in_1__0_, Inst_bSbox_AND_M52_U1_s_in_0__1_,
         Inst_bSbox_AND_M52_U1_s_in_1__0_, Inst_bSbox_AND_M53_U1_n23,
         Inst_bSbox_AND_M53_U1_n22, Inst_bSbox_AND_M53_U1_n21,
         Inst_bSbox_AND_M53_U1_n20, Inst_bSbox_AND_M53_U1_n19,
         Inst_bSbox_AND_M53_U1_n18, Inst_bSbox_AND_M53_U1_n17,
         Inst_bSbox_AND_M53_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M53_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M53_U1_s_out_0__1_, Inst_bSbox_AND_M53_U1_s_out_1__0_,
         Inst_bSbox_AND_M53_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M53_U1_p_0_in_1__0_, Inst_bSbox_AND_M53_U1_s_in_0__1_,
         Inst_bSbox_AND_M53_U1_s_in_1__0_, Inst_bSbox_AND_M54_U1_n23,
         Inst_bSbox_AND_M54_U1_n22, Inst_bSbox_AND_M54_U1_n21,
         Inst_bSbox_AND_M54_U1_n20, Inst_bSbox_AND_M54_U1_n19,
         Inst_bSbox_AND_M54_U1_n18, Inst_bSbox_AND_M54_U1_n17,
         Inst_bSbox_AND_M54_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M54_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M54_U1_s_out_0__1_, Inst_bSbox_AND_M54_U1_s_out_1__0_,
         Inst_bSbox_AND_M54_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M54_U1_p_0_in_1__0_, Inst_bSbox_AND_M54_U1_s_in_0__1_,
         Inst_bSbox_AND_M54_U1_s_in_1__0_, Inst_bSbox_AND_M55_U1_n23,
         Inst_bSbox_AND_M55_U1_n22, Inst_bSbox_AND_M55_U1_n21,
         Inst_bSbox_AND_M55_U1_n20, Inst_bSbox_AND_M55_U1_n19,
         Inst_bSbox_AND_M55_U1_n18, Inst_bSbox_AND_M55_U1_n17,
         Inst_bSbox_AND_M55_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M55_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M55_U1_s_out_0__1_, Inst_bSbox_AND_M55_U1_s_out_1__0_,
         Inst_bSbox_AND_M55_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M55_U1_p_0_in_1__0_, Inst_bSbox_AND_M55_U1_s_in_0__1_,
         Inst_bSbox_AND_M55_U1_s_in_1__0_, Inst_bSbox_AND_M56_U1_n23,
         Inst_bSbox_AND_M56_U1_n22, Inst_bSbox_AND_M56_U1_n21,
         Inst_bSbox_AND_M56_U1_n20, Inst_bSbox_AND_M56_U1_n19,
         Inst_bSbox_AND_M56_U1_n18, Inst_bSbox_AND_M56_U1_n17,
         Inst_bSbox_AND_M56_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M56_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M56_U1_s_out_0__1_, Inst_bSbox_AND_M56_U1_s_out_1__0_,
         Inst_bSbox_AND_M56_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M56_U1_p_0_in_1__0_, Inst_bSbox_AND_M56_U1_s_in_0__1_,
         Inst_bSbox_AND_M56_U1_s_in_1__0_, Inst_bSbox_AND_M57_U1_n23,
         Inst_bSbox_AND_M57_U1_n22, Inst_bSbox_AND_M57_U1_n21,
         Inst_bSbox_AND_M57_U1_n20, Inst_bSbox_AND_M57_U1_n19,
         Inst_bSbox_AND_M57_U1_n18, Inst_bSbox_AND_M57_U1_n17,
         Inst_bSbox_AND_M57_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M57_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M57_U1_s_out_0__1_, Inst_bSbox_AND_M57_U1_s_out_1__0_,
         Inst_bSbox_AND_M57_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M57_U1_p_0_in_1__0_, Inst_bSbox_AND_M57_U1_s_in_0__1_,
         Inst_bSbox_AND_M57_U1_s_in_1__0_, Inst_bSbox_AND_M58_U1_n23,
         Inst_bSbox_AND_M58_U1_n22, Inst_bSbox_AND_M58_U1_n21,
         Inst_bSbox_AND_M58_U1_n20, Inst_bSbox_AND_M58_U1_n19,
         Inst_bSbox_AND_M58_U1_n18, Inst_bSbox_AND_M58_U1_n17,
         Inst_bSbox_AND_M58_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M58_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M58_U1_s_out_0__1_, Inst_bSbox_AND_M58_U1_s_out_1__0_,
         Inst_bSbox_AND_M58_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M58_U1_p_0_in_1__0_, Inst_bSbox_AND_M58_U1_s_in_0__1_,
         Inst_bSbox_AND_M58_U1_s_in_1__0_, Inst_bSbox_AND_M59_U1_n23,
         Inst_bSbox_AND_M59_U1_n22, Inst_bSbox_AND_M59_U1_n21,
         Inst_bSbox_AND_M59_U1_n20, Inst_bSbox_AND_M59_U1_n19,
         Inst_bSbox_AND_M59_U1_n18, Inst_bSbox_AND_M59_U1_n17,
         Inst_bSbox_AND_M59_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M59_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M59_U1_s_out_0__1_, Inst_bSbox_AND_M59_U1_s_out_1__0_,
         Inst_bSbox_AND_M59_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M59_U1_p_0_in_1__0_, Inst_bSbox_AND_M59_U1_s_in_0__1_,
         Inst_bSbox_AND_M59_U1_s_in_1__0_, Inst_bSbox_AND_M60_U1_n23,
         Inst_bSbox_AND_M60_U1_n22, Inst_bSbox_AND_M60_U1_n21,
         Inst_bSbox_AND_M60_U1_n20, Inst_bSbox_AND_M60_U1_n19,
         Inst_bSbox_AND_M60_U1_n18, Inst_bSbox_AND_M60_U1_n17,
         Inst_bSbox_AND_M60_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M60_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M60_U1_s_out_0__1_, Inst_bSbox_AND_M60_U1_s_out_1__0_,
         Inst_bSbox_AND_M60_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M60_U1_p_0_in_1__0_, Inst_bSbox_AND_M60_U1_s_in_0__1_,
         Inst_bSbox_AND_M60_U1_s_in_1__0_, Inst_bSbox_AND_M61_U1_n23,
         Inst_bSbox_AND_M61_U1_n22, Inst_bSbox_AND_M61_U1_n21,
         Inst_bSbox_AND_M61_U1_n20, Inst_bSbox_AND_M61_U1_n19,
         Inst_bSbox_AND_M61_U1_n18, Inst_bSbox_AND_M61_U1_n17,
         Inst_bSbox_AND_M61_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M61_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M61_U1_s_out_0__1_, Inst_bSbox_AND_M61_U1_s_out_1__0_,
         Inst_bSbox_AND_M61_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M61_U1_p_0_in_1__0_, Inst_bSbox_AND_M61_U1_s_in_0__1_,
         Inst_bSbox_AND_M61_U1_s_in_1__0_, Inst_bSbox_AND_M62_U1_n23,
         Inst_bSbox_AND_M62_U1_n22, Inst_bSbox_AND_M62_U1_n21,
         Inst_bSbox_AND_M62_U1_n20, Inst_bSbox_AND_M62_U1_n19,
         Inst_bSbox_AND_M62_U1_n18, Inst_bSbox_AND_M62_U1_n17,
         Inst_bSbox_AND_M62_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M62_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M62_U1_s_out_0__1_, Inst_bSbox_AND_M62_U1_s_out_1__0_,
         Inst_bSbox_AND_M62_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M62_U1_p_0_in_1__0_, Inst_bSbox_AND_M62_U1_s_in_0__1_,
         Inst_bSbox_AND_M62_U1_s_in_1__0_, Inst_bSbox_AND_M63_U1_n23,
         Inst_bSbox_AND_M63_U1_n22, Inst_bSbox_AND_M63_U1_n21,
         Inst_bSbox_AND_M63_U1_n20, Inst_bSbox_AND_M63_U1_n19,
         Inst_bSbox_AND_M63_U1_n18, Inst_bSbox_AND_M63_U1_n17,
         Inst_bSbox_AND_M63_U1_p_0_out_0__1_,
         Inst_bSbox_AND_M63_U1_p_0_out_1__0_,
         Inst_bSbox_AND_M63_U1_s_out_0__1_, Inst_bSbox_AND_M63_U1_s_out_1__0_,
         Inst_bSbox_AND_M63_U1_p_0_in_0__1_,
         Inst_bSbox_AND_M63_U1_p_0_in_1__0_, Inst_bSbox_AND_M63_U1_s_in_0__1_,
         Inst_bSbox_AND_M63_U1_s_in_1__0_;
  wire   [7:0] StateOutXORroundKey;
  wire   [7:0] keyStateIn;
  wire   [7:0] stateArray_inS00ser;
  wire   [7:0] stateArray_inS01ser;
  wire   [7:0] stateArray_inS02ser;
  wire   [7:0] stateArray_inS03ser;
  wire   [7:0] stateArray_inS10ser;
  wire   [7:0] stateArray_inS11ser;
  wire   [7:0] stateArray_inS12ser;
  wire   [7:0] stateArray_inS13ser;
  wire   [7:0] stateArray_inS20ser;
  wire   [7:0] stateArray_inS21ser;
  wire   [7:0] stateArray_inS22ser;
  wire   [7:0] stateArray_inS23ser;
  wire   [7:0] stateArray_inS30ser;
  wire   [7:0] stateArray_inS31ser;
  wire   [7:0] stateArray_inS32ser;
  wire   [7:0] stateArray_outS10ser_MC;
  wire   [31:0] StateInMC;
  wire   [7:0] stateArray_outS20ser_MC;
  wire   [7:0] stateArray_outS30ser_MC;
  wire   [31:0] MCout;
  wire   [7:0] KeyArray_outS01ser_XOR_00;
  wire   [7:0] KeyArray_outS10ser;
  wire   [7:0] KeyArray_inS00ser;
  wire   [7:0] KeyArray_outS11ser;
  wire   [7:0] KeyArray_inS01ser;
  wire   [7:0] KeyArray_outS02ser;
  wire   [7:0] KeyArray_outS12ser;
  wire   [7:0] KeyArray_inS02ser;
  wire   [7:0] KeyArray_outS03ser;
  wire   [7:0] keySBIn;
  wire   [7:0] KeyArray_inS03ser;
  wire   [7:0] KeyArray_outS20ser;
  wire   [7:0] KeyArray_inS10ser;
  wire   [7:0] KeyArray_outS21ser;
  wire   [7:0] KeyArray_inS11ser;
  wire   [7:0] KeyArray_outS22ser;
  wire   [7:0] KeyArray_inS12ser;
  wire   [7:0] KeyArray_outS23ser;
  wire   [7:0] KeyArray_inS13ser;
  wire   [7:0] KeyArray_outS30ser;
  wire   [7:0] KeyArray_inS20ser;
  wire   [7:0] KeyArray_outS31ser;
  wire   [7:0] KeyArray_inS21ser;
  wire   [7:0] KeyArray_outS32ser;
  wire   [7:0] KeyArray_inS22ser;
  wire   [7:0] KeyArray_outS33ser;
  wire   [7:0] KeyArray_inS23ser;
  wire   [7:0] KeyArray_inS31ser;
  wire   [7:0] KeyArray_inS32ser;
  wire   [7:0] KeyArray_inS33ser;
  wire   [7:0] KeyArray_outS01ser_p;
  wire   [7:0] KeyArray_inS30ser;
  wire   [7:0] MixColumns_line0_S13;
  wire   [4:3] MixColumns_line0_S02;
  wire   [4:3] MixColumns_line0_timesTHREE_input2;
  wire   [7:0] MixColumns_line1_S13;
  wire   [4:3] MixColumns_line1_timesTHREE_input2;
  wire   [7:0] MixColumns_line2_S13;
  wire   [4:3] MixColumns_line2_timesTHREE_input2;
  wire   [7:0] MixColumns_line3_S13;
  wire   [7:0] roundConstant;
  wire   [7:0] SboxIn;
  wire   [7:0] StateIn;
  wire   [7:0] SboxOut;
  wire   [7:0] stateArray_inS33ser;
  wire   [7:0] stateArray_input_MC;
  wire   [7:0] KeyArray_inS30par;
  wire   [1:0] Inst_bSbox_AND_M1_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M1_U1_z;
  wire   [1:0] Inst_bSbox_AND_M1_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M2_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M2_U1_z;
  wire   [1:0] Inst_bSbox_AND_M2_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M4_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M4_U1_z;
  wire   [1:0] Inst_bSbox_AND_M4_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M6_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M6_U1_z;
  wire   [1:0] Inst_bSbox_AND_M6_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M7_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M7_U1_z;
  wire   [1:0] Inst_bSbox_AND_M7_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M9_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M9_U1_z;
  wire   [1:0] Inst_bSbox_AND_M9_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M11_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M11_U1_z;
  wire   [1:0] Inst_bSbox_AND_M11_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M12_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M12_U1_z;
  wire   [1:0] Inst_bSbox_AND_M12_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M14_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M14_U1_z;
  wire   [1:0] Inst_bSbox_AND_M14_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M25_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M25_U1_z;
  wire   [1:0] Inst_bSbox_AND_M25_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M31_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M31_U1_z;
  wire   [1:0] Inst_bSbox_AND_M31_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M34_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M34_U1_z;
  wire   [1:0] Inst_bSbox_AND_M34_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M29_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M29_U1_z;
  wire   [1:0] Inst_bSbox_AND_M29_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M30_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M30_U1_z;
  wire   [1:0] Inst_bSbox_AND_M30_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M32_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M32_U1_z;
  wire   [1:0] Inst_bSbox_AND_M32_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M35_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M35_U1_z;
  wire   [1:0] Inst_bSbox_AND_M35_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M46_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M46_U1_z;
  wire   [1:0] Inst_bSbox_AND_M46_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M47_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M47_U1_z;
  wire   [1:0] Inst_bSbox_AND_M47_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M48_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M48_U1_z;
  wire   [1:0] Inst_bSbox_AND_M48_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M49_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M49_U1_z;
  wire   [1:0] Inst_bSbox_AND_M49_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M50_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M50_U1_z;
  wire   [1:0] Inst_bSbox_AND_M50_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M51_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M51_U1_z;
  wire   [1:0] Inst_bSbox_AND_M51_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M52_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M52_U1_z;
  wire   [1:0] Inst_bSbox_AND_M52_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M53_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M53_U1_z;
  wire   [1:0] Inst_bSbox_AND_M53_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M54_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M54_U1_z;
  wire   [1:0] Inst_bSbox_AND_M54_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M55_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M55_U1_z;
  wire   [1:0] Inst_bSbox_AND_M55_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M56_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M56_U1_z;
  wire   [1:0] Inst_bSbox_AND_M56_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M57_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M57_U1_z;
  wire   [1:0] Inst_bSbox_AND_M57_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M58_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M58_U1_z;
  wire   [1:0] Inst_bSbox_AND_M58_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M59_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M59_U1_z;
  wire   [1:0] Inst_bSbox_AND_M59_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M60_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M60_U1_z;
  wire   [1:0] Inst_bSbox_AND_M60_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M61_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M61_U1_z;
  wire   [1:0] Inst_bSbox_AND_M61_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M62_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M62_U1_z;
  wire   [1:0] Inst_bSbox_AND_M62_U1_mul;
  wire   [1:0] Inst_bSbox_AND_M63_U1_a_reg;
  wire   [1:0] Inst_bSbox_AND_M63_U1_z;
  wire   [1:0] Inst_bSbox_AND_M63_U1_mul;

  DFF_X1 ctrl_seq6_SFF_0_Q_reg_FF_FF ( .D(new_AGEMA_signal_4241), .CK(clk),
        .QN(n57) );
  DFF_X1 ctrl_seq6_SFF_1_Q_reg_FF_FF ( .D(new_AGEMA_signal_4245), .CK(clk),
        .QN(n59) );
  DFF_X1 ctrl_seq6_SFF_2_Q_reg_FF_FF ( .D(new_AGEMA_signal_4249), .CK(clk),
        .QN(n56) );
  DFF_X1 ctrl_seq6_SFF_3_Q_reg_FF_FF ( .D(new_AGEMA_signal_4253), .CK(clk),
        .QN(n58) );
  DFF_X1 ctrl_seq6_SFF_4_Q_reg_FF_FF ( .D(new_AGEMA_signal_4257), .CK(clk),
        .QN(n44) );
  DFF_X1 ctrl_seq4_SFF_0_Q_reg_FF_FF ( .D(new_AGEMA_signal_4261), .CK(clk),
        .Q(n281), .QN(n55) );
  DFF_X1 ctrl_seq4_SFF_1_Q_reg_FF_FF ( .D(new_AGEMA_signal_4265), .CK(clk),
        .Q(n66) );
  DFF_X1 ctrl_CSselMC_reg_FF_FF ( .D(new_AGEMA_signal_4269), .CK(clk), .Q(
        ctrl_n6) );
  DFF_X1 ctrl_CSenRC_reg_FF_FF ( .D(new_AGEMA_signal_4273), .CK(clk), .QN(n53)
         );
  DFF_X1 calcRCon_s_current_state_reg_0__FF_FF ( .D(new_AGEMA_signal_6197),
        .CK(clk), .Q(n275), .QN(n52) );
  DFF_X1 calcRCon_s_current_state_reg_1__FF_FF ( .D(new_AGEMA_signal_6201),
        .CK(clk), .Q(n279), .QN(n51) );
  DFF_X1 calcRCon_s_current_state_reg_2__FF_FF ( .D(new_AGEMA_signal_6205),
        .CK(clk), .Q(n272), .QN(n50) );
  DFF_X1 calcRCon_s_current_state_reg_3__FF_FF ( .D(new_AGEMA_signal_6209),
        .CK(clk), .Q(n277), .QN(n49) );
  DFF_X1 calcRCon_s_current_state_reg_4__FF_FF ( .D(new_AGEMA_signal_6213),
        .CK(clk), .Q(n276), .QN(n45) );
  DFF_X1 calcRCon_s_current_state_reg_5__FF_FF ( .D(new_AGEMA_signal_6217),
        .CK(clk), .Q(n274), .QN(n46) );
  DFF_X1 calcRCon_s_current_state_reg_6__FF_FF ( .D(new_AGEMA_signal_6221),
        .CK(clk), .Q(n280), .QN(n48) );
  DFF_X1 calcRCon_s_current_state_reg_7__FF_FF ( .D(new_AGEMA_signal_6225),
        .CK(clk), .Q(n273), .QN(n47) );
  DFF_X1 nReset_reg_FF_FF ( .D(new_AGEMA_signal_6229), .CK(clk), .Q(n14), .QN(
        n278) );
  INV_X4 U157 ( .A(n202), .ZN(n204) );
  INV_X4 U158 ( .A(n239), .ZN(n188) );
  BUF_X1 U159 ( .A(n210), .Z(n190) );
  INV_X1 U160 ( .A(n278), .ZN(n191) );
  INV_X2 U161 ( .A(n278), .ZN(n291) );
  INV_X2 U162 ( .A(n278), .ZN(n296) );
  INV_X2 U163 ( .A(n278), .ZN(n297) );
  INV_X2 U164 ( .A(n278), .ZN(n298) );
  INV_X1 U165 ( .A(n317), .ZN(n192) );
  INV_X4 U166 ( .A(n192), .ZN(n193) );
  INV_X2 U167 ( .A(n237), .ZN(n194) );
  INV_X2 U168 ( .A(n237), .ZN(n195) );
  INV_X2 U169 ( .A(n237), .ZN(n308) );
  INV_X2 U170 ( .A(n237), .ZN(n306) );
  INV_X2 U171 ( .A(n237), .ZN(n307) );
  BUF_X2 U172 ( .A(n278), .Z(n237) );
  INV_X2 U173 ( .A(n192), .ZN(n196) );
  INV_X2 U174 ( .A(n192), .ZN(n197) );
  INV_X2 U175 ( .A(n192), .ZN(n198) );
  INV_X2 U176 ( .A(n192), .ZN(n199) );
  INV_X2 U177 ( .A(n192), .ZN(n200) );
  INV_X2 U178 ( .A(n237), .ZN(n311) );
  INV_X4 U179 ( .A(n237), .ZN(n295) );
  INV_X2 U180 ( .A(n237), .ZN(n310) );
  INV_X2 U181 ( .A(n237), .ZN(n309) );
  BUF_X2 U182 ( .A(new_AGEMA_signal_4009), .Z(n282) );
  BUF_X2 U183 ( .A(new_AGEMA_signal_3833), .Z(n284) );
  BUF_X2 U184 ( .A(new_AGEMA_signal_3765), .Z(n285) );
  BUF_X2 U185 ( .A(new_AGEMA_signal_3629), .Z(n287) );
  BUF_X2 U186 ( .A(n209), .Z(n288) );
  BUF_X4 U187 ( .A(n188), .Z(n290) );
  BUF_X1 U188 ( .A(n204), .Z(n205) );
  BUF_X1 U189 ( .A(n205), .Z(n268) );
  BUF_X1 U190 ( .A(n205), .Z(n269) );
  BUF_X1 U191 ( .A(n205), .Z(n263) );
  BUF_X1 U192 ( .A(n205), .Z(n264) );
  BUF_X1 U193 ( .A(n205), .Z(n271) );
  BUF_X1 U194 ( .A(n204), .Z(n203) );
  BUF_X1 U195 ( .A(n205), .Z(n251) );
  BUF_X1 U196 ( .A(n205), .Z(n252) );
  BUF_X1 U197 ( .A(n205), .Z(n254) );
  BUF_X1 U198 ( .A(n205), .Z(n255) );
  BUF_X1 U199 ( .A(n203), .Z(n253) );
  BUF_X1 U200 ( .A(n204), .Z(n259) );
  BUF_X1 U201 ( .A(n205), .Z(n261) );
  BUF_X1 U202 ( .A(n205), .Z(n257) );
  BUF_X1 U203 ( .A(n203), .Z(n258) );
  BUF_X1 U204 ( .A(n204), .Z(n256) );
  BUF_X1 U205 ( .A(n205), .Z(n267) );
  BUF_X1 U206 ( .A(n205), .Z(n265) );
  BUF_X1 U207 ( .A(n205), .Z(n270) );
  BUF_X1 U208 ( .A(n205), .Z(n262) );
  BUF_X1 U209 ( .A(n205), .Z(n266) );
  INV_X1 U210 ( .A(n203), .ZN(n250) );
  AND4_X1 U211 ( .A1(n57), .A2(n56), .A3(n44), .A4(n59), .ZN(n201) );
  NAND2_X1 U212 ( .A1(n58), .A2(n201), .ZN(n216) );
  NOR2_X4 U213 ( .A1(n237), .A2(n216), .ZN(n202) );
  INV_X2 U214 ( .A(n204), .ZN(n240) );
  INV_X2 U215 ( .A(n204), .ZN(n241) );
  INV_X2 U216 ( .A(n204), .ZN(n242) );
  INV_X2 U217 ( .A(n203), .ZN(n243) );
  INV_X2 U218 ( .A(n204), .ZN(n244) );
  INV_X2 U219 ( .A(n204), .ZN(n245) );
  INV_X2 U220 ( .A(n204), .ZN(n246) );
  INV_X2 U221 ( .A(n204), .ZN(n247) );
  INV_X2 U222 ( .A(n203), .ZN(n248) );
  INV_X2 U223 ( .A(n203), .ZN(n249) );
  INV_X1 U224 ( .A(start), .ZN(n189) );
  INV_X1 U225 ( .A(n237), .ZN(n312) );
  NAND4_X1 U226 ( .A1(n48), .A2(n273), .A3(n277), .A4(n275), .ZN(n207) );
  NAND4_X1 U227 ( .A1(n51), .A2(n45), .A3(n46), .A4(n272), .ZN(n206) );
  NOR2_X1 U228 ( .A1(n207), .A2(n206), .ZN(n208) );
  NOR2_X1 U229 ( .A1(n281), .A2(n66), .ZN(n221) );
  NOR3_X1 U230 ( .A1(n208), .A2(n237), .A3(n221), .ZN(n209) );
  AND2_X4 U231 ( .A1(n14), .A2(ctrl_n6), .ZN(n210) );
  BUF_X1 U232 ( .A(n210), .Z(n318) );
  BUF_X1 U233 ( .A(n210), .Z(n317) );
  BUF_X1 U234 ( .A(n210), .Z(n319) );
  INV_X1 U235 ( .A(n237), .ZN(n292) );
  BUF_X1 U236 ( .A(n210), .Z(n316) );
  BUF_X1 U237 ( .A(n210), .Z(n315) );
  BUF_X1 U238 ( .A(n210), .Z(n321) );
  BUF_X1 U239 ( .A(n210), .Z(n320) );
  INV_X1 U240 ( .A(n237), .ZN(n293) );
  BUF_X1 U241 ( .A(n210), .Z(n313) );
  BUF_X1 U242 ( .A(n210), .Z(n314) );
  INV_X1 U243 ( .A(n278), .ZN(n301) );
  INV_X1 U244 ( .A(n278), .ZN(n300) );
  BUF_X1 U245 ( .A(n210), .Z(n322) );
  NAND4_X1 U246 ( .A1(n272), .A2(n279), .A3(n276), .A4(n274), .ZN(n239) );
  INV_X1 U247 ( .A(n237), .ZN(n294) );
  BUF_X2 U248 ( .A(new_AGEMA_signal_3697), .Z(n286) );
  BUF_X2 U249 ( .A(new_AGEMA_signal_3997), .Z(n283) );
  INV_X2 U250 ( .A(n278), .ZN(n299) );
  INV_X2 U251 ( .A(n278), .ZN(n302) );
  INV_X2 U252 ( .A(n278), .ZN(n303) );
  INV_X2 U253 ( .A(n278), .ZN(n304) );
  INV_X2 U254 ( .A(n278), .ZN(n305) );
  NAND2_X1 U256 ( .A1(n216), .A2(n275), .ZN(n211) );
  NAND2_X1 U257 ( .A1(n273), .A2(n250), .ZN(n224) );
  NAND3_X1 U258 ( .A1(n211), .A2(n224), .A3(n191), .ZN(calcRCon_n51) );
  NAND2_X1 U259 ( .A1(n272), .A2(n216), .ZN(n213) );
  NAND2_X1 U260 ( .A1(n250), .A2(n279), .ZN(n212) );
  NAND3_X1 U261 ( .A1(n213), .A2(n212), .A3(n293), .ZN(calcRCon_n49) );
  NAND2_X1 U262 ( .A1(n216), .A2(n273), .ZN(n215) );
  NAND2_X1 U263 ( .A1(n250), .A2(n280), .ZN(n214) );
  NAND3_X1 U264 ( .A1(n215), .A2(n214), .A3(n312), .ZN(calcRCon_n44) );
  NAND2_X1 U265 ( .A1(n250), .A2(n276), .ZN(n218) );
  NAND2_X1 U266 ( .A1(n216), .A2(n294), .ZN(n236) );
  INV_X1 U267 ( .A(n236), .ZN(n232) );
  NAND2_X1 U268 ( .A1(n232), .A2(n274), .ZN(n217) );
  NAND2_X1 U269 ( .A1(n218), .A2(n217), .ZN(calcRCon_n46) );
  NAND2_X1 U270 ( .A1(n250), .A2(n274), .ZN(n220) );
  NAND2_X1 U271 ( .A1(n232), .A2(n280), .ZN(n219) );
  NAND2_X1 U272 ( .A1(n220), .A2(n219), .ZN(calcRCon_n45) );
  NAND2_X1 U273 ( .A1(n232), .A2(n66), .ZN(ctrl_seq4_SFF_0_QD) );
  INV_X1 U274 ( .A(n221), .ZN(n222) );
  NAND2_X1 U275 ( .A1(n198), .A2(n222), .ZN(n223) );
  NAND2_X1 U276 ( .A1(n253), .A2(n223), .ZN(ctrl_N14) );
  NAND3_X1 U277 ( .A1(n250), .A2(n47), .A3(n272), .ZN(n227) );
  INV_X1 U278 ( .A(n224), .ZN(n231) );
  NAND2_X1 U279 ( .A1(n50), .A2(n231), .ZN(n226) );
  NAND2_X1 U280 ( .A1(n251), .A2(n277), .ZN(n225) );
  NAND4_X1 U281 ( .A1(n292), .A2(n227), .A3(n226), .A4(n225), .ZN(calcRCon_n48) );
  NAND2_X1 U282 ( .A1(n52), .A2(n231), .ZN(n230) );
  NAND3_X1 U283 ( .A1(n47), .A2(n250), .A3(n275), .ZN(n229) );
  NAND2_X1 U284 ( .A1(n232), .A2(n279), .ZN(n228) );
  NAND3_X1 U285 ( .A1(n230), .A2(n229), .A3(n228), .ZN(calcRCon_n50) );
  NAND2_X1 U286 ( .A1(n49), .A2(n231), .ZN(n235) );
  NAND3_X1 U287 ( .A1(n47), .A2(n250), .A3(n277), .ZN(n234) );
  NAND2_X1 U288 ( .A1(n232), .A2(n276), .ZN(n233) );
  NAND3_X1 U289 ( .A1(n235), .A2(n234), .A3(n233), .ZN(calcRCon_n47) );
  NOR2_X1 U290 ( .A1(n55), .A2(n236), .ZN(ctrl_seq4_SFF_1_QD) );
  NOR2_X1 U291 ( .A1(n57), .A2(n237), .ZN(ctrl_seq6_SFF_1_QD) );
  NOR2_X1 U292 ( .A1(n56), .A2(n237), .ZN(ctrl_seq6_SFF_3_QD) );
  NOR2_X1 U293 ( .A1(n47), .A2(n53), .ZN(roundConstant[7]) );
  NOR2_X1 U294 ( .A1(n48), .A2(n53), .ZN(roundConstant[6]) );
  NOR2_X1 U295 ( .A1(n46), .A2(n53), .ZN(roundConstant[5]) );
  NOR2_X1 U296 ( .A1(n45), .A2(n53), .ZN(roundConstant[4]) );
  NOR2_X1 U297 ( .A1(n49), .A2(n53), .ZN(roundConstant[3]) );
  NOR2_X1 U298 ( .A1(n50), .A2(n53), .ZN(roundConstant[2]) );
  NOR2_X1 U299 ( .A1(n51), .A2(n53), .ZN(roundConstant[1]) );
  NOR2_X1 U300 ( .A1(n52), .A2(n53), .ZN(roundConstant[0]) );
  XOR2_X1 U301 ( .A(n57), .B(n44), .Z(n238) );
  NAND2_X1 U302 ( .A1(n292), .A2(n238), .ZN(ctrl_seq6_SFF_0_QD) );
  NAND2_X1 U303 ( .A1(n312), .A2(n59), .ZN(ctrl_seq6_SFF_2_QD) );
  NAND2_X1 U304 ( .A1(n293), .A2(n58), .ZN(ctrl_seq6_SFF_4_QD) );
  NOR4_X1 U305 ( .A1(n55), .A2(n66), .A3(n253), .A4(n239), .ZN(done) );
  XOR2_X1 U29_Ins_0_U1 ( .A(ciphertext_s0[120]), .B(keyStateIn[0]), .Z(
        StateOutXORroundKey[0]) );
  XOR2_X1 U29_Ins_1_U1 ( .A(ciphertext_s1[120]), .B(new_AGEMA_signal_1983),
        .Z(new_AGEMA_signal_1984) );
  XOR2_X1 U30_Ins_0_U1 ( .A(ciphertext_s0[121]), .B(keyStateIn[1]), .Z(
        StateOutXORroundKey[1]) );
  XOR2_X1 U30_Ins_1_U1 ( .A(ciphertext_s1[121]), .B(new_AGEMA_signal_1986),
        .Z(new_AGEMA_signal_1987) );
  XOR2_X1 U31_Ins_0_U1 ( .A(ciphertext_s0[122]), .B(keyStateIn[2]), .Z(
        StateOutXORroundKey[2]) );
  XOR2_X1 U31_Ins_1_U1 ( .A(ciphertext_s1[122]), .B(new_AGEMA_signal_1989),
        .Z(new_AGEMA_signal_1990) );
  XOR2_X1 U32_Ins_0_U1 ( .A(ciphertext_s0[123]), .B(keyStateIn[3]), .Z(
        StateOutXORroundKey[3]) );
  XOR2_X1 U32_Ins_1_U1 ( .A(ciphertext_s1[123]), .B(new_AGEMA_signal_1992),
        .Z(new_AGEMA_signal_1993) );
  XOR2_X1 U33_Ins_0_U1 ( .A(ciphertext_s0[124]), .B(keyStateIn[4]), .Z(
        StateOutXORroundKey[4]) );
  XOR2_X1 U33_Ins_1_U1 ( .A(ciphertext_s1[124]), .B(new_AGEMA_signal_1995),
        .Z(new_AGEMA_signal_1996) );
  XOR2_X1 U34_Ins_0_U1 ( .A(ciphertext_s0[125]), .B(keyStateIn[5]), .Z(
        StateOutXORroundKey[5]) );
  XOR2_X1 U34_Ins_1_U1 ( .A(ciphertext_s1[125]), .B(new_AGEMA_signal_1998),
        .Z(new_AGEMA_signal_1999) );
  XOR2_X1 U35_Ins_0_U1 ( .A(ciphertext_s0[126]), .B(keyStateIn[6]), .Z(
        StateOutXORroundKey[6]) );
  XOR2_X1 U35_Ins_1_U1 ( .A(ciphertext_s1[126]), .B(new_AGEMA_signal_2001),
        .Z(new_AGEMA_signal_2002) );
  XOR2_X1 U36_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(keyStateIn[7]), .Z(
        StateOutXORroundKey[7]) );
  XOR2_X1 U36_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(new_AGEMA_signal_2004),
        .Z(new_AGEMA_signal_2005) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n4), .A2(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n3), .ZN(
        stateArray_S00reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS00ser[0]), .A2(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n2), .ZN(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n3) );
  INV_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n2) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[120]), .A2(n243), .ZN(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n4) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3126) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2156), .A2(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[120]), .A2(n243), .ZN(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S00reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS00ser[1]), .A2(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[121]), .A2(n241), .ZN(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3127) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2159), .A2(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[121]), .A2(n241), .ZN(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S00reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS00ser[2]), .A2(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[122]), .A2(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3128) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2162), .A2(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[122]), .A2(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S00reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS00ser[3]), .A2(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[123]), .A2(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3129) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2165), .A2(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[123]), .A2(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S00reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS00ser[4]), .A2(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[124]), .A2(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3130) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2168), .A2(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[124]), .A2(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S00reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS00ser[5]), .A2(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[125]), .A2(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3131) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2171), .A2(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[125]), .A2(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S00reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS00ser[6]), .A2(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[126]), .A2(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3132) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2174), .A2(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[126]), .A2(n249), .ZN(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S00reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS00ser[7]), .A2(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[127]), .A2(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3133) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2177), .A2(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[127]), .A2(n248), .ZN(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S01reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS01ser[0]), .A2(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[112]), .A2(n248), .ZN(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3134) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2180), .A2(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[112]), .A2(n248), .ZN(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S01reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS01ser[1]), .A2(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[113]), .A2(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3135) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2183), .A2(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[113]), .A2(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S01reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS01ser[2]), .A2(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n247), .ZN(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[114]), .A2(n247), .ZN(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3136) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2186), .A2(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n247), .ZN(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[114]), .A2(n247), .ZN(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S01reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS01ser[3]), .A2(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[115]), .A2(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3137) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2189), .A2(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[115]), .A2(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S01reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS01ser[4]), .A2(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[116]), .A2(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3138) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2192), .A2(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[116]), .A2(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S01reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS01ser[5]), .A2(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n202), .ZN(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[117]), .A2(n202), .ZN(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3139) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2195), .A2(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n202), .ZN(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[117]), .A2(n202), .ZN(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S01reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS01ser[6]), .A2(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[118]), .A2(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3140) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2198), .A2(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[118]), .A2(n246), .ZN(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S01reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS01ser[7]), .A2(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[119]), .A2(n242), .ZN(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3141) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2201), .A2(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[119]), .A2(n242), .ZN(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S02reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS02ser[0]), .A2(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[104]), .A2(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3142) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2204), .A2(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[104]), .A2(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S02reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS02ser[1]), .A2(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[105]), .A2(n240), .ZN(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3143) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2207), .A2(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[105]), .A2(n240), .ZN(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S02reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS02ser[2]), .A2(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[106]), .A2(n243), .ZN(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3144) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2210), .A2(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[106]), .A2(n243), .ZN(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S02reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS02ser[3]), .A2(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[107]), .A2(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3145) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2213), .A2(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[107]), .A2(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S02reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS02ser[4]), .A2(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[108]), .A2(n248), .ZN(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3146) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2216), .A2(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[108]), .A2(n248), .ZN(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S02reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS02ser[5]), .A2(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[109]), .A2(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3147) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2219), .A2(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[109]), .A2(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S02reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS02ser[6]), .A2(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[110]), .A2(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3148) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2222), .A2(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[110]), .A2(n249), .ZN(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S02reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS02ser[7]), .A2(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[111]), .A2(n248), .ZN(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3149) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2225), .A2(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[111]), .A2(n248), .ZN(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S03reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS03ser[0]), .A2(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n249), .ZN(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[96]), .A2(n249), .ZN(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3150) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3046), .A2(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n249), .ZN(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[96]), .A2(n249), .ZN(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S03reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS03ser[1]), .A2(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n249), .ZN(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[97]), .A2(n249), .ZN(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3151) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3048), .A2(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n249), .ZN(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[97]), .A2(n249), .ZN(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S03reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS03ser[2]), .A2(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n247), .ZN(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[98]), .A2(n247), .ZN(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3152) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3050), .A2(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n247), .ZN(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[98]), .A2(n247), .ZN(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S03reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS03ser[3]), .A2(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[99]), .A2(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3153) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3052), .A2(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[99]), .A2(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S03reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS03ser[4]), .A2(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[100]), .A2(n244), .ZN(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3154) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3054), .A2(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[100]), .A2(n244), .ZN(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S03reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS03ser[5]), .A2(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[101]), .A2(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3155) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3056), .A2(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[101]), .A2(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S03reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS03ser[6]), .A2(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[102]), .A2(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3156) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3058), .A2(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[102]), .A2(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S03reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS03ser[7]), .A2(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[103]), .A2(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3157) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3060), .A2(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[103]), .A2(n202), .ZN(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S10reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS10ser[0]), .A2(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[80]), .A2(n240), .ZN(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3158) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2228), .A2(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[80]), .A2(n240), .ZN(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S10reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS10ser[1]), .A2(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n202), .ZN(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[81]), .A2(n202), .ZN(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3159) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2231), .A2(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n202), .ZN(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[81]), .A2(n202), .ZN(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S10reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS10ser[2]), .A2(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[82]), .A2(n245), .ZN(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3160) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2234), .A2(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[82]), .A2(n245), .ZN(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S10reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS10ser[3]), .A2(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[83]), .A2(n245), .ZN(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3161) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2237), .A2(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[83]), .A2(n245), .ZN(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S10reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS10ser[4]), .A2(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[84]), .A2(n244), .ZN(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3162) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2240), .A2(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[84]), .A2(n244), .ZN(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S10reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS10ser[5]), .A2(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n249), .ZN(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[85]), .A2(n249), .ZN(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3163) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2243), .A2(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n249), .ZN(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[85]), .A2(n249), .ZN(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S10reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS10ser[6]), .A2(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n247), .ZN(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[86]), .A2(n247), .ZN(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3164) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2246), .A2(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n247), .ZN(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[86]), .A2(n247), .ZN(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S10reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS10ser[7]), .A2(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[87]), .A2(n246), .ZN(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3165) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2249), .A2(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[87]), .A2(n246), .ZN(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S11reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS11ser[0]), .A2(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[72]), .A2(n246), .ZN(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3166) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2252), .A2(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[72]), .A2(n246), .ZN(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S11reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS11ser[1]), .A2(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[73]), .A2(n246), .ZN(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3167) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2255), .A2(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[73]), .A2(n246), .ZN(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S11reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS11ser[2]), .A2(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[74]), .A2(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3168) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2258), .A2(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[74]), .A2(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S11reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS11ser[3]), .A2(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[75]), .A2(n248), .ZN(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3169) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2261), .A2(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[75]), .A2(n248), .ZN(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S11reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS11ser[4]), .A2(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[76]), .A2(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3170) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2264), .A2(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[76]), .A2(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S11reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS11ser[5]), .A2(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[77]), .A2(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3171) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2267), .A2(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[77]), .A2(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S11reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS11ser[6]), .A2(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[78]), .A2(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3172) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2270), .A2(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[78]), .A2(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S11reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS11ser[7]), .A2(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[79]), .A2(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3173) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2273), .A2(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[79]), .A2(n247), .ZN(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S12reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS12ser[0]), .A2(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[64]), .A2(n246), .ZN(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3174) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2276), .A2(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[64]), .A2(n246), .ZN(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S12reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS12ser[1]), .A2(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n247), .ZN(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[65]), .A2(n247), .ZN(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3175) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2279), .A2(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n247), .ZN(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[65]), .A2(n247), .ZN(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S12reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS12ser[2]), .A2(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[66]), .A2(n241), .ZN(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3176) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2282), .A2(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[66]), .A2(n241), .ZN(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S12reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS12ser[3]), .A2(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[67]), .A2(n243), .ZN(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3177) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2285), .A2(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[67]), .A2(n243), .ZN(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S12reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS12ser[4]), .A2(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[68]), .A2(n240), .ZN(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3178) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2288), .A2(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[68]), .A2(n240), .ZN(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S12reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS12ser[5]), .A2(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n247), .ZN(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[69]), .A2(n247), .ZN(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3179) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2291), .A2(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n247), .ZN(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[69]), .A2(n247), .ZN(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S12reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS12ser[6]), .A2(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[70]), .A2(n241), .ZN(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3180) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2294), .A2(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[70]), .A2(n241), .ZN(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S12reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS12ser[7]), .A2(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[71]), .A2(n245), .ZN(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3181) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2297), .A2(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[71]), .A2(n245), .ZN(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S13reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS13ser[0]), .A2(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n202), .ZN(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[88]), .A2(n202), .ZN(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3182) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3062), .A2(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n202), .ZN(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[88]), .A2(n202), .ZN(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S13reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS13ser[1]), .A2(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[89]), .A2(n242), .ZN(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3183) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3064), .A2(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[89]), .A2(n242), .ZN(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S13reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS13ser[2]), .A2(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[90]), .A2(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3184) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3066), .A2(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[90]), .A2(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S13reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS13ser[3]), .A2(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[91]), .A2(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3185) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3068), .A2(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[91]), .A2(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S13reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS13ser[4]), .A2(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n250), .ZN(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[92]), .A2(n250), .ZN(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3186) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3070), .A2(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n250), .ZN(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[92]), .A2(n250), .ZN(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S13reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS13ser[5]), .A2(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[93]), .A2(n241), .ZN(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3187) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3072), .A2(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[93]), .A2(n241), .ZN(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S13reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS13ser[6]), .A2(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n250), .ZN(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[94]), .A2(n250), .ZN(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3188) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3074), .A2(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n250), .ZN(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[94]), .A2(n250), .ZN(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S13reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS13ser[7]), .A2(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[95]), .A2(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3189) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3076), .A2(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[95]), .A2(n248), .ZN(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S20reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS20ser[0]), .A2(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[40]), .A2(n246), .ZN(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3190) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2300), .A2(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[40]), .A2(n246), .ZN(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S20reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS20ser[1]), .A2(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[41]), .A2(n244), .ZN(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3191) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2303), .A2(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[41]), .A2(n244), .ZN(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S20reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS20ser[2]), .A2(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[42]), .A2(n246), .ZN(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3192) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2306), .A2(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[42]), .A2(n246), .ZN(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S20reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS20ser[3]), .A2(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[43]), .A2(n243), .ZN(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3193) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2309), .A2(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[43]), .A2(n243), .ZN(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S20reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS20ser[4]), .A2(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n202), .ZN(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[44]), .A2(n202), .ZN(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3194) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2312), .A2(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n202), .ZN(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[44]), .A2(n202), .ZN(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S20reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS20ser[5]), .A2(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[45]), .A2(n242), .ZN(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3195) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2315), .A2(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[45]), .A2(n242), .ZN(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S20reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS20ser[6]), .A2(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n248), .ZN(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[46]), .A2(n248), .ZN(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3196) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2318), .A2(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n248), .ZN(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[46]), .A2(n248), .ZN(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S20reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS20ser[7]), .A2(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[47]), .A2(n240), .ZN(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3197) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2321), .A2(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[47]), .A2(n240), .ZN(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S21reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS21ser[0]), .A2(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n246), .ZN(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[32]), .A2(n246), .ZN(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3198) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2324), .A2(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n246), .ZN(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[32]), .A2(n246), .ZN(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S21reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS21ser[1]), .A2(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[33]), .A2(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3199) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2327), .A2(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[33]), .A2(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S21reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS21ser[2]), .A2(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[34]), .A2(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3200) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2330), .A2(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[34]), .A2(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S21reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS21ser[3]), .A2(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[35]), .A2(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3201) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2333), .A2(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[35]), .A2(n243), .ZN(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S21reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS21ser[4]), .A2(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[36]), .A2(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3202) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2336), .A2(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[36]), .A2(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S21reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS21ser[5]), .A2(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[37]), .A2(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3203) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2339), .A2(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[37]), .A2(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S21reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS21ser[6]), .A2(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[38]), .A2(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3204) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2342), .A2(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[38]), .A2(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S21reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS21ser[7]), .A2(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[39]), .A2(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3205) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2345), .A2(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[39]), .A2(n242), .ZN(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S22reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS22ser[0]), .A2(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[56]), .A2(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3206) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2348), .A2(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[56]), .A2(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S22reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS22ser[1]), .A2(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[57]), .A2(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3207) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2351), .A2(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[57]), .A2(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S22reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS22ser[2]), .A2(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[58]), .A2(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3208) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2354), .A2(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[58]), .A2(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S22reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS22ser[3]), .A2(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[59]), .A2(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3209) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2357), .A2(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[59]), .A2(n242), .ZN(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S22reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS22ser[4]), .A2(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[60]), .A2(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3210) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2360), .A2(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[60]), .A2(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S22reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS22ser[5]), .A2(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[61]), .A2(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3211) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2363), .A2(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[61]), .A2(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S22reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS22ser[6]), .A2(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[62]), .A2(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3212) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2366), .A2(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[62]), .A2(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S22reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS22ser[7]), .A2(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[63]), .A2(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3213) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2369), .A2(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[63]), .A2(n241), .ZN(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S23reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS23ser[0]), .A2(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[48]), .A2(n241), .ZN(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3214) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3078), .A2(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[48]), .A2(n241), .ZN(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S23reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS23ser[1]), .A2(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[49]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3215) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3080), .A2(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[49]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S23reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS23ser[2]), .A2(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[50]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3216) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3082), .A2(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[50]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S23reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS23ser[3]), .A2(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[51]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3217) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3084), .A2(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[51]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S23reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS23ser[4]), .A2(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[52]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3218) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3086), .A2(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[52]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S23reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS23ser[5]), .A2(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[53]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3219) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3088), .A2(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[53]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S23reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS23ser[6]), .A2(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[54]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3220) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3090), .A2(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[54]), .A2(n245), .ZN(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S23reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS23ser[7]), .A2(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[55]), .A2(n244), .ZN(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3221) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3092), .A2(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[55]), .A2(n244), .ZN(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S30reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS30ser[0]), .A2(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[0]), .A2(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3222) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2372), .A2(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[0]), .A2(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S30reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS30ser[1]), .A2(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n250), .ZN(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[1]), .A2(n250), .ZN(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3223) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2375), .A2(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n250), .ZN(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[1]), .A2(n250), .ZN(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S30reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS30ser[2]), .A2(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[2]), .A2(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3224) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2378), .A2(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[2]), .A2(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S30reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS30ser[3]), .A2(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[3]), .A2(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3225) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2381), .A2(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[3]), .A2(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S30reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS30ser[4]), .A2(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[4]), .A2(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3226) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2384), .A2(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[4]), .A2(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S30reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS30ser[5]), .A2(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[5]), .A2(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3227) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2387), .A2(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[5]), .A2(n244), .ZN(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S30reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS30ser[6]), .A2(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[6]), .A2(n243), .ZN(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3228) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2390), .A2(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[6]), .A2(n243), .ZN(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S30reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS30ser[7]), .A2(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[7]), .A2(n243), .ZN(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3229) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2393), .A2(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[7]), .A2(n243), .ZN(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S31reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS31ser[0]), .A2(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[24]), .A2(n243), .ZN(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3230) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2396), .A2(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[24]), .A2(n243), .ZN(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S31reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS31ser[1]), .A2(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n243), .ZN(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[25]), .A2(n243), .ZN(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3231) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2399), .A2(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n243), .ZN(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[25]), .A2(n243), .ZN(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S31reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS31ser[2]), .A2(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[26]), .A2(n241), .ZN(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3232) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2402), .A2(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[26]), .A2(n241), .ZN(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S31reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS31ser[3]), .A2(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[27]), .A2(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3233) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2405), .A2(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[27]), .A2(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S31reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS31ser[4]), .A2(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[28]), .A2(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3234) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2408), .A2(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[28]), .A2(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S31reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS31ser[5]), .A2(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[29]), .A2(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3235) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2411), .A2(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[29]), .A2(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S31reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS31ser[6]), .A2(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[30]), .A2(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3236) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2414), .A2(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[30]), .A2(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S31reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS31ser[7]), .A2(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[31]), .A2(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3237) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2417), .A2(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[31]), .A2(n240), .ZN(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S32reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS32ser[0]), .A2(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[16]), .A2(n240), .ZN(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3238) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2420), .A2(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[16]), .A2(n240), .ZN(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S32reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS32ser[1]), .A2(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n240), .ZN(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[17]), .A2(n240), .ZN(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3239) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2423), .A2(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n240), .ZN(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[17]), .A2(n240), .ZN(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S32reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS32ser[2]), .A2(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[18]), .A2(n244), .ZN(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3240) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2426), .A2(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[18]), .A2(n244), .ZN(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S32reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS32ser[3]), .A2(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[19]), .A2(n245), .ZN(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3241) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2429), .A2(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[19]), .A2(n245), .ZN(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S32reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS32ser[4]), .A2(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n241), .ZN(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[20]), .A2(n241), .ZN(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3242) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2432), .A2(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n241), .ZN(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[20]), .A2(n241), .ZN(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S32reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS32ser[5]), .A2(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n202), .ZN(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[21]), .A2(n202), .ZN(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3243) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2435), .A2(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n202), .ZN(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[21]), .A2(n202), .ZN(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S32reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS32ser[6]), .A2(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n244), .ZN(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[22]), .A2(n244), .ZN(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3244) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2438), .A2(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n244), .ZN(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[22]), .A2(n244), .ZN(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S32reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS32ser[7]), .A2(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n245), .ZN(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[23]), .A2(n245), .ZN(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3245) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2441), .A2(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n245), .ZN(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[23]), .A2(n245), .ZN(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS00ser[0]) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[120]), .A2(stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_U2 ( .A(n14), .ZN(
        stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[112]), .A2(n14), .ZN(
        stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2156) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[120]), .A2(stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_U2 ( .A(n14), .ZN(
        stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[112]), .A2(n14), .ZN(
        stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS00ser[1]) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[121]), .A2(stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[113]), .A2(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2159) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[121]), .A2(stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[113]), .A2(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS00ser[2]) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[122]), .A2(stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[114]), .A2(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2162) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[122]), .A2(stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[114]), .A2(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS00ser[3]) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[123]), .A2(stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[115]), .A2(n299), .ZN(
        stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2165) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[123]), .A2(stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[115]), .A2(n299), .ZN(
        stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS00ser[4]) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[124]), .A2(stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[116]), .A2(n304), .ZN(
        stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2168) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[124]), .A2(stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[116]), .A2(n304), .ZN(
        stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS00ser[5]) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[125]), .A2(stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[117]), .A2(n303), .ZN(
        stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2171) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[125]), .A2(stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[117]), .A2(n303), .ZN(
        stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS00ser[6]) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[126]), .A2(stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[118]), .A2(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2174) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[126]), .A2(stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[118]), .A2(n302), .ZN(
        stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS00ser[7]) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[127]), .A2(stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[119]), .A2(n299), .ZN(
        stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2177) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[127]), .A2(stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n6), .ZN(stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[119]), .A2(n299), .ZN(
        stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS01ser[0]) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[112]), .A2(stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[104]), .A2(n303), .ZN(
        stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2180) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[112]), .A2(stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[104]), .A2(n303), .ZN(
        stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS01ser[1]) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[113]), .A2(stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[105]), .A2(n302), .ZN(
        stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2183) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[113]), .A2(stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[105]), .A2(n302), .ZN(
        stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS01ser[2]) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[114]), .A2(stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[106]), .A2(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2186) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[114]), .A2(stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[106]), .A2(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS01ser[3]) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[115]), .A2(stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[107]), .A2(n298), .ZN(
        stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2189) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[115]), .A2(stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[107]), .A2(n298), .ZN(
        stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS01ser[4]) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[116]), .A2(stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[108]), .A2(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2192) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[116]), .A2(stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[108]), .A2(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS01ser[5]) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[117]), .A2(stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[109]), .A2(n296), .ZN(
        stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2195) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[117]), .A2(stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[109]), .A2(n296), .ZN(
        stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS01ser[6]) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[118]), .A2(stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[110]), .A2(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2198) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[118]), .A2(stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[110]), .A2(n304), .ZN(
        stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS01ser[7]) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[119]), .A2(stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[111]), .A2(n299), .ZN(
        stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2201) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[119]), .A2(stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n6), .ZN(stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[111]), .A2(n299), .ZN(
        stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS02ser[0]) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[104]), .A2(stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[96]), .A2(n305), .ZN(
        stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2204) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[104]), .A2(stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[96]), .A2(n305), .ZN(
        stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS02ser[1]) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[105]), .A2(stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[97]), .A2(n303), .ZN(
        stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2207) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[105]), .A2(stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[97]), .A2(n303), .ZN(
        stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS02ser[2]) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[106]), .A2(stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[98]), .A2(n298), .ZN(
        stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2210) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[106]), .A2(stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[98]), .A2(n298), .ZN(
        stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS02ser[3]) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[107]), .A2(stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[99]), .A2(n296), .ZN(
        stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2213) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[107]), .A2(stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[99]), .A2(n296), .ZN(
        stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS02ser[4]) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[108]), .A2(stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[100]), .A2(n304), .ZN(
        stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2216) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[108]), .A2(stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[100]), .A2(n304), .ZN(
        stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS02ser[5]) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[109]), .A2(stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[101]), .A2(n304), .ZN(
        stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2219) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[109]), .A2(stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[101]), .A2(n304), .ZN(
        stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS02ser[6]) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[110]), .A2(stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[102]), .A2(n299), .ZN(
        stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2222) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[110]), .A2(stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[102]), .A2(n299), .ZN(
        stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS02ser[7]) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[111]), .A2(stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[103]), .A2(n298), .ZN(
        stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2225) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[111]), .A2(stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n6), .ZN(stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[103]), .A2(n298), .ZN(
        stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_outS10ser_MC[0]) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[88]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_U1 ( .A1(StateInMC[24]), .A2(n210), .ZN(stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3008) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[88]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2880), .A2(n210), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_outS10ser_MC[1]) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[89]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_U1 ( .A1(StateInMC[25]), .A2(n193), .ZN(stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3009) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[89]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2881), .A2(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_outS10ser_MC[2]) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[90]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_U1 ( .A1(StateInMC[26]), .A2(n210), .ZN(stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3010) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[90]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2882), .A2(n210), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_outS10ser_MC[3]) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[91]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_U1 ( .A1(StateInMC[27]), .A2(n193), .ZN(stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3011) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[91]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2883), .A2(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_outS10ser_MC[4]) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[92]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_U2 ( .A(n321), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_U1 ( .A1(StateInMC[28]), .A2(n321), .ZN(stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3012) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[92]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_U2 ( .A(n321), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2884), .A2(n321), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_outS10ser_MC[5]) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[93]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_U1 ( .A1(StateInMC[29]), .A2(n193), .ZN(stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3013) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[93]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2885), .A2(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_outS10ser_MC[6]) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[94]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_U2 ( .A(n320), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_U1 ( .A1(StateInMC[30]), .A2(n320), .ZN(stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3014) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[94]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_U2 ( .A(n320), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2886), .A2(n320), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_outS10ser_MC[7]) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[95]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_U1 ( .A1(StateInMC[31]), .A2(n193), .ZN(stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3015) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[95]), .A2(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2887), .A2(n193), .ZN(
        stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS03ser[0]) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[96]), .A2(stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        stateArray_outS10ser_MC[0]), .A2(n297), .ZN(
        stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3046) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[96]), .A2(stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3008), .A2(n297), .ZN(
        stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS03ser[1]) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[97]), .A2(stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        stateArray_outS10ser_MC[1]), .A2(n291), .ZN(
        stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3048) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[97]), .A2(stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3009), .A2(n291), .ZN(
        stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS03ser[2]) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[98]), .A2(stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        stateArray_outS10ser_MC[2]), .A2(n304), .ZN(
        stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3050) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[98]), .A2(stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_U2 ( .A(n304), .ZN(
        stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3010), .A2(n304), .ZN(
        stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS03ser[3]) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[99]), .A2(stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        stateArray_outS10ser_MC[3]), .A2(n291), .ZN(
        stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3052) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[99]), .A2(stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3011), .A2(n291), .ZN(
        stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS03ser[4]) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[100]), .A2(stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n6), .ZN(stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        stateArray_outS10ser_MC[4]), .A2(n297), .ZN(
        stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3054) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[100]), .A2(stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n6), .ZN(stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3012), .A2(n297), .ZN(
        stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS03ser[5]) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[101]), .A2(stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n6), .ZN(stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        stateArray_outS10ser_MC[5]), .A2(n305), .ZN(
        stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3056) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[101]), .A2(stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n6), .ZN(stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3013), .A2(n305), .ZN(
        stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS03ser[6]) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[102]), .A2(stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n6), .ZN(stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_U2 ( .A(n301), .ZN(
        stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        stateArray_outS10ser_MC[6]), .A2(n301), .ZN(
        stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3058) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[102]), .A2(stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n6), .ZN(stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_U2 ( .A(n301), .ZN(
        stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3014), .A2(n301), .ZN(
        stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS03ser[7]) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[103]), .A2(stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n6), .ZN(stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_U2 ( .A(n310), .ZN(
        stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        stateArray_outS10ser_MC[7]), .A2(n310), .ZN(
        stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3060) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[103]), .A2(stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n6), .ZN(stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_U2 ( .A(n310), .ZN(
        stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3015), .A2(n310), .ZN(
        stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS10ser[0]) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[88]), .A2(stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[80]), .A2(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2228) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[88]), .A2(stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[80]), .A2(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS10ser[1]) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[89]), .A2(stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_U2 ( .A(n191), .ZN(
        stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[81]), .A2(n191), .ZN(
        stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2231) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[89]), .A2(stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_U2 ( .A(n191), .ZN(
        stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[81]), .A2(n191), .ZN(
        stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS10ser[2]) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[90]), .A2(stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[82]), .A2(n299), .ZN(
        stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2234) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[90]), .A2(stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[82]), .A2(n299), .ZN(
        stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS10ser[3]) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[91]), .A2(stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[83]), .A2(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2237) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[91]), .A2(stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[83]), .A2(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS10ser[4]) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[92]), .A2(stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[84]), .A2(n297), .ZN(
        stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2240) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[92]), .A2(stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[84]), .A2(n297), .ZN(
        stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS10ser[5]) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[93]), .A2(stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[85]), .A2(n298), .ZN(
        stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2243) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[93]), .A2(stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[85]), .A2(n298), .ZN(
        stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS10ser[6]) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[94]), .A2(stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[86]), .A2(n303), .ZN(
        stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2246) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[94]), .A2(stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[86]), .A2(n303), .ZN(
        stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS10ser[7]) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[95]), .A2(stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[87]), .A2(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2249) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[95]), .A2(stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[87]), .A2(n296), .ZN(
        stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS11ser[0]) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[80]), .A2(stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[72]), .A2(n291), .ZN(
        stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2252) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[80]), .A2(stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[72]), .A2(n291), .ZN(
        stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS11ser[1]) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[81]), .A2(stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[73]), .A2(n305), .ZN(
        stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2255) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[81]), .A2(stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[73]), .A2(n305), .ZN(
        stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS11ser[2]) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[82]), .A2(stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[74]), .A2(n302), .ZN(
        stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2258) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[82]), .A2(stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[74]), .A2(n302), .ZN(
        stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS11ser[3]) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[83]), .A2(stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[75]), .A2(n297), .ZN(
        stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2261) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[83]), .A2(stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[75]), .A2(n297), .ZN(
        stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS11ser[4]) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[84]), .A2(stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[76]), .A2(n299), .ZN(
        stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2264) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[84]), .A2(stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[76]), .A2(n299), .ZN(
        stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS11ser[5]) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[85]), .A2(stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[77]), .A2(n298), .ZN(
        stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2267) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[85]), .A2(stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[77]), .A2(n298), .ZN(
        stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS11ser[6]) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[86]), .A2(stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[78]), .A2(n297), .ZN(
        stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2270) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[86]), .A2(stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[78]), .A2(n297), .ZN(
        stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS11ser[7]) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[87]), .A2(stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[79]), .A2(n296), .ZN(
        stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2273) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[87]), .A2(stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[79]), .A2(n296), .ZN(
        stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS12ser[0]) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[72]), .A2(stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[64]), .A2(n303), .ZN(
        stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2276) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[72]), .A2(stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[64]), .A2(n303), .ZN(
        stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS12ser[1]) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[73]), .A2(stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[65]), .A2(n291), .ZN(
        stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2279) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[73]), .A2(stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[65]), .A2(n291), .ZN(
        stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS12ser[2]) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[74]), .A2(stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[66]), .A2(n302), .ZN(
        stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2282) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[74]), .A2(stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[66]), .A2(n302), .ZN(
        stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS12ser[3]) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[75]), .A2(stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[67]), .A2(n296), .ZN(
        stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2285) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[75]), .A2(stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[67]), .A2(n296), .ZN(
        stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS12ser[4]) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[76]), .A2(stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_U2 ( .A(n191), .ZN(
        stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[68]), .A2(n191), .ZN(
        stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2288) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[76]), .A2(stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_U2 ( .A(n191), .ZN(
        stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[68]), .A2(n191), .ZN(
        stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS12ser[5]) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[77]), .A2(stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[69]), .A2(n305), .ZN(
        stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2291) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[77]), .A2(stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[69]), .A2(n305), .ZN(
        stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS12ser[6]) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[78]), .A2(stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_U2 ( .A(n301), .ZN(
        stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[70]), .A2(n301), .ZN(
        stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2294) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[78]), .A2(stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_U2 ( .A(n301), .ZN(
        stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[70]), .A2(n301), .ZN(
        stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS12ser[7]) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[79]), .A2(stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_U2 ( .A(n300), .ZN(
        stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[71]), .A2(n300), .ZN(
        stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2297) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[79]), .A2(stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_U2 ( .A(n300), .ZN(
        stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[71]), .A2(n300), .ZN(
        stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_outS20ser_MC[0]) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[56]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_U1 ( .A1(StateInMC[16]), .A2(n193), .ZN(stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3016) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[56]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2872), .A2(n193), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_outS20ser_MC[1]) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[57]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_U1 ( .A1(StateInMC[17]), .A2(n210), .ZN(stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3017) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[57]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2873), .A2(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_outS20ser_MC[2]) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[58]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_U1 ( .A1(StateInMC[18]), .A2(n210), .ZN(stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3018) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[58]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2874), .A2(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_outS20ser_MC[3]) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[59]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_U1 ( .A1(StateInMC[19]), .A2(n193), .ZN(stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3019) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[59]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2875), .A2(n193), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_outS20ser_MC[4]) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[60]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_U1 ( .A1(StateInMC[20]), .A2(n210), .ZN(stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3020) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[60]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2876), .A2(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_outS20ser_MC[5]) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[61]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_U1 ( .A1(StateInMC[21]), .A2(n193), .ZN(stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3021) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[61]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2877), .A2(n193), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_outS20ser_MC[6]) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[62]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_U2 ( .A(n313), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_U1 ( .A1(StateInMC[22]), .A2(n313), .ZN(stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3022) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[62]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_U2 ( .A(n313), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2878), .A2(n313), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_outS20ser_MC[7]) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[63]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_U1 ( .A1(StateInMC[23]), .A2(n210), .ZN(stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3023) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[63]), .A2(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2879), .A2(n210), .ZN(
        stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS13ser[0]) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[64]), .A2(stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        stateArray_outS20ser_MC[0]), .A2(n291), .ZN(
        stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3062) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[64]), .A2(stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3016), .A2(n291), .ZN(
        stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS13ser[1]) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[65]), .A2(stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        stateArray_outS20ser_MC[1]), .A2(n298), .ZN(
        stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3064) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[65]), .A2(stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3017), .A2(n298), .ZN(
        stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS13ser[2]) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[66]), .A2(stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        stateArray_outS20ser_MC[2]), .A2(n291), .ZN(
        stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3066) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[66]), .A2(stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3018), .A2(n291), .ZN(
        stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS13ser[3]) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[67]), .A2(stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        stateArray_outS20ser_MC[3]), .A2(n305), .ZN(
        stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3068) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[67]), .A2(stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3019), .A2(n305), .ZN(
        stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS13ser[4]) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[68]), .A2(stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        stateArray_outS20ser_MC[4]), .A2(n303), .ZN(
        stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3070) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[68]), .A2(stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3020), .A2(n303), .ZN(
        stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS13ser[5]) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[69]), .A2(stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        stateArray_outS20ser_MC[5]), .A2(n299), .ZN(
        stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3072) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[69]), .A2(stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_U2 ( .A(n299), .ZN(
        stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3021), .A2(n299), .ZN(
        stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS13ser[6]) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[70]), .A2(stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_U2 ( .A(n300), .ZN(
        stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        stateArray_outS20ser_MC[6]), .A2(n300), .ZN(
        stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3074) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[70]), .A2(stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_U2 ( .A(n300), .ZN(
        stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3022), .A2(n300), .ZN(
        stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS13ser[7]) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[71]), .A2(stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        stateArray_outS20ser_MC[7]), .A2(n302), .ZN(
        stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3076) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[71]), .A2(stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_U2 ( .A(n302), .ZN(
        stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3023), .A2(n302), .ZN(
        stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS20ser[0]) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[56]), .A2(stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[48]), .A2(n297), .ZN(
        stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2300) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[56]), .A2(stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[48]), .A2(n297), .ZN(
        stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS20ser[1]) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[57]), .A2(stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[49]), .A2(n296), .ZN(
        stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2303) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[57]), .A2(stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_U2 ( .A(n296), .ZN(
        stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[49]), .A2(n296), .ZN(
        stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS20ser[2]) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[58]), .A2(stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[50]), .A2(n291), .ZN(
        stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2306) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[58]), .A2(stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_U2 ( .A(n291), .ZN(
        stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[50]), .A2(n291), .ZN(
        stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS20ser[3]) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[59]), .A2(stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[51]), .A2(n303), .ZN(
        stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2309) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[59]), .A2(stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_U2 ( .A(n303), .ZN(
        stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[51]), .A2(n303), .ZN(
        stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS20ser[4]) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[60]), .A2(stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[52]), .A2(n305), .ZN(
        stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2312) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[60]), .A2(stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[52]), .A2(n305), .ZN(
        stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS20ser[5]) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[61]), .A2(stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[53]), .A2(n305), .ZN(
        stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2315) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[61]), .A2(stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_U2 ( .A(n305), .ZN(
        stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[53]), .A2(n305), .ZN(
        stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS20ser[6]) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[62]), .A2(stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_U2 ( .A(n195), .ZN(
        stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[54]), .A2(n195), .ZN(
        stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2318) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[62]), .A2(stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_U2 ( .A(n195), .ZN(
        stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[54]), .A2(n195), .ZN(
        stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS20ser[7]) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[63]), .A2(stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_U2 ( .A(n311), .ZN(
        stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[55]), .A2(n311), .ZN(
        stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2321) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[63]), .A2(stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_U2 ( .A(n311), .ZN(
        stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[55]), .A2(n311), .ZN(
        stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS21ser[0]) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[48]), .A2(stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[40]), .A2(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2324) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[48]), .A2(stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[40]), .A2(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS21ser[1]) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[49]), .A2(stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[41]), .A2(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2327) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[49]), .A2(stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[41]), .A2(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS21ser[2]) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[50]), .A2(stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_U2 ( .A(n311), .ZN(
        stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[42]), .A2(n311), .ZN(
        stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2330) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[50]), .A2(stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_U2 ( .A(n311), .ZN(
        stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[42]), .A2(n311), .ZN(
        stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS21ser[3]) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[51]), .A2(stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_U2 ( .A(n306), .ZN(
        stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[43]), .A2(n306), .ZN(
        stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2333) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[51]), .A2(stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_U2 ( .A(n306), .ZN(
        stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[43]), .A2(n306), .ZN(
        stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS21ser[4]) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[52]), .A2(stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_U2 ( .A(n308), .ZN(
        stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[44]), .A2(n308), .ZN(
        stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2336) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[52]), .A2(stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_U2 ( .A(n308), .ZN(
        stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[44]), .A2(n308), .ZN(
        stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS21ser[5]) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[53]), .A2(stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[45]), .A2(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2339) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[53]), .A2(stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[45]), .A2(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS21ser[6]) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[54]), .A2(stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_U2 ( .A(n308), .ZN(
        stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[46]), .A2(n308), .ZN(
        stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2342) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[54]), .A2(stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_U2 ( .A(n308), .ZN(
        stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[46]), .A2(n308), .ZN(
        stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS21ser[7]) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[55]), .A2(stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[47]), .A2(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2345) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[55]), .A2(stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[47]), .A2(n295), .ZN(
        stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS22ser[0]) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[40]), .A2(stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_U2 ( .A(n307), .ZN(
        stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[32]), .A2(n307), .ZN(
        stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2348) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[40]), .A2(stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_U2 ( .A(n307), .ZN(
        stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[32]), .A2(n307), .ZN(
        stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS22ser[1]) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[41]), .A2(stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_U2 ( .A(n309), .ZN(
        stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[33]), .A2(n309), .ZN(
        stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2351) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[41]), .A2(stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_U2 ( .A(n309), .ZN(
        stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[33]), .A2(n309), .ZN(
        stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS22ser[2]) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[42]), .A2(stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[34]), .A2(n295), .ZN(
        stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2354) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[42]), .A2(stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[34]), .A2(n295), .ZN(
        stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS22ser[3]) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[43]), .A2(stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_U2 ( .A(n306), .ZN(
        stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[35]), .A2(n306), .ZN(
        stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2357) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[43]), .A2(stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_U2 ( .A(n306), .ZN(
        stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[35]), .A2(n306), .ZN(
        stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS22ser[4]) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[44]), .A2(stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_U2 ( .A(n308), .ZN(
        stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[36]), .A2(n308), .ZN(
        stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2360) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[44]), .A2(stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_U2 ( .A(n308), .ZN(
        stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[36]), .A2(n308), .ZN(
        stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS22ser[5]) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[45]), .A2(stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_U2 ( .A(n308), .ZN(
        stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[37]), .A2(n308), .ZN(
        stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2363) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[45]), .A2(stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_U2 ( .A(n308), .ZN(
        stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[37]), .A2(n308), .ZN(
        stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS22ser[6]) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[46]), .A2(stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_U2 ( .A(n194), .ZN(
        stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[38]), .A2(n194), .ZN(
        stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2366) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[46]), .A2(stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_U2 ( .A(n194), .ZN(
        stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[38]), .A2(n194), .ZN(
        stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS22ser[7]) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[47]), .A2(stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_U2 ( .A(n294), .ZN(
        stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[39]), .A2(n294), .ZN(
        stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2369) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[47]), .A2(stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_U2 ( .A(n294), .ZN(
        stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[39]), .A2(n294), .ZN(
        stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_outS30ser_MC[0]) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[24]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_U2 ( .A(n313), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_U1 ( .A1(StateInMC[8]),
        .A2(n313), .ZN(stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3024) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[24]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_U2 ( .A(n313), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2864), .A2(n313), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_outS30ser_MC[1]) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[25]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_U1 ( .A1(StateInMC[9]),
        .A2(n210), .ZN(stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3025) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[25]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2865), .A2(n210), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_outS30ser_MC[2]) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[26]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_U1 ( .A1(StateInMC[10]), .A2(n193), .ZN(stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3026) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[26]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2866), .A2(n193), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_outS30ser_MC[3]) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[27]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_U2 ( .A(n320), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_U1 ( .A1(StateInMC[11]), .A2(n320), .ZN(stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3027) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[27]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_U2 ( .A(n320), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2867), .A2(n320), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_outS30ser_MC[4]) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[28]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_U2 ( .A(n322), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_U1 ( .A1(StateInMC[12]), .A2(n322), .ZN(stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3028) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[28]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_U2 ( .A(n322), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2868), .A2(n322), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_outS30ser_MC[5]) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[29]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_U1 ( .A1(StateInMC[13]), .A2(n193), .ZN(stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3029) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[29]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2869), .A2(n193), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_outS30ser_MC[6]) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[30]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_U1 ( .A1(StateInMC[14]), .A2(n210), .ZN(stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3030) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[30]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_U2 ( .A(n210), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2870), .A2(n210), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_outS30ser_MC[7]) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_U3 ( .A1(
        ciphertext_s0[31]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_U1 ( .A1(StateInMC[15]), .A2(n193), .ZN(stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3031) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_U3 ( .A1(
        ciphertext_s1[31]), .A2(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_n6), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_U2 ( .A(n193), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2871), .A2(n193), .ZN(
        stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS23ser[0]) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[32]), .A2(stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_U2 ( .A(n194), .ZN(
        stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        stateArray_outS30ser_MC[0]), .A2(n194), .ZN(
        stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3078) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[32]), .A2(stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_U2 ( .A(n194), .ZN(
        stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3024), .A2(n194), .ZN(
        stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS23ser[1]) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[33]), .A2(stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_U2 ( .A(n310), .ZN(
        stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        stateArray_outS30ser_MC[1]), .A2(n310), .ZN(
        stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3080) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[33]), .A2(stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_U2 ( .A(n310), .ZN(
        stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3025), .A2(n310), .ZN(
        stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS23ser[2]) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[34]), .A2(stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_U2 ( .A(n306), .ZN(
        stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        stateArray_outS30ser_MC[2]), .A2(n306), .ZN(
        stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3082) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[34]), .A2(stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_U2 ( .A(n306), .ZN(
        stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3026), .A2(n306), .ZN(
        stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS23ser[3]) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[35]), .A2(stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_U2 ( .A(n307), .ZN(
        stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        stateArray_outS30ser_MC[3]), .A2(n307), .ZN(
        stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3084) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[35]), .A2(stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_U2 ( .A(n307), .ZN(
        stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3027), .A2(n307), .ZN(
        stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS23ser[4]) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[36]), .A2(stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        stateArray_outS30ser_MC[4]), .A2(n295), .ZN(
        stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3086) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[36]), .A2(stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3028), .A2(n295), .ZN(
        stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS23ser[5]) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[37]), .A2(stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        stateArray_outS30ser_MC[5]), .A2(n298), .ZN(
        stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3088) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[37]), .A2(stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_U2 ( .A(n298), .ZN(
        stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3029), .A2(n298), .ZN(
        stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS23ser[6]) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[38]), .A2(stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        stateArray_outS30ser_MC[6]), .A2(n297), .ZN(
        stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3090) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[38]), .A2(stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_U2 ( .A(n297), .ZN(
        stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3030), .A2(n297), .ZN(
        stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS23ser[7]) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[39]), .A2(stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_U2 ( .A(n310), .ZN(
        stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        stateArray_outS30ser_MC[7]), .A2(n310), .ZN(
        stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3092) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[39]), .A2(stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_U2 ( .A(n310), .ZN(
        stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3031), .A2(n310), .ZN(
        stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS30ser[0]) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[24]), .A2(stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_U2 ( .A(n195), .ZN(
        stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[16]), .A2(n195), .ZN(
        stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2372) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[24]), .A2(stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_U2 ( .A(n195), .ZN(
        stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[16]), .A2(n195), .ZN(
        stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS30ser[1]) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[25]), .A2(stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_U2 ( .A(n310), .ZN(
        stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[17]), .A2(n310), .ZN(
        stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2375) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[25]), .A2(stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_U2 ( .A(n310), .ZN(
        stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[17]), .A2(n310), .ZN(
        stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS30ser[2]) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[26]), .A2(stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_U2 ( .A(n310), .ZN(
        stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[18]), .A2(n310), .ZN(
        stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2378) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[26]), .A2(stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_U2 ( .A(n310), .ZN(
        stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[18]), .A2(n310), .ZN(
        stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS30ser[3]) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[27]), .A2(stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_U2 ( .A(n306), .ZN(
        stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[19]), .A2(n306), .ZN(
        stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2381) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[27]), .A2(stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_U2 ( .A(n306), .ZN(
        stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[19]), .A2(n306), .ZN(
        stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS30ser[4]) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[28]), .A2(stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_U2 ( .A(n309), .ZN(
        stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[20]), .A2(n309), .ZN(
        stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2384) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[28]), .A2(stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_U2 ( .A(n309), .ZN(
        stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[20]), .A2(n309), .ZN(
        stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS30ser[5]) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[29]), .A2(stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[21]), .A2(n295), .ZN(
        stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2387) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[29]), .A2(stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[21]), .A2(n295), .ZN(
        stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS30ser[6]) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[30]), .A2(stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_U2 ( .A(n309), .ZN(
        stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[22]), .A2(n309), .ZN(
        stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2390) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[30]), .A2(stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_U2 ( .A(n309), .ZN(
        stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[22]), .A2(n309), .ZN(
        stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS30ser[7]) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[31]), .A2(stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_U2 ( .A(n307), .ZN(
        stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[23]), .A2(n307), .ZN(
        stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2393) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[31]), .A2(stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_U2 ( .A(n307), .ZN(
        stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[23]), .A2(n307), .ZN(
        stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS31ser[0]) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[16]), .A2(stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_U2 ( .A(n311), .ZN(
        stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[8]), .A2(n311), .ZN(
        stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2396) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[16]), .A2(stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_U2 ( .A(n311), .ZN(
        stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[8]), .A2(n311), .ZN(
        stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS31ser[1]) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[17]), .A2(stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_U2 ( .A(n311), .ZN(
        stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[9]), .A2(n311), .ZN(
        stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2399) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[17]), .A2(stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_U2 ( .A(n311), .ZN(
        stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[9]), .A2(n311), .ZN(
        stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS31ser[2]) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[18]), .A2(stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_U2 ( .A(n307), .ZN(
        stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[10]), .A2(n307), .ZN(
        stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2402) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[18]), .A2(stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_U2 ( .A(n307), .ZN(
        stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[10]), .A2(n307), .ZN(
        stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS31ser[3]) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[19]), .A2(stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_U2 ( .A(n309), .ZN(
        stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[11]), .A2(n309), .ZN(
        stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2405) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[19]), .A2(stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_U2 ( .A(n309), .ZN(
        stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[11]), .A2(n309), .ZN(
        stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS31ser[4]) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[20]), .A2(stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_U2 ( .A(n309), .ZN(
        stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[12]), .A2(n309), .ZN(
        stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2408) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[20]), .A2(stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_U2 ( .A(n309), .ZN(
        stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[12]), .A2(n309), .ZN(
        stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS31ser[5]) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[21]), .A2(stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_U2 ( .A(n195), .ZN(
        stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[13]), .A2(n195), .ZN(
        stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2411) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[21]), .A2(stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_U2 ( .A(n195), .ZN(
        stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[13]), .A2(n195), .ZN(
        stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS31ser[6]) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[22]), .A2(stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_U2 ( .A(n194), .ZN(
        stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[14]), .A2(n194), .ZN(
        stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2414) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[22]), .A2(stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_U2 ( .A(n194), .ZN(
        stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[14]), .A2(n194), .ZN(
        stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS31ser[7]) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[23]), .A2(stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_U2 ( .A(n307), .ZN(
        stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[15]), .A2(n307), .ZN(
        stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2417) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[23]), .A2(stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_U2 ( .A(n307), .ZN(
        stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[15]), .A2(n307), .ZN(
        stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS32ser[0]) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        plaintext_s0[8]), .A2(stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_U2 ( .A(n195), .ZN(
        stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[0]), .A2(n195), .ZN(
        stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2420) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        plaintext_s1[8]), .A2(stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_U2 ( .A(n195), .ZN(
        stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[0]), .A2(n195), .ZN(
        stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS32ser[1]) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        plaintext_s0[9]), .A2(stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_U2 ( .A(n194), .ZN(
        stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[1]), .A2(n194), .ZN(
        stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2423) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        plaintext_s1[9]), .A2(stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_U2 ( .A(n194), .ZN(
        stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[1]), .A2(n194), .ZN(
        stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS32ser[2]) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        plaintext_s0[10]), .A2(stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_U2 ( .A(n311), .ZN(
        stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[2]), .A2(n311), .ZN(
        stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2426) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        plaintext_s1[10]), .A2(stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_U2 ( .A(n311), .ZN(
        stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[2]), .A2(n311), .ZN(
        stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS32ser[3]) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        plaintext_s0[11]), .A2(stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_U2 ( .A(n306), .ZN(
        stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[3]), .A2(n306), .ZN(
        stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2429) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        plaintext_s1[11]), .A2(stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_U2 ( .A(n306), .ZN(
        stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[3]), .A2(n306), .ZN(
        stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS32ser[4]) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        plaintext_s0[12]), .A2(stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[4]), .A2(n295), .ZN(
        stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2432) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        plaintext_s1[12]), .A2(stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_U2 ( .A(n295), .ZN(
        stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[4]), .A2(n295), .ZN(
        stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS32ser[5]) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        plaintext_s0[13]), .A2(stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_U2 ( .A(n195), .ZN(
        stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[5]), .A2(n195), .ZN(
        stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2435) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        plaintext_s1[13]), .A2(stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_U2 ( .A(n195), .ZN(
        stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[5]), .A2(n195), .ZN(
        stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS32ser[6]) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        plaintext_s0[14]), .A2(stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_U2 ( .A(n194), .ZN(
        stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[6]), .A2(n194), .ZN(
        stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2438) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        plaintext_s1[14]), .A2(stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_U2 ( .A(n194), .ZN(
        stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[6]), .A2(n194), .ZN(
        stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS32ser[7]) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        plaintext_s0[15]), .A2(stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_U2 ( .A(n308), .ZN(
        stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        ciphertext_s0[7]), .A2(n308), .ZN(
        stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2441) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        plaintext_s1[15]), .A2(stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n6),
        .ZN(stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_U2 ( .A(n308), .ZN(
        stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        ciphertext_s1[7]), .A2(n308), .ZN(
        stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_0_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_0_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_0_U1_Ins_0_n7), .ZN(StateInMC[0]) );
  NAND2_X1 MUX_StateInMC_mux_inst_0_U1_Ins_0_U3 ( .A1(MCout[0]), .A2(
        MUX_StateInMC_mux_inst_0_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_0_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_0_U1_Ins_0_U1 ( .A1(ciphertext_s0[24]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_0_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_0_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2860) );
  NAND2_X1 MUX_StateInMC_mux_inst_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2825),
        .A2(MUX_StateInMC_mux_inst_0_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_0_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_0_U1_Ins_1_U1 ( .A1(ciphertext_s1[24]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_1_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_1_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_1_U1_Ins_0_n7), .ZN(StateInMC[1]) );
  NAND2_X1 MUX_StateInMC_mux_inst_1_U1_Ins_0_U3 ( .A1(MCout[1]), .A2(
        MUX_StateInMC_mux_inst_1_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_1_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_1_U1_Ins_0_U1 ( .A1(ciphertext_s0[25]), .A2(
        n188), .ZN(MUX_StateInMC_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_1_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_1_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2861) );
  NAND2_X1 MUX_StateInMC_mux_inst_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2849),
        .A2(MUX_StateInMC_mux_inst_1_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_1_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_1_U1_Ins_1_U1 ( .A1(ciphertext_s1[25]), .A2(
        n188), .ZN(MUX_StateInMC_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_2_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_2_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_2_U1_Ins_0_n7), .ZN(StateInMC[2]) );
  NAND2_X1 MUX_StateInMC_mux_inst_2_U1_Ins_0_U3 ( .A1(MCout[2]), .A2(
        MUX_StateInMC_mux_inst_2_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_2_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_2_U1_Ins_0_U1 ( .A1(ciphertext_s0[26]), .A2(
        n188), .ZN(MUX_StateInMC_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_2_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_2_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2834) );
  NAND2_X1 MUX_StateInMC_mux_inst_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2823),
        .A2(MUX_StateInMC_mux_inst_2_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_2_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_2_U1_Ins_1_U1 ( .A1(ciphertext_s1[26]), .A2(
        n188), .ZN(MUX_StateInMC_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_3_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_3_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_3_U1_Ins_0_n7), .ZN(StateInMC[3]) );
  NAND2_X1 MUX_StateInMC_mux_inst_3_U1_Ins_0_U3 ( .A1(MCout[3]), .A2(
        MUX_StateInMC_mux_inst_3_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_3_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_3_U1_Ins_0_U1 ( .A1(ciphertext_s0[27]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_3_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_3_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2862) );
  NAND2_X1 MUX_StateInMC_mux_inst_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2848),
        .A2(MUX_StateInMC_mux_inst_3_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_3_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_3_U1_Ins_1_U1 ( .A1(ciphertext_s1[27]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_4_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_4_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_4_U1_Ins_0_n7), .ZN(StateInMC[4]) );
  NAND2_X1 MUX_StateInMC_mux_inst_4_U1_Ins_0_U3 ( .A1(MCout[4]), .A2(
        MUX_StateInMC_mux_inst_4_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_4_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_4_U1_Ins_0_U1 ( .A1(ciphertext_s0[28]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_4_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_4_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2863) );
  NAND2_X1 MUX_StateInMC_mux_inst_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2847),
        .A2(MUX_StateInMC_mux_inst_4_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_4_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_4_U1_Ins_1_U1 ( .A1(ciphertext_s1[28]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_5_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_5_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_5_U1_Ins_0_n7), .ZN(StateInMC[5]) );
  NAND2_X1 MUX_StateInMC_mux_inst_5_U1_Ins_0_U3 ( .A1(MCout[5]), .A2(
        MUX_StateInMC_mux_inst_5_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_5_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_5_U1_Ins_0_U1 ( .A1(ciphertext_s0[29]), .A2(
        n188), .ZN(MUX_StateInMC_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_5_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_5_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2835) );
  NAND2_X1 MUX_StateInMC_mux_inst_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2820),
        .A2(MUX_StateInMC_mux_inst_5_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_5_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_5_U1_Ins_1_U1 ( .A1(ciphertext_s1[29]), .A2(
        n188), .ZN(MUX_StateInMC_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_6_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_6_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_6_U1_Ins_0_n7), .ZN(StateInMC[6]) );
  NAND2_X1 MUX_StateInMC_mux_inst_6_U1_Ins_0_U3 ( .A1(MCout[6]), .A2(
        MUX_StateInMC_mux_inst_6_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_6_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_6_U1_Ins_0_U1 ( .A1(ciphertext_s0[30]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_6_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_6_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2836) );
  NAND2_X1 MUX_StateInMC_mux_inst_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2819),
        .A2(MUX_StateInMC_mux_inst_6_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_6_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_6_U1_Ins_1_U1 ( .A1(ciphertext_s1[30]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_7_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_7_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_7_U1_Ins_0_n7), .ZN(StateInMC[7]) );
  NAND2_X1 MUX_StateInMC_mux_inst_7_U1_Ins_0_U3 ( .A1(MCout[7]), .A2(
        MUX_StateInMC_mux_inst_7_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_7_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_7_U1_Ins_0_U1 ( .A1(ciphertext_s0[31]), .A2(
        n188), .ZN(MUX_StateInMC_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_7_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_7_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2837) );
  NAND2_X1 MUX_StateInMC_mux_inst_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2818),
        .A2(MUX_StateInMC_mux_inst_7_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_7_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_7_U1_Ins_1_U1 ( .A1(ciphertext_s1[31]), .A2(
        n188), .ZN(MUX_StateInMC_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_8_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_8_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_8_U1_Ins_0_n7), .ZN(StateInMC[8]) );
  NAND2_X1 MUX_StateInMC_mux_inst_8_U1_Ins_0_U3 ( .A1(MCout[8]), .A2(
        MUX_StateInMC_mux_inst_8_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_8_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_8_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_8_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_8_U1_Ins_0_U1 ( .A1(ciphertext_s0[56]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_8_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_8_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_8_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_8_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2864) );
  NAND2_X1 MUX_StateInMC_mux_inst_8_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2817),
        .A2(MUX_StateInMC_mux_inst_8_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_8_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_8_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_8_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_8_U1_Ins_1_U1 ( .A1(ciphertext_s1[56]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_8_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_9_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_9_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_9_U1_Ins_0_n7), .ZN(StateInMC[9]) );
  NAND2_X1 MUX_StateInMC_mux_inst_9_U1_Ins_0_U3 ( .A1(MCout[9]), .A2(
        MUX_StateInMC_mux_inst_9_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_9_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_9_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_9_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_9_U1_Ins_0_U1 ( .A1(ciphertext_s0[57]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_9_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_9_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_9_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_9_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2865) );
  NAND2_X1 MUX_StateInMC_mux_inst_9_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2846),
        .A2(MUX_StateInMC_mux_inst_9_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_9_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_9_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_9_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_9_U1_Ins_1_U1 ( .A1(ciphertext_s1[57]), .A2(
        n290), .ZN(MUX_StateInMC_mux_inst_9_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_10_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_10_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_10_U1_Ins_0_n7), .ZN(StateInMC[10]) );
  NAND2_X1 MUX_StateInMC_mux_inst_10_U1_Ins_0_U3 ( .A1(MCout[10]), .A2(
        MUX_StateInMC_mux_inst_10_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_10_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_10_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_10_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_10_U1_Ins_0_U1 ( .A1(ciphertext_s0[58]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_10_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_10_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_10_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_10_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2866) );
  NAND2_X1 MUX_StateInMC_mux_inst_10_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2815),
        .A2(MUX_StateInMC_mux_inst_10_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_10_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_10_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_10_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_10_U1_Ins_1_U1 ( .A1(ciphertext_s1[58]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_10_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_11_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_11_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_11_U1_Ins_0_n7), .ZN(StateInMC[11]) );
  NAND2_X1 MUX_StateInMC_mux_inst_11_U1_Ins_0_U3 ( .A1(MCout[11]), .A2(
        MUX_StateInMC_mux_inst_11_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_11_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_11_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_11_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_11_U1_Ins_0_U1 ( .A1(ciphertext_s0[59]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_11_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_11_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_11_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_11_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2867) );
  NAND2_X1 MUX_StateInMC_mux_inst_11_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2845),
        .A2(MUX_StateInMC_mux_inst_11_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_11_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_11_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_11_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_11_U1_Ins_1_U1 ( .A1(ciphertext_s1[59]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_11_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_12_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_12_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_12_U1_Ins_0_n7), .ZN(StateInMC[12]) );
  NAND2_X1 MUX_StateInMC_mux_inst_12_U1_Ins_0_U3 ( .A1(MCout[12]), .A2(
        MUX_StateInMC_mux_inst_12_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_12_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_12_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_12_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_12_U1_Ins_0_U1 ( .A1(ciphertext_s0[60]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_12_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_12_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_12_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_12_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2868) );
  NAND2_X1 MUX_StateInMC_mux_inst_12_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2844),
        .A2(MUX_StateInMC_mux_inst_12_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_12_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_12_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_12_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_12_U1_Ins_1_U1 ( .A1(ciphertext_s1[60]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_12_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_13_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_13_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_13_U1_Ins_0_n7), .ZN(StateInMC[13]) );
  NAND2_X1 MUX_StateInMC_mux_inst_13_U1_Ins_0_U3 ( .A1(MCout[13]), .A2(
        MUX_StateInMC_mux_inst_13_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_13_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_13_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_13_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_13_U1_Ins_0_U1 ( .A1(ciphertext_s0[61]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_13_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_13_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_13_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_13_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2869) );
  NAND2_X1 MUX_StateInMC_mux_inst_13_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2812),
        .A2(MUX_StateInMC_mux_inst_13_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_13_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_13_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_13_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_13_U1_Ins_1_U1 ( .A1(ciphertext_s1[61]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_13_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_14_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_14_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_14_U1_Ins_0_n7), .ZN(StateInMC[14]) );
  NAND2_X1 MUX_StateInMC_mux_inst_14_U1_Ins_0_U3 ( .A1(MCout[14]), .A2(
        MUX_StateInMC_mux_inst_14_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_14_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_14_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_14_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_14_U1_Ins_0_U1 ( .A1(ciphertext_s0[62]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_14_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_14_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_14_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_14_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2870) );
  NAND2_X1 MUX_StateInMC_mux_inst_14_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2811),
        .A2(MUX_StateInMC_mux_inst_14_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_14_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_14_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_14_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_14_U1_Ins_1_U1 ( .A1(ciphertext_s1[62]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_14_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_15_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_15_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_15_U1_Ins_0_n7), .ZN(StateInMC[15]) );
  NAND2_X1 MUX_StateInMC_mux_inst_15_U1_Ins_0_U3 ( .A1(MCout[15]), .A2(
        MUX_StateInMC_mux_inst_15_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_15_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_15_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_15_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_15_U1_Ins_0_U1 ( .A1(ciphertext_s0[63]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_15_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_15_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_15_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_15_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2871) );
  NAND2_X1 MUX_StateInMC_mux_inst_15_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2810),
        .A2(MUX_StateInMC_mux_inst_15_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_15_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_15_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_15_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_15_U1_Ins_1_U1 ( .A1(ciphertext_s1[63]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_15_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_16_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_16_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_16_U1_Ins_0_n7), .ZN(StateInMC[16]) );
  NAND2_X1 MUX_StateInMC_mux_inst_16_U1_Ins_0_U3 ( .A1(MCout[16]), .A2(
        MUX_StateInMC_mux_inst_16_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_16_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_16_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_16_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_16_U1_Ins_0_U1 ( .A1(ciphertext_s0[88]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_16_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_16_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_16_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_16_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2872) );
  NAND2_X1 MUX_StateInMC_mux_inst_16_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2809),
        .A2(MUX_StateInMC_mux_inst_16_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_16_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_16_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_16_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_16_U1_Ins_1_U1 ( .A1(ciphertext_s1[88]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_16_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_17_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_17_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_17_U1_Ins_0_n7), .ZN(StateInMC[17]) );
  NAND2_X1 MUX_StateInMC_mux_inst_17_U1_Ins_0_U3 ( .A1(MCout[17]), .A2(
        MUX_StateInMC_mux_inst_17_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_17_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_17_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_17_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_17_U1_Ins_0_U1 ( .A1(ciphertext_s0[89]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_17_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_17_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_17_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_17_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2873) );
  NAND2_X1 MUX_StateInMC_mux_inst_17_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2843),
        .A2(MUX_StateInMC_mux_inst_17_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_17_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_17_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_17_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_17_U1_Ins_1_U1 ( .A1(ciphertext_s1[89]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_17_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_18_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_18_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_18_U1_Ins_0_n7), .ZN(StateInMC[18]) );
  NAND2_X1 MUX_StateInMC_mux_inst_18_U1_Ins_0_U3 ( .A1(MCout[18]), .A2(
        MUX_StateInMC_mux_inst_18_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_18_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_18_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_18_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_18_U1_Ins_0_U1 ( .A1(ciphertext_s0[90]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_18_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_18_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_18_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_18_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2874) );
  NAND2_X1 MUX_StateInMC_mux_inst_18_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2807),
        .A2(MUX_StateInMC_mux_inst_18_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_18_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_18_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_18_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_18_U1_Ins_1_U1 ( .A1(ciphertext_s1[90]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_18_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_19_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_19_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_19_U1_Ins_0_n7), .ZN(StateInMC[19]) );
  NAND2_X1 MUX_StateInMC_mux_inst_19_U1_Ins_0_U3 ( .A1(MCout[19]), .A2(
        MUX_StateInMC_mux_inst_19_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_19_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_19_U1_Ins_0_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_19_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_19_U1_Ins_0_U1 ( .A1(ciphertext_s0[91]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_19_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_19_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_19_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_19_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2875) );
  NAND2_X1 MUX_StateInMC_mux_inst_19_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2842),
        .A2(MUX_StateInMC_mux_inst_19_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_19_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_19_U1_Ins_1_U2 ( .A(n290), .ZN(
        MUX_StateInMC_mux_inst_19_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_19_U1_Ins_1_U1 ( .A1(ciphertext_s1[91]),
        .A2(n290), .ZN(MUX_StateInMC_mux_inst_19_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_20_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_20_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_20_U1_Ins_0_n7), .ZN(StateInMC[20]) );
  NAND2_X1 MUX_StateInMC_mux_inst_20_U1_Ins_0_U3 ( .A1(MCout[20]), .A2(
        MUX_StateInMC_mux_inst_20_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_20_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_20_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_20_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_20_U1_Ins_0_U1 ( .A1(ciphertext_s0[92]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_20_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_20_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_20_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_20_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2876) );
  NAND2_X1 MUX_StateInMC_mux_inst_20_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2841),
        .A2(MUX_StateInMC_mux_inst_20_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_20_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_20_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_20_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_20_U1_Ins_1_U1 ( .A1(ciphertext_s1[92]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_20_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_21_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_21_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_21_U1_Ins_0_n7), .ZN(StateInMC[21]) );
  NAND2_X1 MUX_StateInMC_mux_inst_21_U1_Ins_0_U3 ( .A1(MCout[21]), .A2(
        MUX_StateInMC_mux_inst_21_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_21_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_21_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_21_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_21_U1_Ins_0_U1 ( .A1(ciphertext_s0[93]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_21_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_21_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_21_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_21_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2877) );
  NAND2_X1 MUX_StateInMC_mux_inst_21_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2804),
        .A2(MUX_StateInMC_mux_inst_21_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_21_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_21_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_21_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_21_U1_Ins_1_U1 ( .A1(ciphertext_s1[93]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_21_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_22_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_22_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_22_U1_Ins_0_n7), .ZN(StateInMC[22]) );
  NAND2_X1 MUX_StateInMC_mux_inst_22_U1_Ins_0_U3 ( .A1(MCout[22]), .A2(
        MUX_StateInMC_mux_inst_22_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_22_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_22_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_22_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_22_U1_Ins_0_U1 ( .A1(ciphertext_s0[94]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_22_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_22_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_22_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_22_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2878) );
  NAND2_X1 MUX_StateInMC_mux_inst_22_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2803),
        .A2(MUX_StateInMC_mux_inst_22_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_22_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_22_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_22_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_22_U1_Ins_1_U1 ( .A1(ciphertext_s1[94]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_22_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_23_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_23_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_23_U1_Ins_0_n7), .ZN(StateInMC[23]) );
  NAND2_X1 MUX_StateInMC_mux_inst_23_U1_Ins_0_U3 ( .A1(MCout[23]), .A2(
        MUX_StateInMC_mux_inst_23_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_23_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_23_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_23_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_23_U1_Ins_0_U1 ( .A1(ciphertext_s0[95]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_23_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_23_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_23_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_23_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2879) );
  NAND2_X1 MUX_StateInMC_mux_inst_23_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2802),
        .A2(MUX_StateInMC_mux_inst_23_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_23_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_23_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_23_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_23_U1_Ins_1_U1 ( .A1(ciphertext_s1[95]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_23_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_24_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_24_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_24_U1_Ins_0_n7), .ZN(StateInMC[24]) );
  NAND2_X1 MUX_StateInMC_mux_inst_24_U1_Ins_0_U3 ( .A1(MCout[24]), .A2(
        MUX_StateInMC_mux_inst_24_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_24_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_24_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_24_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_24_U1_Ins_0_U1 ( .A1(ciphertext_s0[120]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_24_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_24_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_24_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_24_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2880) );
  NAND2_X1 MUX_StateInMC_mux_inst_24_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2801),
        .A2(MUX_StateInMC_mux_inst_24_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_24_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_24_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_24_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_24_U1_Ins_1_U1 ( .A1(ciphertext_s1[120]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_24_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_25_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_25_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_25_U1_Ins_0_n7), .ZN(StateInMC[25]) );
  NAND2_X1 MUX_StateInMC_mux_inst_25_U1_Ins_0_U3 ( .A1(MCout[25]), .A2(
        MUX_StateInMC_mux_inst_25_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_25_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_25_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_25_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_25_U1_Ins_0_U1 ( .A1(ciphertext_s0[121]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_25_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_25_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_25_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_25_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2881) );
  NAND2_X1 MUX_StateInMC_mux_inst_25_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2840),
        .A2(MUX_StateInMC_mux_inst_25_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_25_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_25_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_25_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_25_U1_Ins_1_U1 ( .A1(ciphertext_s1[121]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_25_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_26_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_26_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_26_U1_Ins_0_n7), .ZN(StateInMC[26]) );
  NAND2_X1 MUX_StateInMC_mux_inst_26_U1_Ins_0_U3 ( .A1(MCout[26]), .A2(
        MUX_StateInMC_mux_inst_26_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_26_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_26_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_26_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_26_U1_Ins_0_U1 ( .A1(ciphertext_s0[122]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_26_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_26_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_26_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_26_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2882) );
  NAND2_X1 MUX_StateInMC_mux_inst_26_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2799),
        .A2(MUX_StateInMC_mux_inst_26_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_26_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_26_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_26_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_26_U1_Ins_1_U1 ( .A1(ciphertext_s1[122]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_26_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_27_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_27_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_27_U1_Ins_0_n7), .ZN(StateInMC[27]) );
  NAND2_X1 MUX_StateInMC_mux_inst_27_U1_Ins_0_U3 ( .A1(MCout[27]), .A2(
        MUX_StateInMC_mux_inst_27_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_27_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_27_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_27_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_27_U1_Ins_0_U1 ( .A1(ciphertext_s0[123]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_27_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_27_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_27_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_27_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2883) );
  NAND2_X1 MUX_StateInMC_mux_inst_27_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2839),
        .A2(MUX_StateInMC_mux_inst_27_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_27_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_27_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_27_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_27_U1_Ins_1_U1 ( .A1(ciphertext_s1[123]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_27_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_28_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_28_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_28_U1_Ins_0_n7), .ZN(StateInMC[28]) );
  NAND2_X1 MUX_StateInMC_mux_inst_28_U1_Ins_0_U3 ( .A1(MCout[28]), .A2(
        MUX_StateInMC_mux_inst_28_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_28_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_28_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_28_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_28_U1_Ins_0_U1 ( .A1(ciphertext_s0[124]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_28_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_28_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_28_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_28_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2884) );
  NAND2_X1 MUX_StateInMC_mux_inst_28_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2838),
        .A2(MUX_StateInMC_mux_inst_28_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_28_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_28_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_28_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_28_U1_Ins_1_U1 ( .A1(ciphertext_s1[124]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_28_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_29_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_29_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_29_U1_Ins_0_n7), .ZN(StateInMC[29]) );
  NAND2_X1 MUX_StateInMC_mux_inst_29_U1_Ins_0_U3 ( .A1(MCout[29]), .A2(
        MUX_StateInMC_mux_inst_29_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_29_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_29_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_29_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_29_U1_Ins_0_U1 ( .A1(ciphertext_s0[125]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_29_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_29_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_29_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_29_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2885) );
  NAND2_X1 MUX_StateInMC_mux_inst_29_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2796),
        .A2(MUX_StateInMC_mux_inst_29_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_29_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_29_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_29_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_29_U1_Ins_1_U1 ( .A1(ciphertext_s1[125]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_29_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_30_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_30_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_30_U1_Ins_0_n7), .ZN(StateInMC[30]) );
  NAND2_X1 MUX_StateInMC_mux_inst_30_U1_Ins_0_U3 ( .A1(MCout[30]), .A2(
        MUX_StateInMC_mux_inst_30_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_30_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_30_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_30_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_30_U1_Ins_0_U1 ( .A1(ciphertext_s0[126]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_30_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_30_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_30_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_30_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2886) );
  NAND2_X1 MUX_StateInMC_mux_inst_30_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2795),
        .A2(MUX_StateInMC_mux_inst_30_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_30_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_30_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_30_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_30_U1_Ins_1_U1 ( .A1(ciphertext_s1[126]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_30_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_31_U1_Ins_0_U4 ( .A1(
        MUX_StateInMC_mux_inst_31_U1_Ins_0_n8), .A2(
        MUX_StateInMC_mux_inst_31_U1_Ins_0_n7), .ZN(StateInMC[31]) );
  NAND2_X1 MUX_StateInMC_mux_inst_31_U1_Ins_0_U3 ( .A1(MCout[31]), .A2(
        MUX_StateInMC_mux_inst_31_U1_Ins_0_n6), .ZN(
        MUX_StateInMC_mux_inst_31_U1_Ins_0_n7) );
  INV_X1 MUX_StateInMC_mux_inst_31_U1_Ins_0_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_31_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_31_U1_Ins_0_U1 ( .A1(ciphertext_s0[127]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_31_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateInMC_mux_inst_31_U1_Ins_1_U4 ( .A1(
        MUX_StateInMC_mux_inst_31_U1_Ins_1_n8), .A2(
        MUX_StateInMC_mux_inst_31_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2887) );
  NAND2_X1 MUX_StateInMC_mux_inst_31_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2794),
        .A2(MUX_StateInMC_mux_inst_31_U1_Ins_1_n6), .ZN(
        MUX_StateInMC_mux_inst_31_U1_Ins_1_n7) );
  INV_X1 MUX_StateInMC_mux_inst_31_U1_Ins_1_U2 ( .A(n188), .ZN(
        MUX_StateInMC_mux_inst_31_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateInMC_mux_inst_31_U1_Ins_1_U1 ( .A1(ciphertext_s1[127]),
        .A2(n188), .ZN(MUX_StateInMC_mux_inst_31_U1_Ins_1_n8) );
  XOR2_X1 KeyArray_U50_Ins_0_U1 ( .A(KeyArray_outS01ser_7_), .B(keyStateIn[7]),
        .Z(KeyArray_outS01ser_XOR_00[7]) );
  XOR2_X1 KeyArray_U50_Ins_1_U1 ( .A(new_AGEMA_signal_2006), .B(
        new_AGEMA_signal_2004), .Z(new_AGEMA_signal_2007) );
  XOR2_X1 KeyArray_U49_Ins_0_U1 ( .A(KeyArray_outS01ser_6_), .B(keyStateIn[6]),
        .Z(KeyArray_outS01ser_XOR_00[6]) );
  XOR2_X1 KeyArray_U49_Ins_1_U1 ( .A(new_AGEMA_signal_2008), .B(
        new_AGEMA_signal_2001), .Z(new_AGEMA_signal_2009) );
  XOR2_X1 KeyArray_U48_Ins_0_U1 ( .A(KeyArray_outS01ser_5_), .B(keyStateIn[5]),
        .Z(KeyArray_outS01ser_XOR_00[5]) );
  XOR2_X1 KeyArray_U48_Ins_1_U1 ( .A(new_AGEMA_signal_2010), .B(
        new_AGEMA_signal_1998), .Z(new_AGEMA_signal_2011) );
  XOR2_X1 KeyArray_U47_Ins_0_U1 ( .A(KeyArray_outS01ser_4_), .B(keyStateIn[4]),
        .Z(KeyArray_outS01ser_XOR_00[4]) );
  XOR2_X1 KeyArray_U47_Ins_1_U1 ( .A(new_AGEMA_signal_2012), .B(
        new_AGEMA_signal_1995), .Z(new_AGEMA_signal_2013) );
  XOR2_X1 KeyArray_U46_Ins_0_U1 ( .A(KeyArray_outS01ser_3_), .B(keyStateIn[3]),
        .Z(KeyArray_outS01ser_XOR_00[3]) );
  XOR2_X1 KeyArray_U46_Ins_1_U1 ( .A(new_AGEMA_signal_2014), .B(
        new_AGEMA_signal_1992), .Z(new_AGEMA_signal_2015) );
  XOR2_X1 KeyArray_U45_Ins_0_U1 ( .A(KeyArray_outS01ser_2_), .B(keyStateIn[2]),
        .Z(KeyArray_outS01ser_XOR_00[2]) );
  XOR2_X1 KeyArray_U45_Ins_1_U1 ( .A(new_AGEMA_signal_2016), .B(
        new_AGEMA_signal_1989), .Z(new_AGEMA_signal_2017) );
  XOR2_X1 KeyArray_U44_Ins_0_U1 ( .A(KeyArray_outS01ser_1_), .B(keyStateIn[1]),
        .Z(KeyArray_outS01ser_XOR_00[1]) );
  XOR2_X1 KeyArray_U44_Ins_1_U1 ( .A(new_AGEMA_signal_2018), .B(
        new_AGEMA_signal_1986), .Z(new_AGEMA_signal_2019) );
  XOR2_X1 KeyArray_U43_Ins_0_U1 ( .A(KeyArray_outS01ser_0_), .B(keyStateIn[0]),
        .Z(KeyArray_outS01ser_XOR_00[0]) );
  XOR2_X1 KeyArray_U43_Ins_1_U1 ( .A(new_AGEMA_signal_2020), .B(
        new_AGEMA_signal_1983), .Z(new_AGEMA_signal_2021) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_n5) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(keyStateIn[0]), .A2(
        KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n256), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S00reg_gff_1_SFF_0_QD), .A2(n256), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3375)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1983), .A2(KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n256), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3267), .A2(n256), .ZN(KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS00ser[0]), .A2(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n319), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[0]), .A2(n319), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3267) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3247), .A2(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n319), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2491), .A2(n319), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(keyStateIn[1]), .A2(
        KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n259), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S00reg_gff_1_SFF_1_QD), .A2(n259), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3376)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1986), .A2(KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n259), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3268), .A2(n259), .ZN(KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS00ser[1]), .A2(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[1]), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3268) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3249), .A2(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2494), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(keyStateIn[2]), .A2(
        KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n259), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S00reg_gff_1_SFF_2_QD), .A2(n259), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3377)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1989), .A2(KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n259), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3269), .A2(n259), .ZN(KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS00ser[2]), .A2(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[2]), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3269) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3251), .A2(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2497), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(keyStateIn[3]), .A2(
        KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n258), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S00reg_gff_1_SFF_3_QD), .A2(n258), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3378)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1992), .A2(KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n258), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3270), .A2(n258), .ZN(KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS00ser[3]), .A2(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[3]), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3270) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3253), .A2(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2500), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(keyStateIn[4]), .A2(
        KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n265), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S00reg_gff_1_SFF_4_QD), .A2(n265), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3379)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1995), .A2(KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n265), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3271), .A2(n265), .ZN(KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS00ser[4]), .A2(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[4]), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3271) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3255), .A2(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2503), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(keyStateIn[5]), .A2(
        KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n271), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S00reg_gff_1_SFF_5_QD), .A2(n271), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3380)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1998), .A2(KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n271), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3272), .A2(n271), .ZN(KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS00ser[5]), .A2(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[5]), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3272) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3257), .A2(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2506), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(keyStateIn[6]), .A2(
        KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n205), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S00reg_gff_1_SFF_6_QD), .A2(n205), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3381)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2001), .A2(KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n205), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3273), .A2(n205), .ZN(KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS00ser[6]), .A2(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[6]), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3273) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3259), .A2(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2509), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(keyStateIn[7]), .A2(
        KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n253), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S00reg_gff_1_SFF_7_QD), .A2(n253), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3382)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2004), .A2(KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n253), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3274), .A2(n253), .ZN(KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS00ser[7]), .A2(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[7]), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3274) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3261), .A2(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2512), .A2(n210), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS01ser_0_), .A2(KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S01reg_gff_1_SFF_0_QD), .A2(n204), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3275)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2020), .A2(KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2888), .A2(n204), .ZN(KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS01ser[0]), .A2(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n322), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[0]), .A2(n322), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2888) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2444), .A2(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n322), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2515), .A2(n322), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS01ser_1_), .A2(KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n203), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S01reg_gff_1_SFF_1_QD), .A2(n203), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3276)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2018), .A2(KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n203), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2889), .A2(n203), .ZN(KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS01ser[1]), .A2(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n317), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[1]), .A2(n317), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2889) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2447), .A2(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n317), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2518), .A2(n317), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS01ser_2_), .A2(KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n264), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S01reg_gff_1_SFF_2_QD), .A2(n264), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3277)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2016), .A2(KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n264), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2890), .A2(n264), .ZN(KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS01ser[2]), .A2(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n317), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[2]), .A2(n317), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2890) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2450), .A2(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n317), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2521), .A2(n317), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS01ser_3_), .A2(KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n205), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S01reg_gff_1_SFF_3_QD), .A2(n205), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3278)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2014), .A2(KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n205), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2891), .A2(n205), .ZN(KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS01ser[3]), .A2(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[3]), .A2(n198), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2891) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2453), .A2(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2524), .A2(n198), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS01ser_4_), .A2(KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n255), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S01reg_gff_1_SFF_4_QD), .A2(n255), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3279)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2012), .A2(KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n255), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2892), .A2(n255), .ZN(KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS01ser[4]), .A2(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n320), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[4]), .A2(n320), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2892) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2456), .A2(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n320), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2527), .A2(n320), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS01ser_5_), .A2(KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n261), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S01reg_gff_1_SFF_5_QD), .A2(n261), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3280)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2010), .A2(KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n261), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2893), .A2(n261), .ZN(KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS01ser[5]), .A2(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[5]), .A2(n193), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2893) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2459), .A2(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2530), .A2(n193), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS01ser_6_), .A2(KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n261), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S01reg_gff_1_SFF_6_QD), .A2(n261), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3281)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2008), .A2(KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n261), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2894), .A2(n261), .ZN(KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS01ser[6]), .A2(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n322), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[6]), .A2(n322), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2894) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2462), .A2(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n322), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2533), .A2(n322), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS01ser_7_), .A2(KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S01reg_gff_1_SFF_7_QD), .A2(n204), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3282)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2006), .A2(KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2895), .A2(n204), .ZN(KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS01ser[7]), .A2(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[7]), .A2(n193), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2895) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2465), .A2(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2536), .A2(n193), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS02ser[0]), .A2(KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n256), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S02reg_gff_1_SFF_0_QD), .A2(n256), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3283)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2443), .A2(KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n256), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2896), .A2(n256), .ZN(KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS02ser[0]), .A2(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n320), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[0]), .A2(n320), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2896) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2468), .A2(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n320), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2539), .A2(n320), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS02ser[1]), .A2(KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n269), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S02reg_gff_1_SFF_1_QD), .A2(n269), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3284)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2446), .A2(KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n269), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2897), .A2(n269), .ZN(KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS02ser[1]), .A2(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[1]), .A2(n210), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2897) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2471), .A2(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2542), .A2(n210), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS02ser[2]), .A2(KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n269), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S02reg_gff_1_SFF_2_QD), .A2(n269), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3285)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2449), .A2(KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n269), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2898), .A2(n269), .ZN(KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS02ser[2]), .A2(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[2]), .A2(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2898) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2474), .A2(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2545), .A2(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS02ser[3]), .A2(KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n203), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S02reg_gff_1_SFF_3_QD), .A2(n203), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3286)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2452), .A2(KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n203), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2899), .A2(n203), .ZN(KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS02ser[3]), .A2(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n313), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[3]), .A2(n313), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2899) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2477), .A2(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n313), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2548), .A2(n313), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS02ser[4]), .A2(KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n268), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S02reg_gff_1_SFF_4_QD), .A2(n268), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3287)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2455), .A2(KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n268), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2900), .A2(n268), .ZN(KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS02ser[4]), .A2(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n318), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[4]), .A2(n318), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2900) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2480), .A2(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n318), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2551), .A2(n318), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS02ser[5]), .A2(KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n265), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S02reg_gff_1_SFF_5_QD), .A2(n265), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3288)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2458), .A2(KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n265), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2901), .A2(n265), .ZN(KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS02ser[5]), .A2(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n314), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[5]), .A2(n314), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2901) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2483), .A2(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n314), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2554), .A2(n314), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS02ser[6]), .A2(KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n267), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S02reg_gff_1_SFF_6_QD), .A2(n267), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3289)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2461), .A2(KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n267), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2902), .A2(n267), .ZN(KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS02ser[6]), .A2(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[6]), .A2(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2902) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2486), .A2(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2557), .A2(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS02ser[7]), .A2(KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n267), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S02reg_gff_1_SFF_7_QD), .A2(n267), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3290)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2464), .A2(KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n267), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2903), .A2(n267), .ZN(KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS02ser[7]), .A2(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[7]), .A2(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2903) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2489), .A2(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2560), .A2(n316), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS03ser[0]), .A2(KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n271), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S03reg_gff_1_SFF_0_QD), .A2(n271), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3291)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2467), .A2(KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n271), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2904), .A2(n271), .ZN(KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS03ser[0]), .A2(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n315), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(keySBIn[0]),
        .A2(n315), .ZN(KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2904) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2492), .A2(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n315), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2563), .A2(n315), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS03ser[1]), .A2(KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n271), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S03reg_gff_1_SFF_1_QD), .A2(n271), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3292)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2470), .A2(KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n271), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2905), .A2(n271), .ZN(KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS03ser[1]), .A2(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n317), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(keySBIn[1]),
        .A2(n317), .ZN(KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2905) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2495), .A2(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n317), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2566), .A2(n317), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS03ser[2]), .A2(KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n257), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S03reg_gff_1_SFF_2_QD), .A2(n257), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3293)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2473), .A2(KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n257), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2906), .A2(n257), .ZN(KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS03ser[2]), .A2(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(keySBIn[2]),
        .A2(n193), .ZN(KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2906) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2498), .A2(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2569), .A2(n193), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS03ser[3]), .A2(KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n258), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S03reg_gff_1_SFF_3_QD), .A2(n258), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3294)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2476), .A2(KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n258), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2907), .A2(n258), .ZN(KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS03ser[3]), .A2(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n319), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(keySBIn[3]),
        .A2(n319), .ZN(KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2907) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2501), .A2(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n319), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2572), .A2(n319), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS03ser[4]), .A2(KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n258), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S03reg_gff_1_SFF_4_QD), .A2(n258), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3295)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2479), .A2(KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n258), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2908), .A2(n258), .ZN(KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS03ser[4]), .A2(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n315), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(keySBIn[4]),
        .A2(n315), .ZN(KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2908) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2504), .A2(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n315), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2575), .A2(n315), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_n5) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS03ser[5]), .A2(KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n263), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S03reg_gff_1_SFF_5_QD), .A2(n263), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3296)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2482), .A2(KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n263), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2909), .A2(n263), .ZN(KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS03ser[5]), .A2(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n190), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(keySBIn[5]),
        .A2(n190), .ZN(KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2909) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2507), .A2(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n190), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2578), .A2(n190), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_n5) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS03ser[6]), .A2(KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n257), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S03reg_gff_1_SFF_6_QD), .A2(n257), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3297)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2485), .A2(KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n257), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2910), .A2(n257), .ZN(KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS03ser[6]), .A2(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n317), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(keySBIn[6]),
        .A2(n317), .ZN(KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2910) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2510), .A2(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n317), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2581), .A2(n317), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_n5) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS03ser[7]), .A2(KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n271), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S03reg_gff_1_SFF_7_QD), .A2(n271), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3298)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2488), .A2(KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n271), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2911), .A2(n271), .ZN(KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS03ser[7]), .A2(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n319), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(keySBIn[7]),
        .A2(n319), .ZN(KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2911) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2513), .A2(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n319), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2584), .A2(n319), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_n5) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS10ser[0]), .A2(KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n270), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S10reg_gff_1_SFF_0_QD), .A2(n270), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3299)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2491), .A2(KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n270), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2912), .A2(n270), .ZN(KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS10ser[0]), .A2(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[0]), .A2(n193), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2912) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2516), .A2(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2587), .A2(n193), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_n5) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS10ser[1]), .A2(KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n251), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S10reg_gff_1_SFF_1_QD), .A2(n251), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3300)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2494), .A2(KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n251), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2913), .A2(n251), .ZN(KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS10ser[1]), .A2(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n320), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[1]), .A2(n320), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2913) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2519), .A2(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n320), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2590), .A2(n320), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_n5) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS10ser[2]), .A2(KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n251), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S10reg_gff_1_SFF_2_QD), .A2(n251), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3301)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2497), .A2(KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n251), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2914), .A2(n251), .ZN(KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS10ser[2]), .A2(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[2]), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2914) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2522), .A2(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2593), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_n5) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS10ser[3]), .A2(KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S10reg_gff_1_SFF_3_QD), .A2(n204), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3302)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2500), .A2(KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2915), .A2(n204), .ZN(KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS10ser[3]), .A2(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[3]), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2915) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2525), .A2(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2596), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_n5) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS10ser[4]), .A2(KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n269), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S10reg_gff_1_SFF_4_QD), .A2(n269), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3303)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2503), .A2(KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n269), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2916), .A2(n269), .ZN(KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS10ser[4]), .A2(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[4]), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2916) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2528), .A2(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2599), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_n5) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS10ser[5]), .A2(KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n256), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S10reg_gff_1_SFF_5_QD), .A2(n256), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3304)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2506), .A2(KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n256), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2917), .A2(n256), .ZN(KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS10ser[5]), .A2(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[5]), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2917) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2531), .A2(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2602), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_n5) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS10ser[6]), .A2(KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n256), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S10reg_gff_1_SFF_6_QD), .A2(n256), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3305)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2509), .A2(KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n256), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2918), .A2(n256), .ZN(KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS10ser[6]), .A2(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[6]), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2918) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2534), .A2(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2605), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_n5) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS10ser[7]), .A2(KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n269), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S10reg_gff_1_SFF_7_QD), .A2(n269), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3306)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2512), .A2(KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n269), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2919), .A2(n269), .ZN(KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS10ser[7]), .A2(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[7]), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2919) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2537), .A2(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2608), .A2(n198), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS11ser[0]), .A2(KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n267), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S11reg_gff_1_SFF_0_QD), .A2(n267), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3307)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2515), .A2(KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n267), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2920), .A2(n267), .ZN(KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS11ser[0]), .A2(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[0]), .A2(n198), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2920) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2540), .A2(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2611), .A2(n198), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS11ser[1]), .A2(KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n267), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S11reg_gff_1_SFF_1_QD), .A2(n267), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3308)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2518), .A2(KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n267), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2921), .A2(n267), .ZN(KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS11ser[1]), .A2(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[1]), .A2(n198), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2921) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2543), .A2(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2614), .A2(n198), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS11ser[2]), .A2(KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n267), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S11reg_gff_1_SFF_2_QD), .A2(n267), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3309)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2521), .A2(KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n267), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2922), .A2(n267), .ZN(KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS11ser[2]), .A2(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[2]), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2922) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2546), .A2(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2617), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS11ser[3]), .A2(KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n251), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S11reg_gff_1_SFF_3_QD), .A2(n251), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3310)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2524), .A2(KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n251), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2923), .A2(n251), .ZN(KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS11ser[3]), .A2(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[3]), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2923) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2549), .A2(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2620), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS11ser[4]), .A2(KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n252), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S11reg_gff_1_SFF_4_QD), .A2(n252), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3311)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2527), .A2(KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n252), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2924), .A2(n252), .ZN(KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS11ser[4]), .A2(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[4]), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2924) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2552), .A2(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2623), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS11ser[5]), .A2(KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n259), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S11reg_gff_1_SFF_5_QD), .A2(n259), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3312)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2530), .A2(KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n259), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2925), .A2(n259), .ZN(KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS11ser[5]), .A2(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[5]), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2925) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2555), .A2(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2626), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS11ser[6]), .A2(KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n261), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S11reg_gff_1_SFF_6_QD), .A2(n261), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3313)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2533), .A2(KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n261), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2926), .A2(n261), .ZN(KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS11ser[6]), .A2(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[6]), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2926) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2558), .A2(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2629), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS11ser[7]), .A2(KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n257), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S11reg_gff_1_SFF_7_QD), .A2(n257), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3314)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2536), .A2(KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n257), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2927), .A2(n257), .ZN(KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS11ser[7]), .A2(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[7]), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2927) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2561), .A2(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2632), .A2(n197), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS12ser[0]), .A2(KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n203), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S12reg_gff_1_SFF_0_QD), .A2(n203), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3093)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2539), .A2(KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n203), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2928), .A2(n203), .ZN(KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS12ser[0]), .A2(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[0]), .A2(n197), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2928) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2564), .A2(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2635), .A2(n197), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS12ser[1]), .A2(KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n254), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S12reg_gff_1_SFF_1_QD), .A2(n254), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3094)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2542), .A2(KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n254), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2929), .A2(n254), .ZN(KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS12ser[1]), .A2(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[1]), .A2(n197), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2929) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2567), .A2(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2638), .A2(n197), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS12ser[2]), .A2(KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n262), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S12reg_gff_1_SFF_2_QD), .A2(n262), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3095)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2545), .A2(KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n262), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2930), .A2(n262), .ZN(KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS12ser[2]), .A2(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n315), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[2]), .A2(n315), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2930) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2570), .A2(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n315), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2641), .A2(n315), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS12ser[3]), .A2(KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S12reg_gff_1_SFF_3_QD), .A2(n204), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3096)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2548), .A2(KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2931), .A2(n204), .ZN(KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS12ser[3]), .A2(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n321), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[3]), .A2(n321), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2931) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2573), .A2(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n321), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2644), .A2(n321), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS12ser[4]), .A2(KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S12reg_gff_1_SFF_4_QD), .A2(n204), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3097)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2551), .A2(KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2932), .A2(n204), .ZN(KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS12ser[4]), .A2(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n322), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[4]), .A2(n322), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2932) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2576), .A2(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n322), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2647), .A2(n322), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS12ser[5]), .A2(KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n265), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S12reg_gff_1_SFF_5_QD), .A2(n265), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3098)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2554), .A2(KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n265), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2933), .A2(n265), .ZN(KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS12ser[5]), .A2(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n190), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[5]), .A2(n190), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2933) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2579), .A2(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n190), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2650), .A2(n190), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS12ser[6]), .A2(KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n265), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S12reg_gff_1_SFF_6_QD), .A2(n265), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3099)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2557), .A2(KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n265), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2934), .A2(n265), .ZN(KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS12ser[6]), .A2(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[6]), .A2(n193), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2934) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2582), .A2(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2653), .A2(n193), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS12ser[7]), .A2(KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n264), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S12reg_gff_1_SFF_7_QD), .A2(n264), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3100)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2560), .A2(KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n264), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2935), .A2(n264), .ZN(KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS12ser[7]), .A2(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[7]), .A2(n193), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2935) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2585), .A2(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2656), .A2(n193), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(keySBIn[0]), .A2(
        KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n262), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S13reg_gff_1_SFF_0_QD), .A2(n262), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3101)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2563), .A2(KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n262), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2936), .A2(n262), .ZN(KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS13ser[0]), .A2(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[0]), .A2(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2936) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2588), .A2(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2659), .A2(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(keySBIn[1]), .A2(
        KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n255), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S13reg_gff_1_SFF_1_QD), .A2(n255), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3102)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2566), .A2(KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n255), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2937), .A2(n255), .ZN(KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS13ser[1]), .A2(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n318), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[1]), .A2(n318), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2937) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2591), .A2(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n318), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2662), .A2(n318), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(keySBIn[2]), .A2(
        KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S13reg_gff_1_SFF_2_QD), .A2(n204), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3103)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2569), .A2(KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2938), .A2(n204), .ZN(KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS13ser[2]), .A2(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n322), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[2]), .A2(n322), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2938) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2594), .A2(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n322), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2665), .A2(n322), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(keySBIn[3]), .A2(
        KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n271), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S13reg_gff_1_SFF_3_QD), .A2(n271), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3104)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2572), .A2(KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n271), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2939), .A2(n271), .ZN(KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS13ser[3]), .A2(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[3]), .A2(n198), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2939) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2597), .A2(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2668), .A2(n198), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(keySBIn[4]), .A2(
        KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n203), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S13reg_gff_1_SFF_4_QD), .A2(n203), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3105)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2575), .A2(KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n203), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2940), .A2(n203), .ZN(KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS13ser[4]), .A2(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[4]), .A2(n197), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2940) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2600), .A2(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2671), .A2(n197), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_n5) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(keySBIn[5]), .A2(
        KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n270), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S13reg_gff_1_SFF_5_QD), .A2(n270), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3106)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2578), .A2(KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n270), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2941), .A2(n270), .ZN(KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS13ser[5]), .A2(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[5]), .A2(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2941) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2603), .A2(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2674), .A2(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_n5) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(keySBIn[6]), .A2(
        KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n270), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S13reg_gff_1_SFF_6_QD), .A2(n270), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3107)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2581), .A2(KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n270), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2942), .A2(n270), .ZN(KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS13ser[6]), .A2(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[6]), .A2(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2942) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2606), .A2(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2677), .A2(n193), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_n5) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(keySBIn[7]), .A2(
        KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S13reg_gff_1_SFF_7_QD), .A2(n204), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3108)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2584), .A2(KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2943), .A2(n204), .ZN(KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS13ser[7]), .A2(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[7]), .A2(n199), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2943) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2609), .A2(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2680), .A2(n199), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_n5) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS20ser[0]), .A2(KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n254), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S20reg_gff_1_SFF_0_QD), .A2(n254), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3315)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2587), .A2(KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n254), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2944), .A2(n254), .ZN(KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS20ser[0]), .A2(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[0]), .A2(n210), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2944) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2612), .A2(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2683), .A2(n210), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_n5) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS20ser[1]), .A2(KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n253), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S20reg_gff_1_SFF_1_QD), .A2(n253), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3316)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2590), .A2(KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n253), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2945), .A2(n253), .ZN(KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS20ser[1]), .A2(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n313), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[1]), .A2(n313), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2945) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2615), .A2(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n313), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2686), .A2(n313), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_n5) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS20ser[2]), .A2(KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n253), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S20reg_gff_1_SFF_2_QD), .A2(n253), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3317)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2593), .A2(KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n253), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2946), .A2(n253), .ZN(KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS20ser[2]), .A2(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n321), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[2]), .A2(n321), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2946) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2618), .A2(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n321), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2689), .A2(n321), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_n5) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS20ser[3]), .A2(KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n268), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S20reg_gff_1_SFF_3_QD), .A2(n268), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3318)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2596), .A2(KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n268), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2947), .A2(n268), .ZN(KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS20ser[3]), .A2(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[3]), .A2(n199), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2947) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2621), .A2(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2692), .A2(n199), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_n5) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS20ser[4]), .A2(KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n268), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S20reg_gff_1_SFF_4_QD), .A2(n268), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3319)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2599), .A2(KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n268), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2948), .A2(n268), .ZN(KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS20ser[4]), .A2(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[4]), .A2(n200), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2948) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2624), .A2(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2695), .A2(n200), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_n5) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS20ser[5]), .A2(KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n263), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S20reg_gff_1_SFF_5_QD), .A2(n263), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3320)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2602), .A2(KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n263), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2949), .A2(n263), .ZN(KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS20ser[5]), .A2(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n314), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[5]), .A2(n314), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2949) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2627), .A2(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n314), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2698), .A2(n314), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_n5) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS20ser[6]), .A2(KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n262), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S20reg_gff_1_SFF_6_QD), .A2(n262), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3321)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2605), .A2(KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n262), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2950), .A2(n262), .ZN(KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS20ser[6]), .A2(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n316), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[6]), .A2(n316), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2950) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2630), .A2(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n316), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2701), .A2(n316), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_n5) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS20ser[7]), .A2(KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n205), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S20reg_gff_1_SFF_7_QD), .A2(n205), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3322)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2608), .A2(KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n205), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2951), .A2(n205), .ZN(KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS20ser[7]), .A2(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[7]), .A2(n200), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2951) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2633), .A2(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2704), .A2(n200), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS21ser[0]), .A2(KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n251), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S21reg_gff_1_SFF_0_QD), .A2(n251), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3323)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2611), .A2(KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n251), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2952), .A2(n251), .ZN(KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS21ser[0]), .A2(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n313), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[0]), .A2(n313), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2952) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2636), .A2(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n313), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2707), .A2(n313), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS21ser[1]), .A2(KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n255), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S21reg_gff_1_SFF_1_QD), .A2(n255), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3324)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2614), .A2(KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n255), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2953), .A2(n255), .ZN(KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS21ser[1]), .A2(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[1]), .A2(n196), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2953) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2639), .A2(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2710), .A2(n196), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS21ser[2]), .A2(KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n259), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S21reg_gff_1_SFF_2_QD), .A2(n259), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3325)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2617), .A2(KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n259), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2954), .A2(n259), .ZN(KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS21ser[2]), .A2(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[2]), .A2(n210), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2954) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2642), .A2(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2713), .A2(n210), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS21ser[3]), .A2(KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n254), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S21reg_gff_1_SFF_3_QD), .A2(n254), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3326)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2620), .A2(KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n254), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2955), .A2(n254), .ZN(KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS21ser[3]), .A2(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[3]), .A2(n199), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2955) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2645), .A2(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2716), .A2(n199), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS21ser[4]), .A2(KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n270), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S21reg_gff_1_SFF_4_QD), .A2(n270), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3327)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2623), .A2(KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n270), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2956), .A2(n270), .ZN(KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS21ser[4]), .A2(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[4]), .A2(n200), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2956) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2648), .A2(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2719), .A2(n200), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS21ser[5]), .A2(KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n262), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S21reg_gff_1_SFF_5_QD), .A2(n262), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3328)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2626), .A2(KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n262), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2957), .A2(n262), .ZN(KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS21ser[5]), .A2(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n321), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[5]), .A2(n321), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2957) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2651), .A2(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n321), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2722), .A2(n321), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS21ser[6]), .A2(KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n255), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S21reg_gff_1_SFF_6_QD), .A2(n255), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3329)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2629), .A2(KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n255), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2958), .A2(n255), .ZN(KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS21ser[6]), .A2(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[6]), .A2(n196), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2958) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2654), .A2(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2725), .A2(n196), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS21ser[7]), .A2(KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S21reg_gff_1_SFF_7_QD), .A2(n204), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3330)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2632), .A2(KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2959), .A2(n204), .ZN(KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS21ser[7]), .A2(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[7]), .A2(n210), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2959) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2657), .A2(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2728), .A2(n210), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS22ser[0]), .A2(KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n270), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S22reg_gff_1_SFF_0_QD), .A2(n270), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3331)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2635), .A2(KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n270), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2960), .A2(n270), .ZN(KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS22ser[0]), .A2(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[0]), .A2(n193), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2960) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2660), .A2(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2731), .A2(n193), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS22ser[1]), .A2(KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n252), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S22reg_gff_1_SFF_1_QD), .A2(n252), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3332)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2638), .A2(KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n252), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2961), .A2(n252), .ZN(KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS22ser[1]), .A2(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n190), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[1]), .A2(n190), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2961) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2663), .A2(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n190), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2734), .A2(n190), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS22ser[2]), .A2(KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n266), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S22reg_gff_1_SFF_2_QD), .A2(n266), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3333)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2641), .A2(KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n266), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2962), .A2(n266), .ZN(KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS22ser[2]), .A2(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[2]), .A2(n196), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2962) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2666), .A2(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2737), .A2(n196), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS22ser[3]), .A2(KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n253), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S22reg_gff_1_SFF_3_QD), .A2(n253), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3334)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2644), .A2(KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n253), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2963), .A2(n253), .ZN(KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS22ser[3]), .A2(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n210), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[3]), .A2(n210), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2963) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2669), .A2(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n210), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2740), .A2(n210), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS22ser[4]), .A2(KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n255), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S22reg_gff_1_SFF_4_QD), .A2(n255), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3335)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2647), .A2(KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n255), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2964), .A2(n255), .ZN(KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS22ser[4]), .A2(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n314), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[4]), .A2(n314), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2964) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2672), .A2(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n314), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2743), .A2(n314), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS22ser[5]), .A2(KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n257), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S22reg_gff_1_SFF_5_QD), .A2(n257), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3336)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2650), .A2(KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n257), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2965), .A2(n257), .ZN(KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS22ser[5]), .A2(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[5]), .A2(n193), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2965) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2675), .A2(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2746), .A2(n193), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS22ser[6]), .A2(KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n252), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S22reg_gff_1_SFF_6_QD), .A2(n252), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3337)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2653), .A2(KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n252), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2966), .A2(n252), .ZN(KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS22ser[6]), .A2(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n198), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[6]), .A2(n198), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2966) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2678), .A2(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n198), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2749), .A2(n198), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS22ser[7]), .A2(KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n258), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S22reg_gff_1_SFF_7_QD), .A2(n258), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3338)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2656), .A2(KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n258), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2967), .A2(n258), .ZN(KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS22ser[7]), .A2(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[7]), .A2(n197), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2967) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2681), .A2(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2752), .A2(n197), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS23ser[0]), .A2(KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n263), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S23reg_gff_1_SFF_0_QD), .A2(n263), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3339)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2659), .A2(KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n263), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2968), .A2(n263), .ZN(KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS23ser[0]), .A2(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n319), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[0]), .A2(n319), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2968) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2684), .A2(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n319), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2755), .A2(n319), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS23ser[1]), .A2(KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n251), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S23reg_gff_1_SFF_1_QD), .A2(n251), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3340)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2662), .A2(KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n251), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2969), .A2(n251), .ZN(KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS23ser[1]), .A2(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n197), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[1]), .A2(n197), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2969) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2687), .A2(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n197), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2758), .A2(n197), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS23ser[2]), .A2(KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n256), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S23reg_gff_1_SFF_2_QD), .A2(n256), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3341)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2665), .A2(KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n256), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2970), .A2(n256), .ZN(KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS23ser[2]), .A2(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[2]), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2970) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2690), .A2(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2761), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS23ser[3]), .A2(KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n265), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S23reg_gff_1_SFF_3_QD), .A2(n265), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3342)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2668), .A2(KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n265), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2971), .A2(n265), .ZN(KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS23ser[3]), .A2(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[3]), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2971) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2693), .A2(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2764), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS23ser[4]), .A2(KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n268), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S23reg_gff_1_SFF_4_QD), .A2(n268), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3343)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2671), .A2(KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n268), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2972), .A2(n268), .ZN(KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS23ser[4]), .A2(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[4]), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2972) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2696), .A2(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2767), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_n5) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS23ser[5]), .A2(KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n262), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S23reg_gff_1_SFF_5_QD), .A2(n262), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3344)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2674), .A2(KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n262), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2973), .A2(n262), .ZN(KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS23ser[5]), .A2(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[5]), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2973) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2699), .A2(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2770), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_n5) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS23ser[6]), .A2(KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S23reg_gff_1_SFF_6_QD), .A2(n204), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3345)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2677), .A2(KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2974), .A2(n204), .ZN(KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS23ser[6]), .A2(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[6]), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2974) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2702), .A2(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2773), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_n5) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS23ser[7]), .A2(KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n261), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S23reg_gff_1_SFF_7_QD), .A2(n261), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3346)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2680), .A2(KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n261), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2975), .A2(n261), .ZN(KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS23ser[7]), .A2(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[7]), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2975) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2705), .A2(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2776), .A2(n199), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS31ser[0]), .A2(KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n257), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S31reg_gff_1_SFF_0_QD), .A2(n257), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3347)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2707), .A2(KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n257), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2976), .A2(n257), .ZN(KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS31ser[0]), .A2(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_0_), .A2(n199), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2976) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2732), .A2(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2020), .A2(n199), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS31ser[1]), .A2(KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n258), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S31reg_gff_1_SFF_1_QD), .A2(n258), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3348)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2710), .A2(KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n258), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2977), .A2(n258), .ZN(KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS31ser[1]), .A2(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n199), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_1_), .A2(n199), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2977) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2735), .A2(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n199), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2018), .A2(n199), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS31ser[2]), .A2(KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n264), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S31reg_gff_1_SFF_2_QD), .A2(n264), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3349)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2713), .A2(KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n264), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2978), .A2(n264), .ZN(KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS31ser[2]), .A2(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_2_), .A2(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2978) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2738), .A2(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2016), .A2(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS31ser[3]), .A2(KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n259), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S31reg_gff_1_SFF_3_QD), .A2(n259), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3350)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2716), .A2(KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n259), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2979), .A2(n259), .ZN(KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS31ser[3]), .A2(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_3_), .A2(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2979) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2741), .A2(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2014), .A2(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS31ser[4]), .A2(KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n268), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S31reg_gff_1_SFF_4_QD), .A2(n268), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3351)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2719), .A2(KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n268), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2980), .A2(n268), .ZN(KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS31ser[4]), .A2(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_4_), .A2(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2980) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2744), .A2(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2012), .A2(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS31ser[5]), .A2(KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S31reg_gff_1_SFF_5_QD), .A2(n204), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3352)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2722), .A2(KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2981), .A2(n204), .ZN(KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS31ser[5]), .A2(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n321), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_5_), .A2(n321), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2981) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2747), .A2(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n321), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2010), .A2(n321), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS31ser[6]), .A2(KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S31reg_gff_1_SFF_6_QD), .A2(n204), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3353)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2725), .A2(KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2982), .A2(n204), .ZN(KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS31ser[6]), .A2(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_6_), .A2(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2982) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2750), .A2(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2008), .A2(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS31ser[7]), .A2(KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n264), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S31reg_gff_1_SFF_7_QD), .A2(n264), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3354)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2728), .A2(KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n264), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2983), .A2(n264), .ZN(KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS31ser[7]), .A2(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_7_), .A2(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2983) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2753), .A2(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2006), .A2(n200), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS32ser[0]), .A2(KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S32reg_gff_1_SFF_0_QD), .A2(n204), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3355)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2731), .A2(KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2984), .A2(n204), .ZN(KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS32ser[0]), .A2(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[0]), .A2(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2984) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2756), .A2(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2443), .A2(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS32ser[1]), .A2(KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n253), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S32reg_gff_1_SFF_1_QD), .A2(n253), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3356)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2734), .A2(KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n253), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2985), .A2(n253), .ZN(KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS32ser[1]), .A2(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[1]), .A2(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2985) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2759), .A2(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2446), .A2(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS32ser[2]), .A2(KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n204), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S32reg_gff_1_SFF_2_QD), .A2(n204), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3357)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2737), .A2(KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n204), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2986), .A2(n204), .ZN(KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS32ser[2]), .A2(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[2]), .A2(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2986) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2762), .A2(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2449), .A2(n200), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS32ser[3]), .A2(KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n266), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S32reg_gff_1_SFF_3_QD), .A2(n266), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3358)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2740), .A2(KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n266), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2987), .A2(n266), .ZN(KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS32ser[3]), .A2(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[3]), .A2(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2987) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2765), .A2(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2452), .A2(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS32ser[4]), .A2(KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n261), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S32reg_gff_1_SFF_4_QD), .A2(n261), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3359)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2743), .A2(KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n261), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2988), .A2(n261), .ZN(KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS32ser[4]), .A2(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[4]), .A2(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2988) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2768), .A2(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2455), .A2(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS32ser[5]), .A2(KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n263), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S32reg_gff_1_SFF_5_QD), .A2(n263), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3360)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2746), .A2(KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n263), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2989), .A2(n263), .ZN(KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS32ser[5]), .A2(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[5]), .A2(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2989) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2771), .A2(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2458), .A2(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_n5) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS32ser[6]), .A2(KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n252), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S32reg_gff_1_SFF_6_QD), .A2(n252), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3361)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2749), .A2(KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n252), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2990), .A2(n252), .ZN(KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS32ser[6]), .A2(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[6]), .A2(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2990) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2774), .A2(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2461), .A2(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_n5) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS32ser[7]), .A2(KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n254), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S32reg_gff_1_SFF_7_QD), .A2(n254), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3362)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2752), .A2(KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n254), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2991), .A2(n254), .ZN(KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS32ser[7]), .A2(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[7]), .A2(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2991) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2777), .A2(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2464), .A2(n196), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_n5) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(KeyArray_outS33ser[0]), .A2(KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n252), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S33reg_gff_1_SFF_0_QD), .A2(n252), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3363)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2755), .A2(KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n252), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2992), .A2(n252), .ZN(KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS33ser[0]), .A2(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[0]), .A2(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2992) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2779), .A2(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2467), .A2(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_n5) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(KeyArray_outS33ser[1]), .A2(KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n269), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S33reg_gff_1_SFF_1_QD), .A2(n269), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3364)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2758), .A2(KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n269), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2993), .A2(n269), .ZN(KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS33ser[1]), .A2(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[1]), .A2(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2993) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2781), .A2(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2470), .A2(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_n5) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(KeyArray_outS33ser[2]), .A2(KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n266), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S33reg_gff_1_SFF_2_QD), .A2(n266), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3365)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2761), .A2(KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n266), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2994), .A2(n266), .ZN(KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS33ser[2]), .A2(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[2]), .A2(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2994) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2783), .A2(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2473), .A2(n196), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_n5) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(KeyArray_outS33ser[3]), .A2(KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n266), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S33reg_gff_1_SFF_3_QD), .A2(n266), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3366)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2764), .A2(KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n266), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2995), .A2(n266), .ZN(KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS33ser[3]), .A2(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n190), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[3]), .A2(n190), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2995) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2785), .A2(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n190), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2476), .A2(n190), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_n5) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(KeyArray_outS33ser[4]), .A2(KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n266), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S33reg_gff_1_SFF_4_QD), .A2(n266), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3367)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2767), .A2(KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n266), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2996), .A2(n266), .ZN(KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS33ser[4]), .A2(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n314), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[4]), .A2(n314), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2996) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2787), .A2(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n314), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2479), .A2(n314), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_n5) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(KeyArray_outS33ser[5]), .A2(KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n264), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S33reg_gff_1_SFF_5_QD), .A2(n264), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3368)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2770), .A2(KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n264), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2997), .A2(n264), .ZN(KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS33ser[5]), .A2(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n318), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[5]), .A2(n318), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2997) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2789), .A2(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n318), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2482), .A2(n318), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_n5) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(KeyArray_outS33ser[6]), .A2(KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n254), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S33reg_gff_1_SFF_6_QD), .A2(n254), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3369)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2773), .A2(KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n254), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2998), .A2(n254), .ZN(KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS33ser[6]), .A2(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n193), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[6]), .A2(n193), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2998) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2791), .A2(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n193), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2485), .A2(n193), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_n5) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(KeyArray_outS33ser[7]), .A2(KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n263), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S33reg_gff_1_SFF_7_QD), .A2(n263), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3370)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2776), .A2(KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n263), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2999), .A2(n263), .ZN(KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        KeyArray_inS33ser[7]), .A2(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n318), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[7]), .A2(n318), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2999) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2793), .A2(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n318), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2488), .A2(n318), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_outS01ser_p[0]) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_U3 ( .A1(
        KeyArray_outS01ser_0_), .A2(KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_XOR_00[0]), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3109) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2020), .A2(KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2021), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_outS01ser_p[1]) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_U3 ( .A1(
        KeyArray_outS01ser_1_), .A2(KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_XOR_00[1]), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3110) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2018), .A2(KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2019), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_outS01ser_p[2]) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_U3 ( .A1(
        KeyArray_outS01ser_2_), .A2(KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_XOR_00[2]), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3111) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2016), .A2(KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2017), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_outS01ser_p[3]) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_U3 ( .A1(
        KeyArray_outS01ser_3_), .A2(KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_XOR_00[3]), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3112) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2014), .A2(KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2015), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_outS01ser_p[4]) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_U3 ( .A1(
        KeyArray_outS01ser_4_), .A2(KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_XOR_00[4]), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3113) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2012), .A2(KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2013), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_outS01ser_p[5]) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_U3 ( .A1(
        KeyArray_outS01ser_5_), .A2(KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_XOR_00[5]), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3114) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2010), .A2(KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2011), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_outS01ser_p[6]) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_U3 ( .A1(
        KeyArray_outS01ser_6_), .A2(KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_XOR_00[6]), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3115) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2008), .A2(KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2009), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_outS01ser_p[7]) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_U3 ( .A1(
        KeyArray_outS01ser_7_), .A2(KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_XOR_00[7]), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3116) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_2006), .A2(KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_n6), .ZN(KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_U2 ( .A(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2007), .A2(n288), .ZN(
        KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS00ser[0]) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[120]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_U2 ( .A(n191), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_p[0]), .A2(n191), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3247) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[120]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_U2 ( .A(n191), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3109), .A2(n191), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS00ser[1]) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[121]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_U2 ( .A(n304), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_p[1]), .A2(n304), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3249) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[121]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_U2 ( .A(n304), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3110), .A2(n304), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS00ser[2]) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[122]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_U2 ( .A(n303), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_p[2]), .A2(n303), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3251) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[122]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_U2 ( .A(n303), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3111), .A2(n303), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS00ser[3]) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[123]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_U2 ( .A(n302), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_p[3]), .A2(n302), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3253) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[123]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_U2 ( .A(n302), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3112), .A2(n302), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS00ser[4]) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[124]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_U2 ( .A(n299), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_p[4]), .A2(n299), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3255) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[124]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_U2 ( .A(n299), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3113), .A2(n299), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS00ser[5]) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[125]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_U2 ( .A(n301), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_p[5]), .A2(n301), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3257) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[125]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_U2 ( .A(n301), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3114), .A2(n301), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS00ser[6]) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[126]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_U2 ( .A(n296), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_p[6]), .A2(n296), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3259) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[126]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_U2 ( .A(n296), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3115), .A2(n296), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS00ser[7]) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[127]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_U2 ( .A(n291), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS01ser_p[7]), .A2(n291), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3261) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[127]),
        .A2(KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_U2 ( .A(n291), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3116), .A2(n291), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS01ser[0]) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[112]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_U2 ( .A(n191), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[0]), .A2(n191), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2444) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[112]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_U2 ( .A(n191), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2443), .A2(n191), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS01ser[1]) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[113]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[1]), .A2(n307), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2447) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[113]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2446), .A2(n307), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS01ser[2]) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[114]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[2]), .A2(n308), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2450) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[114]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2449), .A2(n308), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS01ser[3]) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[115]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[3]), .A2(n194), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2453) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[115]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2452), .A2(n194), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS01ser[4]) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[116]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[4]), .A2(n310), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2456) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[116]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2455), .A2(n310), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS01ser[5]) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[117]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[5]), .A2(n195), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2459) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[117]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2458), .A2(n195), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS01ser[6]) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[118]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[6]), .A2(n307), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2462) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[118]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2461), .A2(n307), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS01ser[7]) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[119]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS02ser[7]), .A2(n308), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2465) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[119]),
        .A2(KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2464), .A2(n308), .ZN(
        KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS02ser[0]) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[104]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[0]), .A2(n310), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2468) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[104]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2467), .A2(n310), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS02ser[1]) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[105]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_U2 ( .A(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[1]), .A2(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2471) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[105]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_U2 ( .A(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2470), .A2(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS02ser[2]) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[106]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_U2 ( .A(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[2]), .A2(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2474) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[106]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_U2 ( .A(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2473), .A2(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS02ser[3]) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[107]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_U2 ( .A(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[3]), .A2(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2477) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[107]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_U2 ( .A(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2476), .A2(n14), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS02ser[4]) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[108]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[4]), .A2(n195), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2480) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[108]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2479), .A2(n195), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS02ser[5]) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[109]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[5]), .A2(n295), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2483) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[109]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2482), .A2(n295), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS02ser[6]) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[110]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[6]), .A2(n195), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2486) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[110]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2485), .A2(n195), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS02ser[7]) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[111]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS03ser[7]), .A2(n311), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2489) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[111]),
        .A2(KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2488), .A2(n311), .ZN(
        KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS03ser[0]) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[96]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[0]), .A2(n309), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2492) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[96]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2491), .A2(n309), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS03ser[1]) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[97]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_U2 ( .A(n312), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[1]), .A2(n312), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2495) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[97]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_U2 ( .A(n312), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2494), .A2(n312), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS03ser[2]) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[98]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_U2 ( .A(n292), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[2]), .A2(n292), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2498) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[98]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_U2 ( .A(n292), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2497), .A2(n292), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS03ser[3]) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[99]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[3]), .A2(n194), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2501) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[99]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2500), .A2(n194), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS03ser[4]) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[100]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_U2 ( .A(n293), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[4]), .A2(n293), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2504) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[100]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_U2 ( .A(n293), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2503), .A2(n293), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS03ser[5]) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[101]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_U2 ( .A(n294), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[5]), .A2(n294), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2507) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[101]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_U2 ( .A(n294), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2506), .A2(n294), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS03ser[6]) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[102]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_U2 ( .A(n294), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[6]), .A2(n294), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2510) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[102]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_U2 ( .A(n294), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2509), .A2(n294), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS03ser[7]) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[103]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS10ser[7]), .A2(n311), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2513) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[103]),
        .A2(KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2512), .A2(n311), .ZN(
        KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS10ser[0]) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[88]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[0]), .A2(n309), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2516) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[88]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2515), .A2(n309), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS10ser[1]) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[89]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[1]), .A2(n195), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2519) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[89]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2518), .A2(n195), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS10ser[2]) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[90]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_U2 ( .A(n312), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[2]), .A2(n312), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2522) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[90]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_U2 ( .A(n312), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2521), .A2(n312), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS10ser[3]) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[91]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[3]), .A2(n194), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2525) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[91]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2524), .A2(n194), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS10ser[4]) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[92]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[4]), .A2(n195), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2528) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[92]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2527), .A2(n195), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS10ser[5]) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[93]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_U2 ( .A(n294), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[5]), .A2(n294), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2531) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[93]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_U2 ( .A(n294), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2530), .A2(n294), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS10ser[6]) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[94]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[6]), .A2(n194), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2534) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[94]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2533), .A2(n194), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS10ser[7]) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[95]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_U2 ( .A(n293), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS11ser[7]), .A2(n293), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2537) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[95]),
        .A2(KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_U2 ( .A(n293), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2536), .A2(n293), .ZN(
        KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS11ser[0]) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[80]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[0]), .A2(n311), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2540) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[80]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2539), .A2(n311), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS11ser[1]) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[81]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[1]), .A2(n195), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2543) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[81]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_U2 ( .A(n195), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2542), .A2(n195), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS11ser[2]) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[82]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_U2 ( .A(n292), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[2]), .A2(n292), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2546) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[82]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_U2 ( .A(n292), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2545), .A2(n292), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS11ser[3]) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[83]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_U2 ( .A(n298), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[3]), .A2(n298), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2549) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[83]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_U2 ( .A(n298), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2548), .A2(n298), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS11ser[4]) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[84]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[4]), .A2(n311), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2552) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[84]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2551), .A2(n311), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS11ser[5]) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[85]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_U2 ( .A(n297), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[5]), .A2(n297), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2555) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[85]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_U2 ( .A(n297), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2554), .A2(n297), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS11ser[6]) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[86]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[6]), .A2(n310), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2558) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[86]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2557), .A2(n310), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS11ser[7]) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[87]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS12ser[7]), .A2(n306), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2561) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[87]),
        .A2(KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2560), .A2(n306), .ZN(
        KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS12ser[0]) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[72]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_U2 ( .A(n191), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_U1 ( .A1(keySBIn[0]),
        .A2(n191), .ZN(KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2564) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[72]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_U2 ( .A(n191), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2563), .A2(n191), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS12ser[1]) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[73]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_U2 ( .A(n304), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_U1 ( .A1(keySBIn[1]),
        .A2(n304), .ZN(KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2567) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[73]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_U2 ( .A(n304), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2566), .A2(n304), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS12ser[2]) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[74]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_U2 ( .A(n301), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_U1 ( .A1(keySBIn[2]),
        .A2(n301), .ZN(KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2570) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[74]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_U2 ( .A(n301), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2569), .A2(n301), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS12ser[3]) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[75]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_U2 ( .A(n305), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_U1 ( .A1(keySBIn[3]),
        .A2(n305), .ZN(KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2573) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[75]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_U2 ( .A(n305), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2572), .A2(n305), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS12ser[4]) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[76]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_U2 ( .A(n304), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_U1 ( .A1(keySBIn[4]),
        .A2(n304), .ZN(KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2576) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[76]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_U2 ( .A(n304), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2575), .A2(n304), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS12ser[5]) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[77]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_U2 ( .A(n291), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_U1 ( .A1(keySBIn[5]),
        .A2(n291), .ZN(KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2579) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[77]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_U2 ( .A(n291), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2578), .A2(n291), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS12ser[6]) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[78]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_U2 ( .A(n291), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_U1 ( .A1(keySBIn[6]),
        .A2(n291), .ZN(KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2582) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[78]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_U2 ( .A(n291), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2581), .A2(n291), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS12ser[7]) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[79]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_U2 ( .A(n305), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_U1 ( .A1(keySBIn[7]),
        .A2(n305), .ZN(KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2585) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[79]),
        .A2(KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_U2 ( .A(n305), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2584), .A2(n305), .ZN(
        KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS13ser[0]) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[64]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[0]), .A2(n309), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2588) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[64]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2587), .A2(n309), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS13ser[1]) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[65]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[1]), .A2(n306), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2591) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[65]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2590), .A2(n306), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS13ser[2]) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[66]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[2]), .A2(n295), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2594) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[66]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2593), .A2(n295), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS13ser[3]) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[67]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[3]), .A2(n310), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2597) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[67]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2596), .A2(n310), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS13ser[4]) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[68]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_U2 ( .A(n292), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[4]), .A2(n292), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2600) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[68]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_U2 ( .A(n292), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2599), .A2(n292), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS13ser[5]) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[69]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[5]), .A2(n295), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2603) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[69]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2602), .A2(n295), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS13ser[6]) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[70]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[6]), .A2(n306), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2606) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[70]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2605), .A2(n306), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS13ser[7]) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[71]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_U2 ( .A(n293), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS20ser[7]), .A2(n293), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2609) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[71]),
        .A2(KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_U2 ( .A(n293), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2608), .A2(n293), .ZN(
        KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS20ser[0]) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[56]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_U2 ( .A(n312), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[0]), .A2(n312), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2612) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[56]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_U2 ( .A(n312), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2611), .A2(n312), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS20ser[1]) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[57]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_U2 ( .A(n293), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[1]), .A2(n293), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2615) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[57]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_U2 ( .A(n293), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2614), .A2(n293), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS20ser[2]) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[58]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[2]), .A2(n307), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2618) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[58]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2617), .A2(n307), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS20ser[3]) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[59]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[3]), .A2(n194), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2621) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[59]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2620), .A2(n194), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS20ser[4]) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[60]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_U2 ( .A(n293), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[4]), .A2(n293), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2624) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[60]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_U2 ( .A(n293), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2623), .A2(n293), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS20ser[5]) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[61]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[5]), .A2(n306), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2627) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[61]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2626), .A2(n306), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS20ser[6]) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[62]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[6]), .A2(n309), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2630) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[62]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2629), .A2(n309), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS20ser[7]) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[63]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS21ser[7]), .A2(n308), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2633) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[63]),
        .A2(KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2632), .A2(n308), .ZN(
        KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS21ser[0]) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[48]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[0]), .A2(n307), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2636) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[48]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2635), .A2(n307), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS21ser[1]) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[49]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_U2 ( .A(n312), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[1]), .A2(n312), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2639) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[49]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_U2 ( .A(n312), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2638), .A2(n312), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS21ser[2]) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[50]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[2]), .A2(n310), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2642) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[50]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2641), .A2(n310), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS21ser[3]) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[51]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[3]), .A2(n310), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2645) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[51]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_U2 ( .A(n310), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2644), .A2(n310), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS21ser[4]) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[52]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[4]), .A2(n306), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2648) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[52]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2647), .A2(n306), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS21ser[5]) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[53]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[5]), .A2(n308), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2651) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[53]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2650), .A2(n308), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS21ser[6]) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[54]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_U2 ( .A(n292), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[6]), .A2(n292), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2654) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[54]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_U2 ( .A(n292), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2653), .A2(n292), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS21ser[7]) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[55]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS22ser[7]), .A2(n309), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2657) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[55]),
        .A2(KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2656), .A2(n309), .ZN(
        KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS22ser[0]) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[40]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[0]), .A2(n307), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2660) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[40]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2659), .A2(n307), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS22ser[1]) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[41]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[1]), .A2(n194), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2663) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[41]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_U2 ( .A(n194), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2662), .A2(n194), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS22ser[2]) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[42]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[2]), .A2(n295), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2666) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[42]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2665), .A2(n295), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS22ser[3]) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[43]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_U2 ( .A(n312), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[3]), .A2(n312), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2669) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[43]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_U2 ( .A(n312), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2668), .A2(n312), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS22ser[4]) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[44]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[4]), .A2(n308), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2672) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[44]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2671), .A2(n308), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS22ser[5]) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[45]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_U2 ( .A(n300), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[5]), .A2(n300), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2675) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[45]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_U2 ( .A(n300), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2674), .A2(n300), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS22ser[6]) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[46]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_U2 ( .A(n294), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[6]), .A2(n294), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2678) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[46]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_U2 ( .A(n294), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2677), .A2(n294), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS22ser[7]) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[47]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS23ser[7]), .A2(n295), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2681) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[47]),
        .A2(KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2680), .A2(n295), .ZN(
        KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS23ser[0]) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[32]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[0]), .A2(n308), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2684) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[32]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_U2 ( .A(n308), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2683), .A2(n308), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS23ser[1]) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[33]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[1]), .A2(n295), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2687) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[33]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2686), .A2(n295), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS23ser[2]) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[34]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[2]), .A2(n311), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2690) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[34]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2689), .A2(n311), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS23ser[3]) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[35]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[3]), .A2(n307), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2693) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[35]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_U2 ( .A(n307), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2692), .A2(n307), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS23ser[4]) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[36]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_U2 ( .A(n292), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[4]), .A2(n292), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2696) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[36]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_U2 ( .A(n292), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2695), .A2(n292), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS23ser[5]) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[37]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[5]), .A2(n309), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2699) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[37]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_U2 ( .A(n309), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2698), .A2(n309), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS23ser[6]) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[38]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[6]), .A2(n311), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2702) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[38]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_U2 ( .A(n311), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2701), .A2(n311), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS23ser[7]) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[39]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS30ser[7]), .A2(n306), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2705) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[39]),
        .A2(KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_U2 ( .A(n306), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2704), .A2(n306), .ZN(
        KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS30ser[0]) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[24]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[0]), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2708) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[24]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2707), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS30ser[1]) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[25]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[1]), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2711) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[25]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2710), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS30ser[2]) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[26]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[2]), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2714) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[26]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2713), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS30ser[3]) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[27]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[3]), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2717) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[27]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2716), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS30ser[4]) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[28]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[4]), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2720) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[28]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2719), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS30ser[5]) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[29]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[5]), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2723) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[29]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2722), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS30ser[6]) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[30]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[6]), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2726) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[30]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2725), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS30ser[7]) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[31]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS31ser[7]), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2729) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[31]),
        .A2(KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_U2 ( .A(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2728), .A2(n295), .ZN(
        KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS31ser[0]) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[16]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_U2 ( .A(n304), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[0]), .A2(n304), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2732) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[16]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_U2 ( .A(n304), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2731), .A2(n304), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS31ser[1]) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[17]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_U2 ( .A(n303), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[1]), .A2(n303), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2735) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[17]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_U2 ( .A(n303), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2734), .A2(n303), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS31ser[2]) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[18]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_U2 ( .A(n299), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[2]), .A2(n299), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2738) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[18]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_U2 ( .A(n299), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2737), .A2(n299), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS31ser[3]) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[19]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_U2 ( .A(n302), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[3]), .A2(n302), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2741) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[19]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_U2 ( .A(n302), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2740), .A2(n302), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS31ser[4]) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[20]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_U2 ( .A(n298), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[4]), .A2(n298), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2744) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[20]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_U2 ( .A(n298), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2743), .A2(n298), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS31ser[5]) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[21]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_U2 ( .A(n300), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[5]), .A2(n300), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2747) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[21]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_U2 ( .A(n300), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2746), .A2(n300), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS31ser[6]) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[22]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_U2 ( .A(n302), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[6]), .A2(n302), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2750) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[22]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_U2 ( .A(n302), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2749), .A2(n302), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS31ser[7]) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[23]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_U2 ( .A(n297), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS32ser[7]), .A2(n297), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2753) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[23]),
        .A2(KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_U2 ( .A(n297), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2752), .A2(n297), .ZN(
        KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS32ser[0]) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[8]), .A2(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_U2 ( .A(n299), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[0]), .A2(n299), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2756) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[8]), .A2(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_U2 ( .A(n299), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2755), .A2(n299), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS32ser[1]) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[9]), .A2(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_U2 ( .A(n303), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[1]), .A2(n303), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2759) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[9]), .A2(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_U2 ( .A(n303), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2758), .A2(n303), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS32ser[2]) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[10]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_U2 ( .A(n301), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[2]), .A2(n301), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2762) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[10]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_U2 ( .A(n301), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2761), .A2(n301), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS32ser[3]) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[11]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_U2 ( .A(n297), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[3]), .A2(n297), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2765) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[11]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_U2 ( .A(n297), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2764), .A2(n297), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS32ser[4]) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[12]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_U2 ( .A(n298), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[4]), .A2(n298), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2768) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[12]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_U2 ( .A(n298), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2767), .A2(n298), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS32ser[5]) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[13]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_U2 ( .A(n296), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[5]), .A2(n296), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2771) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[13]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_U2 ( .A(n296), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2770), .A2(n296), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS32ser[6]) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[14]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_U2 ( .A(n291), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[6]), .A2(n291), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2774) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[14]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_U2 ( .A(n291), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2773), .A2(n291), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS32ser[7]) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[15]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_U2 ( .A(n305), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        KeyArray_outS33ser[7]), .A2(n305), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2777) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[15]),
        .A2(KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_U2 ( .A(n305), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2776), .A2(n305), .ZN(
        KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        KeyArray_inS33ser[0]) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_U3 ( .A1(key_s0[0]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_U2 ( .A(n303), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_U1 ( .A1(keyStateIn[0]),
        .A2(n303), .ZN(KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2779) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_U3 ( .A1(key_s1[0]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_U2 ( .A(n303), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_1983), .A2(n303), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        KeyArray_inS33ser[1]) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_U3 ( .A1(key_s0[1]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_U2 ( .A(n302), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_U1 ( .A1(keyStateIn[1]),
        .A2(n302), .ZN(KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2781) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_U3 ( .A1(key_s1[1]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_U2 ( .A(n302), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_1986), .A2(n302), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        KeyArray_inS33ser[2]) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_U3 ( .A1(key_s0[2]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_U2 ( .A(n299), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_U1 ( .A1(keyStateIn[2]),
        .A2(n299), .ZN(KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2783) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_U3 ( .A1(key_s1[2]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_U2 ( .A(n299), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_1989), .A2(n299), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        KeyArray_inS33ser[3]) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_U3 ( .A1(key_s0[3]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_U2 ( .A(n300), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_U1 ( .A1(keyStateIn[3]),
        .A2(n300), .ZN(KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2785) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_U3 ( .A1(key_s1[3]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_U2 ( .A(n300), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_1992), .A2(n300), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        KeyArray_inS33ser[4]) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_U3 ( .A1(key_s0[4]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_U2 ( .A(n298), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_U1 ( .A1(keyStateIn[4]),
        .A2(n298), .ZN(KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2787) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_U3 ( .A1(key_s1[4]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_U2 ( .A(n298), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_1995), .A2(n298), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        KeyArray_inS33ser[5]) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_U3 ( .A1(key_s0[5]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_U2 ( .A(n297), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_U1 ( .A1(keyStateIn[5]),
        .A2(n297), .ZN(KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2789) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_U3 ( .A1(key_s1[5]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_U2 ( .A(n297), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_1998), .A2(n297), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        KeyArray_inS33ser[6]) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_U3 ( .A1(key_s0[6]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_U2 ( .A(n296), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_U1 ( .A1(keyStateIn[6]),
        .A2(n296), .ZN(KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2791) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_U3 ( .A1(key_s1[6]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_U2 ( .A(n296), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2001), .A2(n296), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        KeyArray_inS33ser[7]) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_U3 ( .A1(key_s0[7]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_U2 ( .A(n305), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_U1 ( .A1(keyStateIn[7]),
        .A2(n305), .ZN(KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n8), .A2(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_2793) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_U3 ( .A1(key_s1[7]), .A2(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_U2 ( .A(n305), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_2004), .A2(n305), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n8) );
  XNOR2_X1 MixColumns_line0_U24_Ins0_U1 ( .A(MixColumns_line0_n16), .B(
        MixColumns_line0_n15), .ZN(MCout[31]) );
  XOR2_X1 MixColumns_line0_U24_Ins_1_U1 ( .A(new_AGEMA_signal_2122), .B(
        new_AGEMA_signal_2024), .Z(new_AGEMA_signal_2794) );
  XNOR2_X1 MixColumns_line0_U23_Ins0_U1 ( .A(ciphertext_s0[63]), .B(
        ciphertext_s0[31]), .ZN(MixColumns_line0_n15) );
  XOR2_X1 MixColumns_line0_U23_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        ciphertext_s1[31]), .Z(new_AGEMA_signal_2024) );
  XOR2_X1 MixColumns_line0_U22_Ins_0_U1 ( .A(ciphertext_s0[126]), .B(
        MixColumns_line0_S13[7]), .Z(MixColumns_line0_n16) );
  XOR2_X1 MixColumns_line0_U22_Ins_1_U1 ( .A(ciphertext_s1[126]), .B(
        new_AGEMA_signal_2051), .Z(new_AGEMA_signal_2122) );
  XNOR2_X1 MixColumns_line0_U21_Ins0_U1 ( .A(MixColumns_line0_n14), .B(
        MixColumns_line0_n13), .ZN(MCout[30]) );
  XOR2_X1 MixColumns_line0_U21_Ins_1_U1 ( .A(new_AGEMA_signal_2123), .B(
        new_AGEMA_signal_2027), .Z(new_AGEMA_signal_2795) );
  XNOR2_X1 MixColumns_line0_U20_Ins0_U1 ( .A(ciphertext_s0[62]), .B(
        ciphertext_s0[30]), .ZN(MixColumns_line0_n13) );
  XOR2_X1 MixColumns_line0_U20_Ins_1_U1 ( .A(ciphertext_s1[62]), .B(
        ciphertext_s1[30]), .Z(new_AGEMA_signal_2027) );
  XOR2_X1 MixColumns_line0_U19_Ins_0_U1 ( .A(ciphertext_s0[125]), .B(
        MixColumns_line0_S13[6]), .Z(MixColumns_line0_n14) );
  XOR2_X1 MixColumns_line0_U19_Ins_1_U1 ( .A(ciphertext_s1[125]), .B(
        new_AGEMA_signal_2053), .Z(new_AGEMA_signal_2123) );
  XNOR2_X1 MixColumns_line0_U18_Ins0_U1 ( .A(MixColumns_line0_n12), .B(
        MixColumns_line0_n11), .ZN(MCout[29]) );
  XOR2_X1 MixColumns_line0_U18_Ins_1_U1 ( .A(new_AGEMA_signal_2124), .B(
        new_AGEMA_signal_2030), .Z(new_AGEMA_signal_2796) );
  XNOR2_X1 MixColumns_line0_U17_Ins0_U1 ( .A(ciphertext_s0[61]), .B(
        ciphertext_s0[29]), .ZN(MixColumns_line0_n11) );
  XOR2_X1 MixColumns_line0_U17_Ins_1_U1 ( .A(ciphertext_s1[61]), .B(
        ciphertext_s1[29]), .Z(new_AGEMA_signal_2030) );
  XOR2_X1 MixColumns_line0_U16_Ins_0_U1 ( .A(ciphertext_s0[124]), .B(
        MixColumns_line0_S13[5]), .Z(MixColumns_line0_n12) );
  XOR2_X1 MixColumns_line0_U16_Ins_1_U1 ( .A(ciphertext_s1[124]), .B(
        new_AGEMA_signal_2055), .Z(new_AGEMA_signal_2124) );
  XNOR2_X1 MixColumns_line0_U15_Ins0_U1 ( .A(MixColumns_line0_n10), .B(
        MixColumns_line0_n9), .ZN(MCout[28]) );
  XOR2_X1 MixColumns_line0_U15_Ins_1_U1 ( .A(new_AGEMA_signal_2797), .B(
        new_AGEMA_signal_2033), .Z(new_AGEMA_signal_2838) );
  XNOR2_X1 MixColumns_line0_U14_Ins0_U1 ( .A(ciphertext_s0[60]), .B(
        ciphertext_s0[28]), .ZN(MixColumns_line0_n9) );
  XOR2_X1 MixColumns_line0_U14_Ins_1_U1 ( .A(ciphertext_s1[60]), .B(
        ciphertext_s1[28]), .Z(new_AGEMA_signal_2033) );
  XOR2_X1 MixColumns_line0_U13_Ins_0_U1 ( .A(MixColumns_line0_S02[4]), .B(
        MixColumns_line0_S13[4]), .Z(MixColumns_line0_n10) );
  XOR2_X1 MixColumns_line0_U13_Ins_1_U1 ( .A(new_AGEMA_signal_2046), .B(
        new_AGEMA_signal_2127), .Z(new_AGEMA_signal_2797) );
  XNOR2_X1 MixColumns_line0_U12_Ins0_U1 ( .A(MixColumns_line0_n8), .B(
        MixColumns_line0_n7), .ZN(MCout[27]) );
  XOR2_X1 MixColumns_line0_U12_Ins_1_U1 ( .A(new_AGEMA_signal_2798), .B(
        new_AGEMA_signal_2036), .Z(new_AGEMA_signal_2839) );
  XNOR2_X1 MixColumns_line0_U11_Ins0_U1 ( .A(ciphertext_s0[59]), .B(
        ciphertext_s0[27]), .ZN(MixColumns_line0_n7) );
  XOR2_X1 MixColumns_line0_U11_Ins_1_U1 ( .A(ciphertext_s1[59]), .B(
        ciphertext_s1[27]), .Z(new_AGEMA_signal_2036) );
  XOR2_X1 MixColumns_line0_U10_Ins_0_U1 ( .A(MixColumns_line0_S02[3]), .B(
        MixColumns_line0_S13[3]), .Z(MixColumns_line0_n8) );
  XOR2_X1 MixColumns_line0_U10_Ins_1_U1 ( .A(new_AGEMA_signal_2047), .B(
        new_AGEMA_signal_2128), .Z(new_AGEMA_signal_2798) );
  XNOR2_X1 MixColumns_line0_U9_Ins0_U1 ( .A(MixColumns_line0_n6), .B(
        MixColumns_line0_n5), .ZN(MCout[26]) );
  XOR2_X1 MixColumns_line0_U9_Ins_1_U1 ( .A(new_AGEMA_signal_2125), .B(
        new_AGEMA_signal_2039), .Z(new_AGEMA_signal_2799) );
  XNOR2_X1 MixColumns_line0_U8_Ins0_U1 ( .A(ciphertext_s0[58]), .B(
        ciphertext_s0[26]), .ZN(MixColumns_line0_n5) );
  XOR2_X1 MixColumns_line0_U8_Ins_1_U1 ( .A(ciphertext_s1[58]), .B(
        ciphertext_s1[26]), .Z(new_AGEMA_signal_2039) );
  XOR2_X1 MixColumns_line0_U7_Ins_0_U1 ( .A(ciphertext_s0[121]), .B(
        MixColumns_line0_S13[2]), .Z(MixColumns_line0_n6) );
  XOR2_X1 MixColumns_line0_U7_Ins_1_U1 ( .A(ciphertext_s1[121]), .B(
        new_AGEMA_signal_2058), .Z(new_AGEMA_signal_2125) );
  XNOR2_X1 MixColumns_line0_U6_Ins0_U1 ( .A(MixColumns_line0_n4), .B(
        MixColumns_line0_n3), .ZN(MCout[25]) );
  XOR2_X1 MixColumns_line0_U6_Ins_1_U1 ( .A(new_AGEMA_signal_2800), .B(
        new_AGEMA_signal_2042), .Z(new_AGEMA_signal_2840) );
  XNOR2_X1 MixColumns_line0_U5_Ins0_U1 ( .A(ciphertext_s0[25]), .B(
        ciphertext_s0[57]), .ZN(MixColumns_line0_n3) );
  XOR2_X1 MixColumns_line0_U5_Ins_1_U1 ( .A(ciphertext_s1[25]), .B(
        ciphertext_s1[57]), .Z(new_AGEMA_signal_2042) );
  XOR2_X1 MixColumns_line0_U4_Ins_0_U1 ( .A(MixColumns_line0_S02_1), .B(
        MixColumns_line0_S13[1]), .Z(MixColumns_line0_n4) );
  XOR2_X1 MixColumns_line0_U4_Ins_1_U1 ( .A(new_AGEMA_signal_2048), .B(
        new_AGEMA_signal_2129), .Z(new_AGEMA_signal_2800) );
  XNOR2_X1 MixColumns_line0_U3_Ins0_U1 ( .A(MixColumns_line0_n2), .B(
        MixColumns_line0_n1), .ZN(MCout[24]) );
  XOR2_X1 MixColumns_line0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2126), .B(
        new_AGEMA_signal_2045), .Z(new_AGEMA_signal_2801) );
  XNOR2_X1 MixColumns_line0_U2_Ins0_U1 ( .A(ciphertext_s0[24]), .B(
        ciphertext_s0[56]), .ZN(MixColumns_line0_n1) );
  XOR2_X1 MixColumns_line0_U2_Ins_1_U1 ( .A(ciphertext_s1[24]), .B(
        ciphertext_s1[56]), .Z(new_AGEMA_signal_2045) );
  XOR2_X1 MixColumns_line0_U1_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(
        MixColumns_line0_S13[0]), .Z(MixColumns_line0_n2) );
  XOR2_X1 MixColumns_line0_U1_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(
        new_AGEMA_signal_2060), .Z(new_AGEMA_signal_2126) );
  XOR2_X1 MixColumns_line0_timesTWO_U3_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(
        ciphertext_s0[123]), .Z(MixColumns_line0_S02[4]) );
  XOR2_X1 MixColumns_line0_timesTWO_U3_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(
        ciphertext_s1[123]), .Z(new_AGEMA_signal_2046) );
  XOR2_X1 MixColumns_line0_timesTWO_U2_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(
        ciphertext_s0[122]), .Z(MixColumns_line0_S02[3]) );
  XOR2_X1 MixColumns_line0_timesTWO_U2_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(
        ciphertext_s1[122]), .Z(new_AGEMA_signal_2047) );
  XOR2_X1 MixColumns_line0_timesTWO_U1_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(
        ciphertext_s0[120]), .Z(MixColumns_line0_S02_1) );
  XOR2_X1 MixColumns_line0_timesTWO_U1_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(
        ciphertext_s1[120]), .Z(new_AGEMA_signal_2048) );
  XOR2_X1 MixColumns_line0_timesTHREE_U8_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(
        ciphertext_s0[94]), .Z(MixColumns_line0_S13[7]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U8_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        ciphertext_s1[94]), .Z(new_AGEMA_signal_2051) );
  XOR2_X1 MixColumns_line0_timesTHREE_U7_Ins_0_U1 ( .A(ciphertext_s0[94]), .B(
        ciphertext_s0[93]), .Z(MixColumns_line0_S13[6]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U7_Ins_1_U1 ( .A(ciphertext_s1[94]), .B(
        ciphertext_s1[93]), .Z(new_AGEMA_signal_2053) );
  XOR2_X1 MixColumns_line0_timesTHREE_U6_Ins_0_U1 ( .A(ciphertext_s0[93]), .B(
        ciphertext_s0[92]), .Z(MixColumns_line0_S13[5]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U6_Ins_1_U1 ( .A(ciphertext_s1[93]), .B(
        ciphertext_s1[92]), .Z(new_AGEMA_signal_2055) );
  XOR2_X1 MixColumns_line0_timesTHREE_U5_Ins_0_U1 ( .A(ciphertext_s0[92]), .B(
        MixColumns_line0_timesTHREE_input2[4]), .Z(MixColumns_line0_S13[4]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U5_Ins_1_U1 ( .A(ciphertext_s1[92]), .B(
        new_AGEMA_signal_2062), .Z(new_AGEMA_signal_2127) );
  XOR2_X1 MixColumns_line0_timesTHREE_U4_Ins_0_U1 ( .A(ciphertext_s0[91]), .B(
        MixColumns_line0_timesTHREE_input2[3]), .Z(MixColumns_line0_S13[3]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U4_Ins_1_U1 ( .A(ciphertext_s1[91]), .B(
        new_AGEMA_signal_2063), .Z(new_AGEMA_signal_2128) );
  XOR2_X1 MixColumns_line0_timesTHREE_U3_Ins_0_U1 ( .A(ciphertext_s0[90]), .B(
        ciphertext_s0[89]), .Z(MixColumns_line0_S13[2]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U3_Ins_1_U1 ( .A(ciphertext_s1[90]), .B(
        ciphertext_s1[89]), .Z(new_AGEMA_signal_2058) );
  XOR2_X1 MixColumns_line0_timesTHREE_U2_Ins_0_U1 ( .A(ciphertext_s0[89]), .B(
        MixColumns_line0_timesTHREE_input2_1), .Z(MixColumns_line0_S13[1]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U2_Ins_1_U1 ( .A(ciphertext_s1[89]), .B(
        new_AGEMA_signal_2064), .Z(new_AGEMA_signal_2129) );
  XOR2_X1 MixColumns_line0_timesTHREE_U1_Ins_0_U1 ( .A(ciphertext_s0[88]), .B(
        ciphertext_s0[95]), .Z(MixColumns_line0_S13[0]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U1_Ins_1_U1 ( .A(ciphertext_s1[88]), .B(
        ciphertext_s1[95]), .Z(new_AGEMA_signal_2060) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U3_Ins_0_U1 ( .A(
        ciphertext_s0[95]), .B(ciphertext_s0[91]), .Z(
        MixColumns_line0_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U3_Ins_1_U1 ( .A(
        ciphertext_s1[95]), .B(ciphertext_s1[91]), .Z(new_AGEMA_signal_2062)
         );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U2_Ins_0_U1 ( .A(
        ciphertext_s0[95]), .B(ciphertext_s0[90]), .Z(
        MixColumns_line0_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U2_Ins_1_U1 ( .A(
        ciphertext_s1[95]), .B(ciphertext_s1[90]), .Z(new_AGEMA_signal_2063)
         );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U1_Ins_0_U1 ( .A(
        ciphertext_s0[95]), .B(ciphertext_s0[88]), .Z(
        MixColumns_line0_timesTHREE_input2_1) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U1_Ins_1_U1 ( .A(
        ciphertext_s1[95]), .B(ciphertext_s1[88]), .Z(new_AGEMA_signal_2064)
         );
  XNOR2_X1 MixColumns_line1_U24_Ins0_U1 ( .A(MixColumns_line1_n16), .B(
        MixColumns_line1_n15), .ZN(MCout[23]) );
  XOR2_X1 MixColumns_line1_U24_Ins_1_U1 ( .A(new_AGEMA_signal_2130), .B(
        new_AGEMA_signal_2065), .Z(new_AGEMA_signal_2802) );
  XNOR2_X1 MixColumns_line1_U23_Ins0_U1 ( .A(ciphertext_s0[31]), .B(
        ciphertext_s0[127]), .ZN(MixColumns_line1_n15) );
  XOR2_X1 MixColumns_line1_U23_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        ciphertext_s1[127]), .Z(new_AGEMA_signal_2065) );
  XOR2_X1 MixColumns_line1_U22_Ins_0_U1 ( .A(ciphertext_s0[94]), .B(
        MixColumns_line1_S13[7]), .Z(MixColumns_line1_n16) );
  XOR2_X1 MixColumns_line1_U22_Ins_1_U1 ( .A(ciphertext_s1[94]), .B(
        new_AGEMA_signal_2076), .Z(new_AGEMA_signal_2130) );
  XNOR2_X1 MixColumns_line1_U21_Ins0_U1 ( .A(MixColumns_line1_n14), .B(
        MixColumns_line1_n13), .ZN(MCout[22]) );
  XOR2_X1 MixColumns_line1_U21_Ins_1_U1 ( .A(new_AGEMA_signal_2131), .B(
        new_AGEMA_signal_2066), .Z(new_AGEMA_signal_2803) );
  XNOR2_X1 MixColumns_line1_U20_Ins0_U1 ( .A(ciphertext_s0[30]), .B(
        ciphertext_s0[126]), .ZN(MixColumns_line1_n13) );
  XOR2_X1 MixColumns_line1_U20_Ins_1_U1 ( .A(ciphertext_s1[30]), .B(
        ciphertext_s1[126]), .Z(new_AGEMA_signal_2066) );
  XOR2_X1 MixColumns_line1_U19_Ins_0_U1 ( .A(ciphertext_s0[93]), .B(
        MixColumns_line1_S13[6]), .Z(MixColumns_line1_n14) );
  XOR2_X1 MixColumns_line1_U19_Ins_1_U1 ( .A(ciphertext_s1[93]), .B(
        new_AGEMA_signal_2077), .Z(new_AGEMA_signal_2131) );
  XNOR2_X1 MixColumns_line1_U18_Ins0_U1 ( .A(MixColumns_line1_n12), .B(
        MixColumns_line1_n11), .ZN(MCout[21]) );
  XOR2_X1 MixColumns_line1_U18_Ins_1_U1 ( .A(new_AGEMA_signal_2132), .B(
        new_AGEMA_signal_2067), .Z(new_AGEMA_signal_2804) );
  XNOR2_X1 MixColumns_line1_U17_Ins0_U1 ( .A(ciphertext_s0[29]), .B(
        ciphertext_s0[125]), .ZN(MixColumns_line1_n11) );
  XOR2_X1 MixColumns_line1_U17_Ins_1_U1 ( .A(ciphertext_s1[29]), .B(
        ciphertext_s1[125]), .Z(new_AGEMA_signal_2067) );
  XOR2_X1 MixColumns_line1_U16_Ins_0_U1 ( .A(ciphertext_s0[92]), .B(
        MixColumns_line1_S13[5]), .Z(MixColumns_line1_n12) );
  XOR2_X1 MixColumns_line1_U16_Ins_1_U1 ( .A(ciphertext_s1[92]), .B(
        new_AGEMA_signal_2078), .Z(new_AGEMA_signal_2132) );
  XNOR2_X1 MixColumns_line1_U15_Ins0_U1 ( .A(MixColumns_line1_n10), .B(
        MixColumns_line1_n9), .ZN(MCout[20]) );
  XOR2_X1 MixColumns_line1_U15_Ins_1_U1 ( .A(new_AGEMA_signal_2805), .B(
        new_AGEMA_signal_2068), .Z(new_AGEMA_signal_2841) );
  XNOR2_X1 MixColumns_line1_U14_Ins0_U1 ( .A(ciphertext_s0[28]), .B(
        ciphertext_s0[124]), .ZN(MixColumns_line1_n9) );
  XOR2_X1 MixColumns_line1_U14_Ins_1_U1 ( .A(ciphertext_s1[28]), .B(
        ciphertext_s1[124]), .Z(new_AGEMA_signal_2068) );
  XOR2_X1 MixColumns_line1_U13_Ins_0_U1 ( .A(MixColumns_line1_S02_4_), .B(
        MixColumns_line1_S13[4]), .Z(MixColumns_line1_n10) );
  XOR2_X1 MixColumns_line1_U13_Ins_1_U1 ( .A(new_AGEMA_signal_2073), .B(
        new_AGEMA_signal_2135), .Z(new_AGEMA_signal_2805) );
  XNOR2_X1 MixColumns_line1_U12_Ins0_U1 ( .A(MixColumns_line1_n8), .B(
        MixColumns_line1_n7), .ZN(MCout[19]) );
  XOR2_X1 MixColumns_line1_U12_Ins_1_U1 ( .A(new_AGEMA_signal_2806), .B(
        new_AGEMA_signal_2069), .Z(new_AGEMA_signal_2842) );
  XNOR2_X1 MixColumns_line1_U11_Ins0_U1 ( .A(ciphertext_s0[27]), .B(
        ciphertext_s0[123]), .ZN(MixColumns_line1_n7) );
  XOR2_X1 MixColumns_line1_U11_Ins_1_U1 ( .A(ciphertext_s1[27]), .B(
        ciphertext_s1[123]), .Z(new_AGEMA_signal_2069) );
  XOR2_X1 MixColumns_line1_U10_Ins_0_U1 ( .A(MixColumns_line1_S02_3_), .B(
        MixColumns_line1_S13[3]), .Z(MixColumns_line1_n8) );
  XOR2_X1 MixColumns_line1_U10_Ins_1_U1 ( .A(new_AGEMA_signal_2074), .B(
        new_AGEMA_signal_2136), .Z(new_AGEMA_signal_2806) );
  XNOR2_X1 MixColumns_line1_U9_Ins0_U1 ( .A(MixColumns_line1_n6), .B(
        MixColumns_line1_n5), .ZN(MCout[18]) );
  XOR2_X1 MixColumns_line1_U9_Ins_1_U1 ( .A(new_AGEMA_signal_2133), .B(
        new_AGEMA_signal_2070), .Z(new_AGEMA_signal_2807) );
  XNOR2_X1 MixColumns_line1_U8_Ins0_U1 ( .A(ciphertext_s0[26]), .B(
        ciphertext_s0[122]), .ZN(MixColumns_line1_n5) );
  XOR2_X1 MixColumns_line1_U8_Ins_1_U1 ( .A(ciphertext_s1[26]), .B(
        ciphertext_s1[122]), .Z(new_AGEMA_signal_2070) );
  XOR2_X1 MixColumns_line1_U7_Ins_0_U1 ( .A(ciphertext_s0[89]), .B(
        MixColumns_line1_S13[2]), .Z(MixColumns_line1_n6) );
  XOR2_X1 MixColumns_line1_U7_Ins_1_U1 ( .A(ciphertext_s1[89]), .B(
        new_AGEMA_signal_2079), .Z(new_AGEMA_signal_2133) );
  XNOR2_X1 MixColumns_line1_U6_Ins0_U1 ( .A(MixColumns_line1_n4), .B(
        MixColumns_line1_n3), .ZN(MCout[17]) );
  XOR2_X1 MixColumns_line1_U6_Ins_1_U1 ( .A(new_AGEMA_signal_2808), .B(
        new_AGEMA_signal_2071), .Z(new_AGEMA_signal_2843) );
  XNOR2_X1 MixColumns_line1_U5_Ins0_U1 ( .A(ciphertext_s0[121]), .B(
        ciphertext_s0[25]), .ZN(MixColumns_line1_n3) );
  XOR2_X1 MixColumns_line1_U5_Ins_1_U1 ( .A(ciphertext_s1[121]), .B(
        ciphertext_s1[25]), .Z(new_AGEMA_signal_2071) );
  XOR2_X1 MixColumns_line1_U4_Ins_0_U1 ( .A(MixColumns_line1_S02_1_), .B(
        MixColumns_line1_S13[1]), .Z(MixColumns_line1_n4) );
  XOR2_X1 MixColumns_line1_U4_Ins_1_U1 ( .A(new_AGEMA_signal_2075), .B(
        new_AGEMA_signal_2137), .Z(new_AGEMA_signal_2808) );
  XNOR2_X1 MixColumns_line1_U3_Ins0_U1 ( .A(MixColumns_line1_n2), .B(
        MixColumns_line1_n1), .ZN(MCout[16]) );
  XOR2_X1 MixColumns_line1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2134), .B(
        new_AGEMA_signal_2072), .Z(new_AGEMA_signal_2809) );
  XNOR2_X1 MixColumns_line1_U2_Ins0_U1 ( .A(ciphertext_s0[120]), .B(
        ciphertext_s0[24]), .ZN(MixColumns_line1_n1) );
  XOR2_X1 MixColumns_line1_U2_Ins_1_U1 ( .A(ciphertext_s1[120]), .B(
        ciphertext_s1[24]), .Z(new_AGEMA_signal_2072) );
  XOR2_X1 MixColumns_line1_U1_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(
        MixColumns_line1_S13[0]), .Z(MixColumns_line1_n2) );
  XOR2_X1 MixColumns_line1_U1_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        new_AGEMA_signal_2080), .Z(new_AGEMA_signal_2134) );
  XOR2_X1 MixColumns_line1_timesTWO_U3_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(
        ciphertext_s0[91]), .Z(MixColumns_line1_S02_4_) );
  XOR2_X1 MixColumns_line1_timesTWO_U3_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        ciphertext_s1[91]), .Z(new_AGEMA_signal_2073) );
  XOR2_X1 MixColumns_line1_timesTWO_U2_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(
        ciphertext_s0[90]), .Z(MixColumns_line1_S02_3_) );
  XOR2_X1 MixColumns_line1_timesTWO_U2_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        ciphertext_s1[90]), .Z(new_AGEMA_signal_2074) );
  XOR2_X1 MixColumns_line1_timesTWO_U1_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(
        ciphertext_s0[88]), .Z(MixColumns_line1_S02_1_) );
  XOR2_X1 MixColumns_line1_timesTWO_U1_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        ciphertext_s1[88]), .Z(new_AGEMA_signal_2075) );
  XOR2_X1 MixColumns_line1_timesTHREE_U8_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(
        ciphertext_s0[62]), .Z(MixColumns_line1_S13[7]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U8_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        ciphertext_s1[62]), .Z(new_AGEMA_signal_2076) );
  XOR2_X1 MixColumns_line1_timesTHREE_U7_Ins_0_U1 ( .A(ciphertext_s0[62]), .B(
        ciphertext_s0[61]), .Z(MixColumns_line1_S13[6]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U7_Ins_1_U1 ( .A(ciphertext_s1[62]), .B(
        ciphertext_s1[61]), .Z(new_AGEMA_signal_2077) );
  XOR2_X1 MixColumns_line1_timesTHREE_U6_Ins_0_U1 ( .A(ciphertext_s0[61]), .B(
        ciphertext_s0[60]), .Z(MixColumns_line1_S13[5]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U6_Ins_1_U1 ( .A(ciphertext_s1[61]), .B(
        ciphertext_s1[60]), .Z(new_AGEMA_signal_2078) );
  XOR2_X1 MixColumns_line1_timesTHREE_U5_Ins_0_U1 ( .A(ciphertext_s0[60]), .B(
        MixColumns_line1_timesTHREE_input2[4]), .Z(MixColumns_line1_S13[4]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U5_Ins_1_U1 ( .A(ciphertext_s1[60]), .B(
        new_AGEMA_signal_2081), .Z(new_AGEMA_signal_2135) );
  XOR2_X1 MixColumns_line1_timesTHREE_U4_Ins_0_U1 ( .A(ciphertext_s0[59]), .B(
        MixColumns_line1_timesTHREE_input2[3]), .Z(MixColumns_line1_S13[3]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U4_Ins_1_U1 ( .A(ciphertext_s1[59]), .B(
        new_AGEMA_signal_2082), .Z(new_AGEMA_signal_2136) );
  XOR2_X1 MixColumns_line1_timesTHREE_U3_Ins_0_U1 ( .A(ciphertext_s0[58]), .B(
        ciphertext_s0[57]), .Z(MixColumns_line1_S13[2]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U3_Ins_1_U1 ( .A(ciphertext_s1[58]), .B(
        ciphertext_s1[57]), .Z(new_AGEMA_signal_2079) );
  XOR2_X1 MixColumns_line1_timesTHREE_U2_Ins_0_U1 ( .A(ciphertext_s0[57]), .B(
        MixColumns_line1_timesTHREE_input2_1), .Z(MixColumns_line1_S13[1]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U2_Ins_1_U1 ( .A(ciphertext_s1[57]), .B(
        new_AGEMA_signal_2083), .Z(new_AGEMA_signal_2137) );
  XOR2_X1 MixColumns_line1_timesTHREE_U1_Ins_0_U1 ( .A(ciphertext_s0[56]), .B(
        ciphertext_s0[63]), .Z(MixColumns_line1_S13[0]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U1_Ins_1_U1 ( .A(ciphertext_s1[56]), .B(
        ciphertext_s1[63]), .Z(new_AGEMA_signal_2080) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U3_Ins_0_U1 ( .A(
        ciphertext_s0[63]), .B(ciphertext_s0[59]), .Z(
        MixColumns_line1_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U3_Ins_1_U1 ( .A(
        ciphertext_s1[63]), .B(ciphertext_s1[59]), .Z(new_AGEMA_signal_2081)
         );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U2_Ins_0_U1 ( .A(
        ciphertext_s0[63]), .B(ciphertext_s0[58]), .Z(
        MixColumns_line1_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U2_Ins_1_U1 ( .A(
        ciphertext_s1[63]), .B(ciphertext_s1[58]), .Z(new_AGEMA_signal_2082)
         );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U1_Ins_0_U1 ( .A(
        ciphertext_s0[63]), .B(ciphertext_s0[56]), .Z(
        MixColumns_line1_timesTHREE_input2_1) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U1_Ins_1_U1 ( .A(
        ciphertext_s1[63]), .B(ciphertext_s1[56]), .Z(new_AGEMA_signal_2083)
         );
  XNOR2_X1 MixColumns_line2_U24_Ins0_U1 ( .A(MixColumns_line2_n16), .B(
        MixColumns_line2_n15), .ZN(MCout[15]) );
  XOR2_X1 MixColumns_line2_U24_Ins_1_U1 ( .A(new_AGEMA_signal_2138), .B(
        new_AGEMA_signal_2084), .Z(new_AGEMA_signal_2810) );
  XNOR2_X1 MixColumns_line2_U23_Ins0_U1 ( .A(ciphertext_s0[127]), .B(
        ciphertext_s0[95]), .ZN(MixColumns_line2_n15) );
  XOR2_X1 MixColumns_line2_U23_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(
        ciphertext_s1[95]), .Z(new_AGEMA_signal_2084) );
  XOR2_X1 MixColumns_line2_U22_Ins_0_U1 ( .A(ciphertext_s0[62]), .B(
        MixColumns_line2_S13[7]), .Z(MixColumns_line2_n16) );
  XOR2_X1 MixColumns_line2_U22_Ins_1_U1 ( .A(ciphertext_s1[62]), .B(
        new_AGEMA_signal_2095), .Z(new_AGEMA_signal_2138) );
  XNOR2_X1 MixColumns_line2_U21_Ins0_U1 ( .A(MixColumns_line2_n14), .B(
        MixColumns_line2_n13), .ZN(MCout[14]) );
  XOR2_X1 MixColumns_line2_U21_Ins_1_U1 ( .A(new_AGEMA_signal_2139), .B(
        new_AGEMA_signal_2085), .Z(new_AGEMA_signal_2811) );
  XNOR2_X1 MixColumns_line2_U20_Ins0_U1 ( .A(ciphertext_s0[126]), .B(
        ciphertext_s0[94]), .ZN(MixColumns_line2_n13) );
  XOR2_X1 MixColumns_line2_U20_Ins_1_U1 ( .A(ciphertext_s1[126]), .B(
        ciphertext_s1[94]), .Z(new_AGEMA_signal_2085) );
  XOR2_X1 MixColumns_line2_U19_Ins_0_U1 ( .A(ciphertext_s0[61]), .B(
        MixColumns_line2_S13[6]), .Z(MixColumns_line2_n14) );
  XOR2_X1 MixColumns_line2_U19_Ins_1_U1 ( .A(ciphertext_s1[61]), .B(
        new_AGEMA_signal_2096), .Z(new_AGEMA_signal_2139) );
  XNOR2_X1 MixColumns_line2_U18_Ins0_U1 ( .A(MixColumns_line2_n12), .B(
        MixColumns_line2_n11), .ZN(MCout[13]) );
  XOR2_X1 MixColumns_line2_U18_Ins_1_U1 ( .A(new_AGEMA_signal_2140), .B(
        new_AGEMA_signal_2086), .Z(new_AGEMA_signal_2812) );
  XNOR2_X1 MixColumns_line2_U17_Ins0_U1 ( .A(ciphertext_s0[125]), .B(
        ciphertext_s0[93]), .ZN(MixColumns_line2_n11) );
  XOR2_X1 MixColumns_line2_U17_Ins_1_U1 ( .A(ciphertext_s1[125]), .B(
        ciphertext_s1[93]), .Z(new_AGEMA_signal_2086) );
  XOR2_X1 MixColumns_line2_U16_Ins_0_U1 ( .A(ciphertext_s0[60]), .B(
        MixColumns_line2_S13[5]), .Z(MixColumns_line2_n12) );
  XOR2_X1 MixColumns_line2_U16_Ins_1_U1 ( .A(ciphertext_s1[60]), .B(
        new_AGEMA_signal_2097), .Z(new_AGEMA_signal_2140) );
  XNOR2_X1 MixColumns_line2_U15_Ins0_U1 ( .A(MixColumns_line2_n10), .B(
        MixColumns_line2_n9), .ZN(MCout[12]) );
  XOR2_X1 MixColumns_line2_U15_Ins_1_U1 ( .A(new_AGEMA_signal_2813), .B(
        new_AGEMA_signal_2087), .Z(new_AGEMA_signal_2844) );
  XNOR2_X1 MixColumns_line2_U14_Ins0_U1 ( .A(ciphertext_s0[124]), .B(
        ciphertext_s0[92]), .ZN(MixColumns_line2_n9) );
  XOR2_X1 MixColumns_line2_U14_Ins_1_U1 ( .A(ciphertext_s1[124]), .B(
        ciphertext_s1[92]), .Z(new_AGEMA_signal_2087) );
  XOR2_X1 MixColumns_line2_U13_Ins_0_U1 ( .A(MixColumns_line2_S02_4_), .B(
        MixColumns_line2_S13[4]), .Z(MixColumns_line2_n10) );
  XOR2_X1 MixColumns_line2_U13_Ins_1_U1 ( .A(new_AGEMA_signal_2092), .B(
        new_AGEMA_signal_2143), .Z(new_AGEMA_signal_2813) );
  XNOR2_X1 MixColumns_line2_U12_Ins0_U1 ( .A(MixColumns_line2_n8), .B(
        MixColumns_line2_n7), .ZN(MCout[11]) );
  XOR2_X1 MixColumns_line2_U12_Ins_1_U1 ( .A(new_AGEMA_signal_2814), .B(
        new_AGEMA_signal_2088), .Z(new_AGEMA_signal_2845) );
  XNOR2_X1 MixColumns_line2_U11_Ins0_U1 ( .A(ciphertext_s0[123]), .B(
        ciphertext_s0[91]), .ZN(MixColumns_line2_n7) );
  XOR2_X1 MixColumns_line2_U11_Ins_1_U1 ( .A(ciphertext_s1[123]), .B(
        ciphertext_s1[91]), .Z(new_AGEMA_signal_2088) );
  XOR2_X1 MixColumns_line2_U10_Ins_0_U1 ( .A(MixColumns_line2_S02_3_), .B(
        MixColumns_line2_S13[3]), .Z(MixColumns_line2_n8) );
  XOR2_X1 MixColumns_line2_U10_Ins_1_U1 ( .A(new_AGEMA_signal_2093), .B(
        new_AGEMA_signal_2144), .Z(new_AGEMA_signal_2814) );
  XNOR2_X1 MixColumns_line2_U9_Ins0_U1 ( .A(MixColumns_line2_n6), .B(
        MixColumns_line2_n5), .ZN(MCout[10]) );
  XOR2_X1 MixColumns_line2_U9_Ins_1_U1 ( .A(new_AGEMA_signal_2141), .B(
        new_AGEMA_signal_2089), .Z(new_AGEMA_signal_2815) );
  XNOR2_X1 MixColumns_line2_U8_Ins0_U1 ( .A(ciphertext_s0[122]), .B(
        ciphertext_s0[90]), .ZN(MixColumns_line2_n5) );
  XOR2_X1 MixColumns_line2_U8_Ins_1_U1 ( .A(ciphertext_s1[122]), .B(
        ciphertext_s1[90]), .Z(new_AGEMA_signal_2089) );
  XOR2_X1 MixColumns_line2_U7_Ins_0_U1 ( .A(ciphertext_s0[57]), .B(
        MixColumns_line2_S13[2]), .Z(MixColumns_line2_n6) );
  XOR2_X1 MixColumns_line2_U7_Ins_1_U1 ( .A(ciphertext_s1[57]), .B(
        new_AGEMA_signal_2098), .Z(new_AGEMA_signal_2141) );
  XNOR2_X1 MixColumns_line2_U6_Ins0_U1 ( .A(MixColumns_line2_n4), .B(
        MixColumns_line2_n3), .ZN(MCout[9]) );
  XOR2_X1 MixColumns_line2_U6_Ins_1_U1 ( .A(new_AGEMA_signal_2816), .B(
        new_AGEMA_signal_2090), .Z(new_AGEMA_signal_2846) );
  XNOR2_X1 MixColumns_line2_U5_Ins0_U1 ( .A(ciphertext_s0[89]), .B(
        ciphertext_s0[121]), .ZN(MixColumns_line2_n3) );
  XOR2_X1 MixColumns_line2_U5_Ins_1_U1 ( .A(ciphertext_s1[89]), .B(
        ciphertext_s1[121]), .Z(new_AGEMA_signal_2090) );
  XOR2_X1 MixColumns_line2_U4_Ins_0_U1 ( .A(MixColumns_line2_S02_1_), .B(
        MixColumns_line2_S13[1]), .Z(MixColumns_line2_n4) );
  XOR2_X1 MixColumns_line2_U4_Ins_1_U1 ( .A(new_AGEMA_signal_2094), .B(
        new_AGEMA_signal_2145), .Z(new_AGEMA_signal_2816) );
  XNOR2_X1 MixColumns_line2_U3_Ins0_U1 ( .A(MixColumns_line2_n2), .B(
        MixColumns_line2_n1), .ZN(MCout[8]) );
  XOR2_X1 MixColumns_line2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2142), .B(
        new_AGEMA_signal_2091), .Z(new_AGEMA_signal_2817) );
  XNOR2_X1 MixColumns_line2_U2_Ins0_U1 ( .A(ciphertext_s0[88]), .B(
        ciphertext_s0[120]), .ZN(MixColumns_line2_n1) );
  XOR2_X1 MixColumns_line2_U2_Ins_1_U1 ( .A(ciphertext_s1[88]), .B(
        ciphertext_s1[120]), .Z(new_AGEMA_signal_2091) );
  XOR2_X1 MixColumns_line2_U1_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(
        MixColumns_line2_S13[0]), .Z(MixColumns_line2_n2) );
  XOR2_X1 MixColumns_line2_U1_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        new_AGEMA_signal_2099), .Z(new_AGEMA_signal_2142) );
  XOR2_X1 MixColumns_line2_timesTWO_U3_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(
        ciphertext_s0[59]), .Z(MixColumns_line2_S02_4_) );
  XOR2_X1 MixColumns_line2_timesTWO_U3_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        ciphertext_s1[59]), .Z(new_AGEMA_signal_2092) );
  XOR2_X1 MixColumns_line2_timesTWO_U2_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(
        ciphertext_s0[58]), .Z(MixColumns_line2_S02_3_) );
  XOR2_X1 MixColumns_line2_timesTWO_U2_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        ciphertext_s1[58]), .Z(new_AGEMA_signal_2093) );
  XOR2_X1 MixColumns_line2_timesTWO_U1_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(
        ciphertext_s0[56]), .Z(MixColumns_line2_S02_1_) );
  XOR2_X1 MixColumns_line2_timesTWO_U1_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        ciphertext_s1[56]), .Z(new_AGEMA_signal_2094) );
  XOR2_X1 MixColumns_line2_timesTHREE_U8_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(
        ciphertext_s0[30]), .Z(MixColumns_line2_S13[7]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U8_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        ciphertext_s1[30]), .Z(new_AGEMA_signal_2095) );
  XOR2_X1 MixColumns_line2_timesTHREE_U7_Ins_0_U1 ( .A(ciphertext_s0[30]), .B(
        ciphertext_s0[29]), .Z(MixColumns_line2_S13[6]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U7_Ins_1_U1 ( .A(ciphertext_s1[30]), .B(
        ciphertext_s1[29]), .Z(new_AGEMA_signal_2096) );
  XOR2_X1 MixColumns_line2_timesTHREE_U6_Ins_0_U1 ( .A(ciphertext_s0[29]), .B(
        ciphertext_s0[28]), .Z(MixColumns_line2_S13[5]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U6_Ins_1_U1 ( .A(ciphertext_s1[29]), .B(
        ciphertext_s1[28]), .Z(new_AGEMA_signal_2097) );
  XOR2_X1 MixColumns_line2_timesTHREE_U5_Ins_0_U1 ( .A(ciphertext_s0[28]), .B(
        MixColumns_line2_timesTHREE_input2[4]), .Z(MixColumns_line2_S13[4]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U5_Ins_1_U1 ( .A(ciphertext_s1[28]), .B(
        new_AGEMA_signal_2100), .Z(new_AGEMA_signal_2143) );
  XOR2_X1 MixColumns_line2_timesTHREE_U4_Ins_0_U1 ( .A(ciphertext_s0[27]), .B(
        MixColumns_line2_timesTHREE_input2[3]), .Z(MixColumns_line2_S13[3]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U4_Ins_1_U1 ( .A(ciphertext_s1[27]), .B(
        new_AGEMA_signal_2101), .Z(new_AGEMA_signal_2144) );
  XOR2_X1 MixColumns_line2_timesTHREE_U3_Ins_0_U1 ( .A(ciphertext_s0[26]), .B(
        ciphertext_s0[25]), .Z(MixColumns_line2_S13[2]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U3_Ins_1_U1 ( .A(ciphertext_s1[26]), .B(
        ciphertext_s1[25]), .Z(new_AGEMA_signal_2098) );
  XOR2_X1 MixColumns_line2_timesTHREE_U2_Ins_0_U1 ( .A(ciphertext_s0[25]), .B(
        MixColumns_line2_timesTHREE_input2_1), .Z(MixColumns_line2_S13[1]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U2_Ins_1_U1 ( .A(ciphertext_s1[25]), .B(
        new_AGEMA_signal_2102), .Z(new_AGEMA_signal_2145) );
  XOR2_X1 MixColumns_line2_timesTHREE_U1_Ins_0_U1 ( .A(ciphertext_s0[24]), .B(
        ciphertext_s0[31]), .Z(MixColumns_line2_S13[0]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U1_Ins_1_U1 ( .A(ciphertext_s1[24]), .B(
        ciphertext_s1[31]), .Z(new_AGEMA_signal_2099) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U3_Ins_0_U1 ( .A(
        ciphertext_s0[31]), .B(ciphertext_s0[27]), .Z(
        MixColumns_line2_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U3_Ins_1_U1 ( .A(
        ciphertext_s1[31]), .B(ciphertext_s1[27]), .Z(new_AGEMA_signal_2100)
         );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U2_Ins_0_U1 ( .A(
        ciphertext_s0[31]), .B(ciphertext_s0[26]), .Z(
        MixColumns_line2_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U2_Ins_1_U1 ( .A(
        ciphertext_s1[31]), .B(ciphertext_s1[26]), .Z(new_AGEMA_signal_2101)
         );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U1_Ins_0_U1 ( .A(
        ciphertext_s0[31]), .B(ciphertext_s0[24]), .Z(
        MixColumns_line2_timesTHREE_input2_1) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U1_Ins_1_U1 ( .A(
        ciphertext_s1[31]), .B(ciphertext_s1[24]), .Z(new_AGEMA_signal_2102)
         );
  XNOR2_X1 MixColumns_line3_U24_Ins0_U1 ( .A(MixColumns_line3_n16), .B(
        MixColumns_line3_n15), .ZN(MCout[7]) );
  XOR2_X1 MixColumns_line3_U24_Ins_1_U1 ( .A(new_AGEMA_signal_2146), .B(
        new_AGEMA_signal_2103), .Z(new_AGEMA_signal_2818) );
  XNOR2_X1 MixColumns_line3_U23_Ins0_U1 ( .A(ciphertext_s0[95]), .B(
        ciphertext_s0[63]), .ZN(MixColumns_line3_n15) );
  XOR2_X1 MixColumns_line3_U23_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        ciphertext_s1[63]), .Z(new_AGEMA_signal_2103) );
  XOR2_X1 MixColumns_line3_U22_Ins_0_U1 ( .A(ciphertext_s0[30]), .B(
        MixColumns_line3_S13[7]), .Z(MixColumns_line3_n16) );
  XOR2_X1 MixColumns_line3_U22_Ins_1_U1 ( .A(ciphertext_s1[30]), .B(
        new_AGEMA_signal_2114), .Z(new_AGEMA_signal_2146) );
  XNOR2_X1 MixColumns_line3_U21_Ins0_U1 ( .A(MixColumns_line3_n14), .B(
        MixColumns_line3_n13), .ZN(MCout[6]) );
  XOR2_X1 MixColumns_line3_U21_Ins_1_U1 ( .A(new_AGEMA_signal_2147), .B(
        new_AGEMA_signal_2104), .Z(new_AGEMA_signal_2819) );
  XNOR2_X1 MixColumns_line3_U20_Ins0_U1 ( .A(ciphertext_s0[94]), .B(
        ciphertext_s0[62]), .ZN(MixColumns_line3_n13) );
  XOR2_X1 MixColumns_line3_U20_Ins_1_U1 ( .A(ciphertext_s1[94]), .B(
        ciphertext_s1[62]), .Z(new_AGEMA_signal_2104) );
  XOR2_X1 MixColumns_line3_U19_Ins_0_U1 ( .A(ciphertext_s0[29]), .B(
        MixColumns_line3_S13[6]), .Z(MixColumns_line3_n14) );
  XOR2_X1 MixColumns_line3_U19_Ins_1_U1 ( .A(ciphertext_s1[29]), .B(
        new_AGEMA_signal_2115), .Z(new_AGEMA_signal_2147) );
  XNOR2_X1 MixColumns_line3_U18_Ins0_U1 ( .A(MixColumns_line3_n12), .B(
        MixColumns_line3_n11), .ZN(MCout[5]) );
  XOR2_X1 MixColumns_line3_U18_Ins_1_U1 ( .A(new_AGEMA_signal_2148), .B(
        new_AGEMA_signal_2105), .Z(new_AGEMA_signal_2820) );
  XNOR2_X1 MixColumns_line3_U17_Ins0_U1 ( .A(ciphertext_s0[93]), .B(
        ciphertext_s0[61]), .ZN(MixColumns_line3_n11) );
  XOR2_X1 MixColumns_line3_U17_Ins_1_U1 ( .A(ciphertext_s1[93]), .B(
        ciphertext_s1[61]), .Z(new_AGEMA_signal_2105) );
  XOR2_X1 MixColumns_line3_U16_Ins_0_U1 ( .A(ciphertext_s0[28]), .B(
        MixColumns_line3_S13[5]), .Z(MixColumns_line3_n12) );
  XOR2_X1 MixColumns_line3_U16_Ins_1_U1 ( .A(ciphertext_s1[28]), .B(
        new_AGEMA_signal_2116), .Z(new_AGEMA_signal_2148) );
  XNOR2_X1 MixColumns_line3_U15_Ins0_U1 ( .A(MixColumns_line3_n10), .B(
        MixColumns_line3_n9), .ZN(MCout[4]) );
  XOR2_X1 MixColumns_line3_U15_Ins_1_U1 ( .A(new_AGEMA_signal_2821), .B(
        new_AGEMA_signal_2106), .Z(new_AGEMA_signal_2847) );
  XNOR2_X1 MixColumns_line3_U14_Ins0_U1 ( .A(ciphertext_s0[92]), .B(
        ciphertext_s0[60]), .ZN(MixColumns_line3_n9) );
  XOR2_X1 MixColumns_line3_U14_Ins_1_U1 ( .A(ciphertext_s1[92]), .B(
        ciphertext_s1[60]), .Z(new_AGEMA_signal_2106) );
  XOR2_X1 MixColumns_line3_U13_Ins_0_U1 ( .A(MixColumns_line3_S02_4_), .B(
        MixColumns_line3_S13[4]), .Z(MixColumns_line3_n10) );
  XOR2_X1 MixColumns_line3_U13_Ins_1_U1 ( .A(new_AGEMA_signal_2111), .B(
        new_AGEMA_signal_2151), .Z(new_AGEMA_signal_2821) );
  XNOR2_X1 MixColumns_line3_U12_Ins0_U1 ( .A(MixColumns_line3_n8), .B(
        MixColumns_line3_n7), .ZN(MCout[3]) );
  XOR2_X1 MixColumns_line3_U12_Ins_1_U1 ( .A(new_AGEMA_signal_2822), .B(
        new_AGEMA_signal_2107), .Z(new_AGEMA_signal_2848) );
  XNOR2_X1 MixColumns_line3_U11_Ins0_U1 ( .A(ciphertext_s0[91]), .B(
        ciphertext_s0[59]), .ZN(MixColumns_line3_n7) );
  XOR2_X1 MixColumns_line3_U11_Ins_1_U1 ( .A(ciphertext_s1[91]), .B(
        ciphertext_s1[59]), .Z(new_AGEMA_signal_2107) );
  XOR2_X1 MixColumns_line3_U10_Ins_0_U1 ( .A(MixColumns_line3_S02_3_), .B(
        MixColumns_line3_S13[3]), .Z(MixColumns_line3_n8) );
  XOR2_X1 MixColumns_line3_U10_Ins_1_U1 ( .A(new_AGEMA_signal_2112), .B(
        new_AGEMA_signal_2152), .Z(new_AGEMA_signal_2822) );
  XNOR2_X1 MixColumns_line3_U9_Ins0_U1 ( .A(MixColumns_line3_n6), .B(
        MixColumns_line3_n5), .ZN(MCout[2]) );
  XOR2_X1 MixColumns_line3_U9_Ins_1_U1 ( .A(new_AGEMA_signal_2149), .B(
        new_AGEMA_signal_2108), .Z(new_AGEMA_signal_2823) );
  XNOR2_X1 MixColumns_line3_U8_Ins0_U1 ( .A(ciphertext_s0[90]), .B(
        ciphertext_s0[58]), .ZN(MixColumns_line3_n5) );
  XOR2_X1 MixColumns_line3_U8_Ins_1_U1 ( .A(ciphertext_s1[90]), .B(
        ciphertext_s1[58]), .Z(new_AGEMA_signal_2108) );
  XOR2_X1 MixColumns_line3_U7_Ins_0_U1 ( .A(ciphertext_s0[25]), .B(
        MixColumns_line3_S13[2]), .Z(MixColumns_line3_n6) );
  XOR2_X1 MixColumns_line3_U7_Ins_1_U1 ( .A(ciphertext_s1[25]), .B(
        new_AGEMA_signal_2117), .Z(new_AGEMA_signal_2149) );
  XNOR2_X1 MixColumns_line3_U6_Ins0_U1 ( .A(MixColumns_line3_n4), .B(
        MixColumns_line3_n3), .ZN(MCout[1]) );
  XOR2_X1 MixColumns_line3_U6_Ins_1_U1 ( .A(new_AGEMA_signal_2824), .B(
        new_AGEMA_signal_2109), .Z(new_AGEMA_signal_2849) );
  XNOR2_X1 MixColumns_line3_U5_Ins0_U1 ( .A(ciphertext_s0[57]), .B(
        ciphertext_s0[89]), .ZN(MixColumns_line3_n3) );
  XOR2_X1 MixColumns_line3_U5_Ins_1_U1 ( .A(ciphertext_s1[57]), .B(
        ciphertext_s1[89]), .Z(new_AGEMA_signal_2109) );
  XOR2_X1 MixColumns_line3_U4_Ins_0_U1 ( .A(MixColumns_line3_S02_1_), .B(
        MixColumns_line3_S13[1]), .Z(MixColumns_line3_n4) );
  XOR2_X1 MixColumns_line3_U4_Ins_1_U1 ( .A(new_AGEMA_signal_2113), .B(
        new_AGEMA_signal_2153), .Z(new_AGEMA_signal_2824) );
  XNOR2_X1 MixColumns_line3_U3_Ins0_U1 ( .A(MixColumns_line3_n2), .B(
        MixColumns_line3_n1), .ZN(MCout[0]) );
  XOR2_X1 MixColumns_line3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2150), .B(
        new_AGEMA_signal_2110), .Z(new_AGEMA_signal_2825) );
  XNOR2_X1 MixColumns_line3_U2_Ins0_U1 ( .A(ciphertext_s0[56]), .B(
        ciphertext_s0[88]), .ZN(MixColumns_line3_n1) );
  XOR2_X1 MixColumns_line3_U2_Ins_1_U1 ( .A(ciphertext_s1[56]), .B(
        ciphertext_s1[88]), .Z(new_AGEMA_signal_2110) );
  XOR2_X1 MixColumns_line3_U1_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(
        MixColumns_line3_S13[0]), .Z(MixColumns_line3_n2) );
  XOR2_X1 MixColumns_line3_U1_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        new_AGEMA_signal_2118), .Z(new_AGEMA_signal_2150) );
  XOR2_X1 MixColumns_line3_timesTWO_U3_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(
        ciphertext_s0[27]), .Z(MixColumns_line3_S02_4_) );
  XOR2_X1 MixColumns_line3_timesTWO_U3_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        ciphertext_s1[27]), .Z(new_AGEMA_signal_2111) );
  XOR2_X1 MixColumns_line3_timesTWO_U2_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(
        ciphertext_s0[26]), .Z(MixColumns_line3_S02_3_) );
  XOR2_X1 MixColumns_line3_timesTWO_U2_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        ciphertext_s1[26]), .Z(new_AGEMA_signal_2112) );
  XOR2_X1 MixColumns_line3_timesTWO_U1_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(
        ciphertext_s0[24]), .Z(MixColumns_line3_S02_1_) );
  XOR2_X1 MixColumns_line3_timesTWO_U1_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        ciphertext_s1[24]), .Z(new_AGEMA_signal_2113) );
  XOR2_X1 MixColumns_line3_timesTHREE_U8_Ins_0_U1 ( .A(ciphertext_s0[127]),
        .B(ciphertext_s0[126]), .Z(MixColumns_line3_S13[7]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U8_Ins_1_U1 ( .A(ciphertext_s1[127]),
        .B(ciphertext_s1[126]), .Z(new_AGEMA_signal_2114) );
  XOR2_X1 MixColumns_line3_timesTHREE_U7_Ins_0_U1 ( .A(ciphertext_s0[126]),
        .B(ciphertext_s0[125]), .Z(MixColumns_line3_S13[6]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U7_Ins_1_U1 ( .A(ciphertext_s1[126]),
        .B(ciphertext_s1[125]), .Z(new_AGEMA_signal_2115) );
  XOR2_X1 MixColumns_line3_timesTHREE_U6_Ins_0_U1 ( .A(ciphertext_s0[125]),
        .B(ciphertext_s0[124]), .Z(MixColumns_line3_S13[5]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U6_Ins_1_U1 ( .A(ciphertext_s1[125]),
        .B(ciphertext_s1[124]), .Z(new_AGEMA_signal_2116) );
  XOR2_X1 MixColumns_line3_timesTHREE_U5_Ins_0_U1 ( .A(ciphertext_s0[124]),
        .B(MixColumns_line3_timesTHREE_input2_4_), .Z(MixColumns_line3_S13[4])
         );
  XOR2_X1 MixColumns_line3_timesTHREE_U5_Ins_1_U1 ( .A(ciphertext_s1[124]),
        .B(new_AGEMA_signal_2119), .Z(new_AGEMA_signal_2151) );
  XOR2_X1 MixColumns_line3_timesTHREE_U4_Ins_0_U1 ( .A(ciphertext_s0[123]),
        .B(MixColumns_line3_timesTHREE_input2_3_), .Z(MixColumns_line3_S13[3])
         );
  XOR2_X1 MixColumns_line3_timesTHREE_U4_Ins_1_U1 ( .A(ciphertext_s1[123]),
        .B(new_AGEMA_signal_2120), .Z(new_AGEMA_signal_2152) );
  XOR2_X1 MixColumns_line3_timesTHREE_U3_Ins_0_U1 ( .A(ciphertext_s0[122]),
        .B(ciphertext_s0[121]), .Z(MixColumns_line3_S13[2]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U3_Ins_1_U1 ( .A(ciphertext_s1[122]),
        .B(ciphertext_s1[121]), .Z(new_AGEMA_signal_2117) );
  XOR2_X1 MixColumns_line3_timesTHREE_U2_Ins_0_U1 ( .A(ciphertext_s0[121]),
        .B(MixColumns_line3_timesTHREE_input2_1_), .Z(MixColumns_line3_S13[1])
         );
  XOR2_X1 MixColumns_line3_timesTHREE_U2_Ins_1_U1 ( .A(ciphertext_s1[121]),
        .B(new_AGEMA_signal_2121), .Z(new_AGEMA_signal_2153) );
  XOR2_X1 MixColumns_line3_timesTHREE_U1_Ins_0_U1 ( .A(ciphertext_s0[120]),
        .B(ciphertext_s0[127]), .Z(MixColumns_line3_S13[0]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U1_Ins_1_U1 ( .A(ciphertext_s1[120]),
        .B(ciphertext_s1[127]), .Z(new_AGEMA_signal_2118) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U3_Ins_0_U1 ( .A(
        ciphertext_s0[127]), .B(ciphertext_s0[123]), .Z(
        MixColumns_line3_timesTHREE_input2_4_) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U3_Ins_1_U1 ( .A(
        ciphertext_s1[127]), .B(ciphertext_s1[123]), .Z(new_AGEMA_signal_2119)
         );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U2_Ins_0_U1 ( .A(
        ciphertext_s0[127]), .B(ciphertext_s0[122]), .Z(
        MixColumns_line3_timesTHREE_input2_3_) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U2_Ins_1_U1 ( .A(
        ciphertext_s1[127]), .B(ciphertext_s1[122]), .Z(new_AGEMA_signal_2120)
         );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U1_Ins_0_U1 ( .A(
        ciphertext_s0[127]), .B(ciphertext_s0[120]), .Z(
        MixColumns_line3_timesTHREE_input2_1_) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U1_Ins_1_U1 ( .A(
        ciphertext_s1[127]), .B(ciphertext_s1[120]), .Z(new_AGEMA_signal_2121)
         );
  NAND2_X1 MUX_SboxIn_mux_inst_0_U1_Ins_0_U4 ( .A1(
        MUX_SboxIn_mux_inst_0_U1_Ins_0_n8), .A2(
        MUX_SboxIn_mux_inst_0_U1_Ins_0_n7), .ZN(SboxIn[0]) );
  NAND2_X1 MUX_SboxIn_mux_inst_0_U1_Ins_0_U3 ( .A1(StateOutXORroundKey[0]),
        .A2(MUX_SboxIn_mux_inst_0_U1_Ins_0_n6), .ZN(
        MUX_SboxIn_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 MUX_SboxIn_mux_inst_0_U1_Ins_0_U2 ( .A(n190), .ZN(
        MUX_SboxIn_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_0_U1_Ins_0_U1 ( .A1(keySBIn[0]), .A2(n190),
        .ZN(MUX_SboxIn_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_0_U1_Ins_1_U4 ( .A1(
        MUX_SboxIn_mux_inst_0_U1_Ins_1_n8), .A2(
        MUX_SboxIn_mux_inst_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2826) );
  NAND2_X1 MUX_SboxIn_mux_inst_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1984),
        .A2(MUX_SboxIn_mux_inst_0_U1_Ins_1_n6), .ZN(
        MUX_SboxIn_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 MUX_SboxIn_mux_inst_0_U1_Ins_1_U2 ( .A(n190), .ZN(
        MUX_SboxIn_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2563),
        .A2(n190), .ZN(MUX_SboxIn_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_1_U1_Ins_0_U4 ( .A1(
        MUX_SboxIn_mux_inst_1_U1_Ins_0_n8), .A2(
        MUX_SboxIn_mux_inst_1_U1_Ins_0_n7), .ZN(SboxIn[1]) );
  NAND2_X1 MUX_SboxIn_mux_inst_1_U1_Ins_0_U3 ( .A1(StateOutXORroundKey[1]),
        .A2(MUX_SboxIn_mux_inst_1_U1_Ins_0_n6), .ZN(
        MUX_SboxIn_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 MUX_SboxIn_mux_inst_1_U1_Ins_0_U2 ( .A(n317), .ZN(
        MUX_SboxIn_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_1_U1_Ins_0_U1 ( .A1(keySBIn[1]), .A2(n317),
        .ZN(MUX_SboxIn_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_1_U1_Ins_1_U4 ( .A1(
        MUX_SboxIn_mux_inst_1_U1_Ins_1_n8), .A2(
        MUX_SboxIn_mux_inst_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2827) );
  NAND2_X1 MUX_SboxIn_mux_inst_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1987),
        .A2(MUX_SboxIn_mux_inst_1_U1_Ins_1_n6), .ZN(
        MUX_SboxIn_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 MUX_SboxIn_mux_inst_1_U1_Ins_1_U2 ( .A(n317), .ZN(
        MUX_SboxIn_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2566),
        .A2(n317), .ZN(MUX_SboxIn_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_2_U1_Ins_0_U4 ( .A1(
        MUX_SboxIn_mux_inst_2_U1_Ins_0_n8), .A2(
        MUX_SboxIn_mux_inst_2_U1_Ins_0_n7), .ZN(SboxIn[2]) );
  NAND2_X1 MUX_SboxIn_mux_inst_2_U1_Ins_0_U3 ( .A1(StateOutXORroundKey[2]),
        .A2(MUX_SboxIn_mux_inst_2_U1_Ins_0_n6), .ZN(
        MUX_SboxIn_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 MUX_SboxIn_mux_inst_2_U1_Ins_0_U2 ( .A(n318), .ZN(
        MUX_SboxIn_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_2_U1_Ins_0_U1 ( .A1(keySBIn[2]), .A2(n318),
        .ZN(MUX_SboxIn_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_2_U1_Ins_1_U4 ( .A1(
        MUX_SboxIn_mux_inst_2_U1_Ins_1_n8), .A2(
        MUX_SboxIn_mux_inst_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2828) );
  NAND2_X1 MUX_SboxIn_mux_inst_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1990),
        .A2(MUX_SboxIn_mux_inst_2_U1_Ins_1_n6), .ZN(
        MUX_SboxIn_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 MUX_SboxIn_mux_inst_2_U1_Ins_1_U2 ( .A(n318), .ZN(
        MUX_SboxIn_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2569),
        .A2(n318), .ZN(MUX_SboxIn_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_3_U1_Ins_0_U4 ( .A1(
        MUX_SboxIn_mux_inst_3_U1_Ins_0_n8), .A2(
        MUX_SboxIn_mux_inst_3_U1_Ins_0_n7), .ZN(SboxIn[3]) );
  NAND2_X1 MUX_SboxIn_mux_inst_3_U1_Ins_0_U3 ( .A1(StateOutXORroundKey[3]),
        .A2(MUX_SboxIn_mux_inst_3_U1_Ins_0_n6), .ZN(
        MUX_SboxIn_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 MUX_SboxIn_mux_inst_3_U1_Ins_0_U2 ( .A(n314), .ZN(
        MUX_SboxIn_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_3_U1_Ins_0_U1 ( .A1(keySBIn[3]), .A2(n314),
        .ZN(MUX_SboxIn_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_3_U1_Ins_1_U4 ( .A1(
        MUX_SboxIn_mux_inst_3_U1_Ins_1_n8), .A2(
        MUX_SboxIn_mux_inst_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2829) );
  NAND2_X1 MUX_SboxIn_mux_inst_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1993),
        .A2(MUX_SboxIn_mux_inst_3_U1_Ins_1_n6), .ZN(
        MUX_SboxIn_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 MUX_SboxIn_mux_inst_3_U1_Ins_1_U2 ( .A(n314), .ZN(
        MUX_SboxIn_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2572),
        .A2(n314), .ZN(MUX_SboxIn_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_4_U1_Ins_0_U4 ( .A1(
        MUX_SboxIn_mux_inst_4_U1_Ins_0_n8), .A2(
        MUX_SboxIn_mux_inst_4_U1_Ins_0_n7), .ZN(SboxIn[4]) );
  NAND2_X1 MUX_SboxIn_mux_inst_4_U1_Ins_0_U3 ( .A1(StateOutXORroundKey[4]),
        .A2(MUX_SboxIn_mux_inst_4_U1_Ins_0_n6), .ZN(
        MUX_SboxIn_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 MUX_SboxIn_mux_inst_4_U1_Ins_0_U2 ( .A(n315), .ZN(
        MUX_SboxIn_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_4_U1_Ins_0_U1 ( .A1(keySBIn[4]), .A2(n315),
        .ZN(MUX_SboxIn_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_4_U1_Ins_1_U4 ( .A1(
        MUX_SboxIn_mux_inst_4_U1_Ins_1_n8), .A2(
        MUX_SboxIn_mux_inst_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2830) );
  NAND2_X1 MUX_SboxIn_mux_inst_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1996),
        .A2(MUX_SboxIn_mux_inst_4_U1_Ins_1_n6), .ZN(
        MUX_SboxIn_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 MUX_SboxIn_mux_inst_4_U1_Ins_1_U2 ( .A(n315), .ZN(
        MUX_SboxIn_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2575),
        .A2(n315), .ZN(MUX_SboxIn_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_5_U1_Ins_0_U4 ( .A1(
        MUX_SboxIn_mux_inst_5_U1_Ins_0_n8), .A2(
        MUX_SboxIn_mux_inst_5_U1_Ins_0_n7), .ZN(SboxIn[5]) );
  NAND2_X1 MUX_SboxIn_mux_inst_5_U1_Ins_0_U3 ( .A1(StateOutXORroundKey[5]),
        .A2(MUX_SboxIn_mux_inst_5_U1_Ins_0_n6), .ZN(
        MUX_SboxIn_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 MUX_SboxIn_mux_inst_5_U1_Ins_0_U2 ( .A(n316), .ZN(
        MUX_SboxIn_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_5_U1_Ins_0_U1 ( .A1(keySBIn[5]), .A2(n316),
        .ZN(MUX_SboxIn_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_5_U1_Ins_1_U4 ( .A1(
        MUX_SboxIn_mux_inst_5_U1_Ins_1_n8), .A2(
        MUX_SboxIn_mux_inst_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2831) );
  NAND2_X1 MUX_SboxIn_mux_inst_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_1999),
        .A2(MUX_SboxIn_mux_inst_5_U1_Ins_1_n6), .ZN(
        MUX_SboxIn_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 MUX_SboxIn_mux_inst_5_U1_Ins_1_U2 ( .A(n316), .ZN(
        MUX_SboxIn_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2578),
        .A2(n316), .ZN(MUX_SboxIn_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_6_U1_Ins_0_U4 ( .A1(
        MUX_SboxIn_mux_inst_6_U1_Ins_0_n8), .A2(
        MUX_SboxIn_mux_inst_6_U1_Ins_0_n7), .ZN(SboxIn[6]) );
  NAND2_X1 MUX_SboxIn_mux_inst_6_U1_Ins_0_U3 ( .A1(StateOutXORroundKey[6]),
        .A2(MUX_SboxIn_mux_inst_6_U1_Ins_0_n6), .ZN(
        MUX_SboxIn_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 MUX_SboxIn_mux_inst_6_U1_Ins_0_U2 ( .A(n319), .ZN(
        MUX_SboxIn_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_6_U1_Ins_0_U1 ( .A1(keySBIn[6]), .A2(n319),
        .ZN(MUX_SboxIn_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_6_U1_Ins_1_U4 ( .A1(
        MUX_SboxIn_mux_inst_6_U1_Ins_1_n8), .A2(
        MUX_SboxIn_mux_inst_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2832) );
  NAND2_X1 MUX_SboxIn_mux_inst_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2002),
        .A2(MUX_SboxIn_mux_inst_6_U1_Ins_1_n6), .ZN(
        MUX_SboxIn_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 MUX_SboxIn_mux_inst_6_U1_Ins_1_U2 ( .A(n319), .ZN(
        MUX_SboxIn_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2581),
        .A2(n319), .ZN(MUX_SboxIn_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_7_U1_Ins_0_U4 ( .A1(
        MUX_SboxIn_mux_inst_7_U1_Ins_0_n8), .A2(
        MUX_SboxIn_mux_inst_7_U1_Ins_0_n7), .ZN(SboxIn[7]) );
  NAND2_X1 MUX_SboxIn_mux_inst_7_U1_Ins_0_U3 ( .A1(StateOutXORroundKey[7]),
        .A2(MUX_SboxIn_mux_inst_7_U1_Ins_0_n6), .ZN(
        MUX_SboxIn_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 MUX_SboxIn_mux_inst_7_U1_Ins_0_U2 ( .A(n315), .ZN(
        MUX_SboxIn_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_7_U1_Ins_0_U1 ( .A1(keySBIn[7]), .A2(n315),
        .ZN(MUX_SboxIn_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 MUX_SboxIn_mux_inst_7_U1_Ins_1_U4 ( .A1(
        MUX_SboxIn_mux_inst_7_U1_Ins_1_n8), .A2(
        MUX_SboxIn_mux_inst_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_2833) );
  NAND2_X1 MUX_SboxIn_mux_inst_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_2005),
        .A2(MUX_SboxIn_mux_inst_7_U1_Ins_1_n6), .ZN(
        MUX_SboxIn_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 MUX_SboxIn_mux_inst_7_U1_Ins_1_U2 ( .A(n315), .ZN(
        MUX_SboxIn_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 MUX_SboxIn_mux_inst_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_2584),
        .A2(n315), .ZN(MUX_SboxIn_mux_inst_7_U1_Ins_1_n8) );
  XOR2_X1 Inst_bSbox_XOR_T1_U1_Ins_0_U1 ( .A(SboxIn[7]), .B(SboxIn[4]), .Z(
        Inst_bSbox_T1) );
  XOR2_X1 Inst_bSbox_XOR_T1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2833), .B(
        new_AGEMA_signal_2830), .Z(new_AGEMA_signal_2850) );
  XOR2_X1 Inst_bSbox_XOR_T2_U1_Ins_0_U1 ( .A(SboxIn[7]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T2) );
  XOR2_X1 Inst_bSbox_XOR_T2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2833), .B(
        new_AGEMA_signal_2828), .Z(new_AGEMA_signal_2851) );
  XOR2_X1 Inst_bSbox_XOR_T3_U1_Ins_0_U1 ( .A(SboxIn[7]), .B(SboxIn[1]), .Z(
        Inst_bSbox_T3) );
  XOR2_X1 Inst_bSbox_XOR_T3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2833), .B(
        new_AGEMA_signal_2827), .Z(new_AGEMA_signal_2852) );
  XOR2_X1 Inst_bSbox_XOR_T4_U1_Ins_0_U1 ( .A(SboxIn[4]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T4) );
  XOR2_X1 Inst_bSbox_XOR_T4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2830), .B(
        new_AGEMA_signal_2828), .Z(new_AGEMA_signal_2853) );
  XOR2_X1 Inst_bSbox_XOR_T5_U1_Ins_0_U1 ( .A(SboxIn[3]), .B(SboxIn[1]), .Z(
        Inst_bSbox_T5) );
  XOR2_X1 Inst_bSbox_XOR_T5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2829), .B(
        new_AGEMA_signal_2827), .Z(new_AGEMA_signal_2854) );
  XOR2_X1 Inst_bSbox_XOR_T6_U1_Ins_0_U1 ( .A(Inst_bSbox_T1), .B(Inst_bSbox_T5),
        .Z(Inst_bSbox_T6) );
  XOR2_X1 Inst_bSbox_XOR_T6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2850), .B(
        new_AGEMA_signal_2854), .Z(new_AGEMA_signal_3000) );
  XOR2_X1 Inst_bSbox_XOR_T7_U1_Ins_0_U1 ( .A(SboxIn[6]), .B(SboxIn[5]), .Z(
        Inst_bSbox_T7) );
  XOR2_X1 Inst_bSbox_XOR_T7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2832), .B(
        new_AGEMA_signal_2831), .Z(new_AGEMA_signal_2855) );
  XOR2_X1 Inst_bSbox_XOR_T8_U1_Ins_0_U1 ( .A(SboxIn[0]), .B(Inst_bSbox_T6),
        .Z(Inst_bSbox_T8) );
  XOR2_X1 Inst_bSbox_XOR_T8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2826), .B(
        new_AGEMA_signal_3000), .Z(new_AGEMA_signal_3032) );
  XOR2_X1 Inst_bSbox_XOR_T9_U1_Ins_0_U1 ( .A(SboxIn[0]), .B(Inst_bSbox_T7),
        .Z(Inst_bSbox_T9) );
  XOR2_X1 Inst_bSbox_XOR_T9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2826), .B(
        new_AGEMA_signal_2855), .Z(new_AGEMA_signal_3001) );
  XOR2_X1 Inst_bSbox_XOR_T10_U1_Ins_0_U1 ( .A(Inst_bSbox_T6), .B(Inst_bSbox_T7), .Z(Inst_bSbox_T10) );
  XOR2_X1 Inst_bSbox_XOR_T10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3000), .B(
        new_AGEMA_signal_2855), .Z(new_AGEMA_signal_3033) );
  XOR2_X1 Inst_bSbox_XOR_T11_U1_Ins_0_U1 ( .A(SboxIn[6]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T11) );
  XOR2_X1 Inst_bSbox_XOR_T11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2832), .B(
        new_AGEMA_signal_2828), .Z(new_AGEMA_signal_2856) );
  XOR2_X1 Inst_bSbox_XOR_T12_U1_Ins_0_U1 ( .A(SboxIn[5]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T12) );
  XOR2_X1 Inst_bSbox_XOR_T12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2831), .B(
        new_AGEMA_signal_2828), .Z(new_AGEMA_signal_2857) );
  XOR2_X1 Inst_bSbox_XOR_T13_U1_Ins_0_U1 ( .A(Inst_bSbox_T3), .B(Inst_bSbox_T4), .Z(Inst_bSbox_T13) );
  XOR2_X1 Inst_bSbox_XOR_T13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2852), .B(
        new_AGEMA_signal_2853), .Z(new_AGEMA_signal_3002) );
  XOR2_X1 Inst_bSbox_XOR_T14_U1_Ins_0_U1 ( .A(Inst_bSbox_T6), .B(
        Inst_bSbox_T11), .Z(Inst_bSbox_T14) );
  XOR2_X1 Inst_bSbox_XOR_T14_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3000), .B(
        new_AGEMA_signal_2856), .Z(new_AGEMA_signal_3034) );
  XOR2_X1 Inst_bSbox_XOR_T15_U1_Ins_0_U1 ( .A(Inst_bSbox_T5), .B(
        Inst_bSbox_T11), .Z(Inst_bSbox_T15) );
  XOR2_X1 Inst_bSbox_XOR_T15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2854), .B(
        new_AGEMA_signal_2856), .Z(new_AGEMA_signal_3003) );
  XOR2_X1 Inst_bSbox_XOR_T16_U1_Ins_0_U1 ( .A(Inst_bSbox_T5), .B(
        Inst_bSbox_T12), .Z(Inst_bSbox_T16) );
  XOR2_X1 Inst_bSbox_XOR_T16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2854), .B(
        new_AGEMA_signal_2857), .Z(new_AGEMA_signal_3004) );
  XOR2_X1 Inst_bSbox_XOR_T17_U1_Ins_0_U1 ( .A(Inst_bSbox_T9), .B(
        Inst_bSbox_T16), .Z(Inst_bSbox_T17) );
  XOR2_X1 Inst_bSbox_XOR_T17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3001), .B(
        new_AGEMA_signal_3004), .Z(new_AGEMA_signal_3035) );
  XOR2_X1 Inst_bSbox_XOR_T18_U1_Ins_0_U1 ( .A(SboxIn[4]), .B(SboxIn[0]), .Z(
        Inst_bSbox_T18) );
  XOR2_X1 Inst_bSbox_XOR_T18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2830), .B(
        new_AGEMA_signal_2826), .Z(new_AGEMA_signal_2858) );
  XOR2_X1 Inst_bSbox_XOR_T19_U1_Ins_0_U1 ( .A(Inst_bSbox_T7), .B(
        Inst_bSbox_T18), .Z(Inst_bSbox_T19) );
  XOR2_X1 Inst_bSbox_XOR_T19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2855), .B(
        new_AGEMA_signal_2858), .Z(new_AGEMA_signal_3005) );
  XOR2_X1 Inst_bSbox_XOR_T20_U1_Ins_0_U1 ( .A(Inst_bSbox_T1), .B(
        Inst_bSbox_T19), .Z(Inst_bSbox_T20) );
  XOR2_X1 Inst_bSbox_XOR_T20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2850), .B(
        new_AGEMA_signal_3005), .Z(new_AGEMA_signal_3036) );
  XOR2_X1 Inst_bSbox_XOR_T21_U1_Ins_0_U1 ( .A(SboxIn[1]), .B(SboxIn[0]), .Z(
        Inst_bSbox_T21) );
  XOR2_X1 Inst_bSbox_XOR_T21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2827), .B(
        new_AGEMA_signal_2826), .Z(new_AGEMA_signal_2859) );
  XOR2_X1 Inst_bSbox_XOR_T22_U1_Ins_0_U1 ( .A(Inst_bSbox_T7), .B(
        Inst_bSbox_T21), .Z(Inst_bSbox_T22) );
  XOR2_X1 Inst_bSbox_XOR_T22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2855), .B(
        new_AGEMA_signal_2859), .Z(new_AGEMA_signal_3006) );
  XOR2_X1 Inst_bSbox_XOR_T23_U1_Ins_0_U1 ( .A(Inst_bSbox_T2), .B(
        Inst_bSbox_T22), .Z(Inst_bSbox_T23) );
  XOR2_X1 Inst_bSbox_XOR_T23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2851), .B(
        new_AGEMA_signal_3006), .Z(new_AGEMA_signal_3037) );
  XOR2_X1 Inst_bSbox_XOR_T24_U1_Ins_0_U1 ( .A(Inst_bSbox_T2), .B(
        Inst_bSbox_T10), .Z(Inst_bSbox_T24) );
  XOR2_X1 Inst_bSbox_XOR_T24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2851), .B(
        new_AGEMA_signal_3033), .Z(new_AGEMA_signal_3117) );
  XOR2_X1 Inst_bSbox_XOR_T25_U1_Ins_0_U1 ( .A(Inst_bSbox_T20), .B(
        Inst_bSbox_T17), .Z(Inst_bSbox_T25) );
  XOR2_X1 Inst_bSbox_XOR_T25_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3036), .B(
        new_AGEMA_signal_3035), .Z(new_AGEMA_signal_3118) );
  XOR2_X1 Inst_bSbox_XOR_T26_U1_Ins_0_U1 ( .A(Inst_bSbox_T3), .B(
        Inst_bSbox_T16), .Z(Inst_bSbox_T26) );
  XOR2_X1 Inst_bSbox_XOR_T26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2852), .B(
        new_AGEMA_signal_3004), .Z(new_AGEMA_signal_3038) );
  XOR2_X1 Inst_bSbox_XOR_T27_U1_Ins_0_U1 ( .A(Inst_bSbox_T1), .B(
        Inst_bSbox_T12), .Z(Inst_bSbox_T27) );
  XOR2_X1 Inst_bSbox_XOR_T27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2850), .B(
        new_AGEMA_signal_2857), .Z(new_AGEMA_signal_3007) );
  XOR2_X1 Inst_bSbox_AND_M1_U1_U16 ( .A(Fresh[0]), .B(Inst_bSbox_AND_M1_U1_n7),
        .Z(Inst_bSbox_AND_M1_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M1_U1_U15 ( .A1(new_AGEMA_signal_3002), .A2(
        Inst_bSbox_AND_M1_U1_n6), .ZN(Inst_bSbox_AND_M1_U1_n7) );
  XOR2_X1 Inst_bSbox_AND_M1_U1_U14 ( .A(Fresh[0]), .B(Inst_bSbox_AND_M1_U1_n5),
        .Z(Inst_bSbox_AND_M1_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M1_U1_U13 ( .A1(Inst_bSbox_T13), .A2(
        Inst_bSbox_AND_M1_U1_n6), .ZN(Inst_bSbox_AND_M1_U1_n5) );
  XNOR2_X1 Inst_bSbox_AND_M1_U1_U12 ( .A(Inst_bSbox_AND_M1_U1_n4), .B(
        Inst_bSbox_AND_M1_U1_n3), .ZN(Inst_bSbox_M1) );
  NAND2_X1 Inst_bSbox_AND_M1_U1_U11 ( .A1(Inst_bSbox_AND_M1_U1_a_reg[0]), .A2(
        Inst_bSbox_AND_M1_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M1_U1_n3) );
  XOR2_X1 Inst_bSbox_AND_M1_U1_U10 ( .A(Inst_bSbox_AND_M1_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M1_U1_z[0]), .Z(Inst_bSbox_AND_M1_U1_n4) );
  XNOR2_X1 Inst_bSbox_AND_M1_U1_U9 ( .A(Inst_bSbox_AND_M1_U1_n2), .B(
        Inst_bSbox_AND_M1_U1_n1), .ZN(new_AGEMA_signal_3039) );
  NAND2_X1 Inst_bSbox_AND_M1_U1_U8 ( .A1(Inst_bSbox_AND_M1_U1_a_reg[1]), .A2(
        Inst_bSbox_AND_M1_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M1_U1_n1) );
  XOR2_X1 Inst_bSbox_AND_M1_U1_U7 ( .A(Inst_bSbox_AND_M1_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M1_U1_z[1]), .Z(Inst_bSbox_AND_M1_U1_n2) );
  XNOR2_X1 Inst_bSbox_AND_M1_U1_U6 ( .A(new_AGEMA_signal_3000), .B(
        Inst_bSbox_AND_M1_U1_n6), .ZN(Inst_bSbox_AND_M1_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M1_U1_U5 ( .A(Inst_bSbox_T6), .B(
        Inst_bSbox_AND_M1_U1_n6), .ZN(Inst_bSbox_AND_M1_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M1_U1_U4 ( .A(Fresh[1]), .ZN(Inst_bSbox_AND_M1_U1_n6)
         );
  AND2_X1 Inst_bSbox_AND_M1_U1_U3 ( .A1(Inst_bSbox_T13), .A2(Inst_bSbox_T6),
        .ZN(Inst_bSbox_AND_M1_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M1_U1_U2 ( .A1(new_AGEMA_signal_3002), .A2(
        new_AGEMA_signal_3000), .ZN(Inst_bSbox_AND_M1_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M1_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M1_U1_z[0])
         );
  DFF_X1 Inst_bSbox_AND_M1_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_T13),
        .CK(clk), .Q(Inst_bSbox_AND_M1_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M1_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M1_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M1_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M1_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M1_U1_z[1])
         );
  DFF_X1 Inst_bSbox_AND_M1_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3002), .CK(clk), .Q(Inst_bSbox_AND_M1_U1_a_reg[1]) );
  DFF_X1 Inst_bSbox_AND_M1_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M1_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M1_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M2_U1_U16 ( .A(Fresh[2]), .B(Inst_bSbox_AND_M2_U1_n23), .Z(Inst_bSbox_AND_M2_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M2_U1_U15 ( .A1(new_AGEMA_signal_3037), .A2(
        Inst_bSbox_AND_M2_U1_n22), .ZN(Inst_bSbox_AND_M2_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M2_U1_U14 ( .A(Fresh[2]), .B(Inst_bSbox_AND_M2_U1_n21), .Z(Inst_bSbox_AND_M2_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M2_U1_U13 ( .A1(Inst_bSbox_T23), .A2(
        Inst_bSbox_AND_M2_U1_n22), .ZN(Inst_bSbox_AND_M2_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M2_U1_U12 ( .A(Inst_bSbox_AND_M2_U1_n20), .B(
        Inst_bSbox_AND_M2_U1_n19), .ZN(Inst_bSbox_M2) );
  NAND2_X1 Inst_bSbox_AND_M2_U1_U11 ( .A1(Inst_bSbox_AND_M2_U1_a_reg[0]), .A2(
        Inst_bSbox_AND_M2_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M2_U1_n19) );
  XOR2_X1 Inst_bSbox_AND_M2_U1_U10 ( .A(Inst_bSbox_AND_M2_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M2_U1_z[0]), .Z(Inst_bSbox_AND_M2_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M2_U1_U9 ( .A(Inst_bSbox_AND_M2_U1_n18), .B(
        Inst_bSbox_AND_M2_U1_n17), .ZN(new_AGEMA_signal_3119) );
  NAND2_X1 Inst_bSbox_AND_M2_U1_U8 ( .A1(Inst_bSbox_AND_M2_U1_a_reg[1]), .A2(
        Inst_bSbox_AND_M2_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M2_U1_n17) );
  XOR2_X1 Inst_bSbox_AND_M2_U1_U7 ( .A(Inst_bSbox_AND_M2_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M2_U1_z[1]), .Z(Inst_bSbox_AND_M2_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M2_U1_U6 ( .A(new_AGEMA_signal_3032), .B(
        Inst_bSbox_AND_M2_U1_n22), .ZN(Inst_bSbox_AND_M2_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M2_U1_U5 ( .A(Inst_bSbox_T8), .B(
        Inst_bSbox_AND_M2_U1_n22), .ZN(Inst_bSbox_AND_M2_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M2_U1_U4 ( .A(Fresh[3]), .ZN(Inst_bSbox_AND_M2_U1_n22)
         );
  AND2_X1 Inst_bSbox_AND_M2_U1_U3 ( .A1(Inst_bSbox_T23), .A2(Inst_bSbox_T8),
        .ZN(Inst_bSbox_AND_M2_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M2_U1_U2 ( .A1(new_AGEMA_signal_3037), .A2(
        new_AGEMA_signal_3032), .ZN(Inst_bSbox_AND_M2_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M2_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M2_U1_z[0])
         );
  DFF_X1 Inst_bSbox_AND_M2_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_T23),
        .CK(clk), .Q(Inst_bSbox_AND_M2_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M2_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M2_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M2_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M2_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M2_U1_z[1])
         );
  DFF_X1 Inst_bSbox_AND_M2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3037), .CK(clk), .Q(Inst_bSbox_AND_M2_U1_a_reg[1]) );
  DFF_X1 Inst_bSbox_AND_M2_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M2_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M2_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_M3_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3602), .B(
        Inst_bSbox_M1), .Z(Inst_bSbox_M3) );
  XOR2_X1 Inst_bSbox_XOR_M3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3603), .B(
        new_AGEMA_signal_3039), .Z(new_AGEMA_signal_3120) );
  XOR2_X1 Inst_bSbox_AND_M4_U1_U16 ( .A(Fresh[4]), .B(Inst_bSbox_AND_M4_U1_n23), .Z(Inst_bSbox_AND_M4_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M4_U1_U15 ( .A1(new_AGEMA_signal_3005), .A2(
        Inst_bSbox_AND_M4_U1_n22), .ZN(Inst_bSbox_AND_M4_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M4_U1_U14 ( .A(Fresh[4]), .B(Inst_bSbox_AND_M4_U1_n21), .Z(Inst_bSbox_AND_M4_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M4_U1_U13 ( .A1(Inst_bSbox_T19), .A2(
        Inst_bSbox_AND_M4_U1_n22), .ZN(Inst_bSbox_AND_M4_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M4_U1_U12 ( .A(Inst_bSbox_AND_M4_U1_n20), .B(
        Inst_bSbox_AND_M4_U1_n19), .ZN(Inst_bSbox_M4) );
  NAND2_X1 Inst_bSbox_AND_M4_U1_U11 ( .A1(Inst_bSbox_AND_M4_U1_a_reg[0]), .A2(
        Inst_bSbox_AND_M4_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M4_U1_n19) );
  XOR2_X1 Inst_bSbox_AND_M4_U1_U10 ( .A(Inst_bSbox_AND_M4_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M4_U1_z[0]), .Z(Inst_bSbox_AND_M4_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M4_U1_U9 ( .A(Inst_bSbox_AND_M4_U1_n18), .B(
        Inst_bSbox_AND_M4_U1_n17), .ZN(new_AGEMA_signal_3040) );
  NAND2_X1 Inst_bSbox_AND_M4_U1_U8 ( .A1(Inst_bSbox_AND_M4_U1_a_reg[1]), .A2(
        Inst_bSbox_AND_M4_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M4_U1_n17) );
  XOR2_X1 Inst_bSbox_AND_M4_U1_U7 ( .A(Inst_bSbox_AND_M4_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M4_U1_z[1]), .Z(Inst_bSbox_AND_M4_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M4_U1_U6 ( .A(new_AGEMA_signal_2826), .B(
        Inst_bSbox_AND_M4_U1_n22), .ZN(Inst_bSbox_AND_M4_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M4_U1_U5 ( .A(SboxIn[0]), .B(
        Inst_bSbox_AND_M4_U1_n22), .ZN(Inst_bSbox_AND_M4_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M4_U1_U4 ( .A(Fresh[5]), .ZN(Inst_bSbox_AND_M4_U1_n22)
         );
  AND2_X1 Inst_bSbox_AND_M4_U1_U3 ( .A1(new_AGEMA_signal_3005), .A2(
        new_AGEMA_signal_2826), .ZN(Inst_bSbox_AND_M4_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M4_U1_U2 ( .A1(Inst_bSbox_T19), .A2(SboxIn[0]), .ZN(
        Inst_bSbox_AND_M4_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M4_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M4_U1_z[0])
         );
  DFF_X1 Inst_bSbox_AND_M4_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_T19),
        .CK(clk), .Q(Inst_bSbox_AND_M4_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M4_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M4_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M4_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M4_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M4_U1_z[1])
         );
  DFF_X1 Inst_bSbox_AND_M4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3005), .CK(clk), .Q(Inst_bSbox_AND_M4_U1_a_reg[1]) );
  DFF_X1 Inst_bSbox_AND_M4_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M4_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M4_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_M5_U1_Ins_0_U1 ( .A(Inst_bSbox_M4), .B(Inst_bSbox_M1),
        .Z(Inst_bSbox_M5) );
  XOR2_X1 Inst_bSbox_XOR_M5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3040), .B(
        new_AGEMA_signal_3039), .Z(new_AGEMA_signal_3121) );
  XOR2_X1 Inst_bSbox_AND_M6_U1_U16 ( .A(Fresh[6]), .B(Inst_bSbox_AND_M6_U1_n23), .Z(Inst_bSbox_AND_M6_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M6_U1_U15 ( .A1(new_AGEMA_signal_2852), .A2(
        Inst_bSbox_AND_M6_U1_n22), .ZN(Inst_bSbox_AND_M6_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M6_U1_U14 ( .A(Fresh[6]), .B(Inst_bSbox_AND_M6_U1_n21), .Z(Inst_bSbox_AND_M6_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M6_U1_U13 ( .A1(Inst_bSbox_T3), .A2(
        Inst_bSbox_AND_M6_U1_n22), .ZN(Inst_bSbox_AND_M6_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M6_U1_U12 ( .A(Inst_bSbox_AND_M6_U1_n20), .B(
        Inst_bSbox_AND_M6_U1_n19), .ZN(Inst_bSbox_M6) );
  NAND2_X1 Inst_bSbox_AND_M6_U1_U11 ( .A1(Inst_bSbox_AND_M6_U1_a_reg[0]), .A2(
        Inst_bSbox_AND_M6_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M6_U1_n19) );
  XOR2_X1 Inst_bSbox_AND_M6_U1_U10 ( .A(Inst_bSbox_AND_M6_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M6_U1_z[0]), .Z(Inst_bSbox_AND_M6_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M6_U1_U9 ( .A(Inst_bSbox_AND_M6_U1_n18), .B(
        Inst_bSbox_AND_M6_U1_n17), .ZN(new_AGEMA_signal_3041) );
  NAND2_X1 Inst_bSbox_AND_M6_U1_U8 ( .A1(Inst_bSbox_AND_M6_U1_a_reg[1]), .A2(
        Inst_bSbox_AND_M6_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M6_U1_n17) );
  XOR2_X1 Inst_bSbox_AND_M6_U1_U7 ( .A(Inst_bSbox_AND_M6_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M6_U1_z[1]), .Z(Inst_bSbox_AND_M6_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M6_U1_U6 ( .A(new_AGEMA_signal_3004), .B(
        Inst_bSbox_AND_M6_U1_n22), .ZN(Inst_bSbox_AND_M6_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M6_U1_U5 ( .A(Inst_bSbox_T16), .B(
        Inst_bSbox_AND_M6_U1_n22), .ZN(Inst_bSbox_AND_M6_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M6_U1_U4 ( .A(Fresh[7]), .ZN(Inst_bSbox_AND_M6_U1_n22)
         );
  AND2_X1 Inst_bSbox_AND_M6_U1_U3 ( .A1(new_AGEMA_signal_2852), .A2(
        new_AGEMA_signal_3004), .ZN(Inst_bSbox_AND_M6_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M6_U1_U2 ( .A1(Inst_bSbox_T3), .A2(Inst_bSbox_T16),
        .ZN(Inst_bSbox_AND_M6_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M6_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M6_U1_z[0])
         );
  DFF_X1 Inst_bSbox_AND_M6_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_T3),
        .CK(clk), .Q(Inst_bSbox_AND_M6_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M6_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M6_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M6_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M6_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M6_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M6_U1_z[1])
         );
  DFF_X1 Inst_bSbox_AND_M6_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2852), .CK(clk), .Q(Inst_bSbox_AND_M6_U1_a_reg[1]) );
  DFF_X1 Inst_bSbox_AND_M6_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M6_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M6_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M6_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M7_U1_U16 ( .A(Fresh[8]), .B(Inst_bSbox_AND_M7_U1_n23), .Z(Inst_bSbox_AND_M7_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M7_U1_U15 ( .A1(new_AGEMA_signal_3006), .A2(
        Inst_bSbox_AND_M7_U1_n22), .ZN(Inst_bSbox_AND_M7_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M7_U1_U14 ( .A(Fresh[8]), .B(Inst_bSbox_AND_M7_U1_n21), .Z(Inst_bSbox_AND_M7_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M7_U1_U13 ( .A1(Inst_bSbox_T22), .A2(
        Inst_bSbox_AND_M7_U1_n22), .ZN(Inst_bSbox_AND_M7_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M7_U1_U12 ( .A(Inst_bSbox_AND_M7_U1_n20), .B(
        Inst_bSbox_AND_M7_U1_n19), .ZN(Inst_bSbox_M7) );
  NAND2_X1 Inst_bSbox_AND_M7_U1_U11 ( .A1(Inst_bSbox_AND_M7_U1_a_reg[0]), .A2(
        Inst_bSbox_AND_M7_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M7_U1_n19) );
  XOR2_X1 Inst_bSbox_AND_M7_U1_U10 ( .A(Inst_bSbox_AND_M7_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M7_U1_z[0]), .Z(Inst_bSbox_AND_M7_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M7_U1_U9 ( .A(Inst_bSbox_AND_M7_U1_n18), .B(
        Inst_bSbox_AND_M7_U1_n17), .ZN(new_AGEMA_signal_3042) );
  NAND2_X1 Inst_bSbox_AND_M7_U1_U8 ( .A1(Inst_bSbox_AND_M7_U1_a_reg[1]), .A2(
        Inst_bSbox_AND_M7_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M7_U1_n17) );
  XOR2_X1 Inst_bSbox_AND_M7_U1_U7 ( .A(Inst_bSbox_AND_M7_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M7_U1_z[1]), .Z(Inst_bSbox_AND_M7_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M7_U1_U6 ( .A(new_AGEMA_signal_3001), .B(
        Inst_bSbox_AND_M7_U1_n22), .ZN(Inst_bSbox_AND_M7_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M7_U1_U5 ( .A(Inst_bSbox_T9), .B(
        Inst_bSbox_AND_M7_U1_n22), .ZN(Inst_bSbox_AND_M7_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M7_U1_U4 ( .A(Fresh[9]), .ZN(Inst_bSbox_AND_M7_U1_n22)
         );
  AND2_X1 Inst_bSbox_AND_M7_U1_U3 ( .A1(Inst_bSbox_T22), .A2(Inst_bSbox_T9),
        .ZN(Inst_bSbox_AND_M7_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M7_U1_U2 ( .A1(new_AGEMA_signal_3006), .A2(
        new_AGEMA_signal_3001), .ZN(Inst_bSbox_AND_M7_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M7_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M7_U1_z[0])
         );
  DFF_X1 Inst_bSbox_AND_M7_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_T22),
        .CK(clk), .Q(Inst_bSbox_AND_M7_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M7_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M7_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M7_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M7_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M7_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M7_U1_z[1])
         );
  DFF_X1 Inst_bSbox_AND_M7_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3006), .CK(clk), .Q(Inst_bSbox_AND_M7_U1_a_reg[1]) );
  DFF_X1 Inst_bSbox_AND_M7_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M7_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M7_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M7_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_M8_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3604), .B(
        Inst_bSbox_M6), .Z(Inst_bSbox_M8) );
  XOR2_X1 Inst_bSbox_XOR_M8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3605), .B(
        new_AGEMA_signal_3041), .Z(new_AGEMA_signal_3122) );
  XOR2_X1 Inst_bSbox_AND_M9_U1_U16 ( .A(Fresh[10]), .B(
        Inst_bSbox_AND_M9_U1_n23), .Z(Inst_bSbox_AND_M9_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M9_U1_U15 ( .A1(new_AGEMA_signal_3036), .A2(
        Inst_bSbox_AND_M9_U1_n22), .ZN(Inst_bSbox_AND_M9_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M9_U1_U14 ( .A(Fresh[10]), .B(
        Inst_bSbox_AND_M9_U1_n21), .Z(Inst_bSbox_AND_M9_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M9_U1_U13 ( .A1(Inst_bSbox_T20), .A2(
        Inst_bSbox_AND_M9_U1_n22), .ZN(Inst_bSbox_AND_M9_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M9_U1_U12 ( .A(Inst_bSbox_AND_M9_U1_n20), .B(
        Inst_bSbox_AND_M9_U1_n19), .ZN(Inst_bSbox_M9) );
  NAND2_X1 Inst_bSbox_AND_M9_U1_U11 ( .A1(Inst_bSbox_AND_M9_U1_a_reg[0]), .A2(
        Inst_bSbox_AND_M9_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M9_U1_n19) );
  XOR2_X1 Inst_bSbox_AND_M9_U1_U10 ( .A(Inst_bSbox_AND_M9_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M9_U1_z[0]), .Z(Inst_bSbox_AND_M9_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M9_U1_U9 ( .A(Inst_bSbox_AND_M9_U1_n18), .B(
        Inst_bSbox_AND_M9_U1_n17), .ZN(new_AGEMA_signal_3123) );
  NAND2_X1 Inst_bSbox_AND_M9_U1_U8 ( .A1(Inst_bSbox_AND_M9_U1_a_reg[1]), .A2(
        Inst_bSbox_AND_M9_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M9_U1_n17) );
  XOR2_X1 Inst_bSbox_AND_M9_U1_U7 ( .A(Inst_bSbox_AND_M9_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M9_U1_z[1]), .Z(Inst_bSbox_AND_M9_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M9_U1_U6 ( .A(new_AGEMA_signal_3035), .B(
        Inst_bSbox_AND_M9_U1_n22), .ZN(Inst_bSbox_AND_M9_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M9_U1_U5 ( .A(Inst_bSbox_T17), .B(
        Inst_bSbox_AND_M9_U1_n22), .ZN(Inst_bSbox_AND_M9_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M9_U1_U4 ( .A(Fresh[11]), .ZN(Inst_bSbox_AND_M9_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M9_U1_U3 ( .A1(Inst_bSbox_T20), .A2(Inst_bSbox_T17),
        .ZN(Inst_bSbox_AND_M9_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M9_U1_U2 ( .A1(new_AGEMA_signal_3036), .A2(
        new_AGEMA_signal_3035), .ZN(Inst_bSbox_AND_M9_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M9_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M9_U1_z[0])
         );
  DFF_X1 Inst_bSbox_AND_M9_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_T20),
        .CK(clk), .Q(Inst_bSbox_AND_M9_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M9_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M9_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M9_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M9_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M9_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M9_U1_z[1])
         );
  DFF_X1 Inst_bSbox_AND_M9_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3036), .CK(clk), .Q(Inst_bSbox_AND_M9_U1_a_reg[1]) );
  DFF_X1 Inst_bSbox_AND_M9_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M9_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M9_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M9_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_M10_U1_Ins_0_U1 ( .A(Inst_bSbox_M9), .B(Inst_bSbox_M6), .Z(Inst_bSbox_M10) );
  XOR2_X1 Inst_bSbox_XOR_M10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3123), .B(
        new_AGEMA_signal_3041), .Z(new_AGEMA_signal_3262) );
  XOR2_X1 Inst_bSbox_AND_M11_U1_U16 ( .A(Fresh[12]), .B(
        Inst_bSbox_AND_M11_U1_n23), .Z(Inst_bSbox_AND_M11_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M11_U1_U15 ( .A1(new_AGEMA_signal_2850), .A2(
        Inst_bSbox_AND_M11_U1_n22), .ZN(Inst_bSbox_AND_M11_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M11_U1_U14 ( .A(Fresh[12]), .B(
        Inst_bSbox_AND_M11_U1_n21), .Z(Inst_bSbox_AND_M11_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M11_U1_U13 ( .A1(Inst_bSbox_T1), .A2(
        Inst_bSbox_AND_M11_U1_n22), .ZN(Inst_bSbox_AND_M11_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M11_U1_U12 ( .A(Inst_bSbox_AND_M11_U1_n20), .B(
        Inst_bSbox_AND_M11_U1_n19), .ZN(Inst_bSbox_M11) );
  NAND2_X1 Inst_bSbox_AND_M11_U1_U11 ( .A1(Inst_bSbox_AND_M11_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M11_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M11_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M11_U1_U10 ( .A(Inst_bSbox_AND_M11_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M11_U1_z[0]), .Z(Inst_bSbox_AND_M11_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M11_U1_U9 ( .A(Inst_bSbox_AND_M11_U1_n18), .B(
        Inst_bSbox_AND_M11_U1_n17), .ZN(new_AGEMA_signal_3043) );
  NAND2_X1 Inst_bSbox_AND_M11_U1_U8 ( .A1(Inst_bSbox_AND_M11_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M11_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M11_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M11_U1_U7 ( .A(Inst_bSbox_AND_M11_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M11_U1_z[1]), .Z(Inst_bSbox_AND_M11_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M11_U1_U6 ( .A(new_AGEMA_signal_3003), .B(
        Inst_bSbox_AND_M11_U1_n22), .ZN(Inst_bSbox_AND_M11_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M11_U1_U5 ( .A(Inst_bSbox_T15), .B(
        Inst_bSbox_AND_M11_U1_n22), .ZN(Inst_bSbox_AND_M11_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M11_U1_U4 ( .A(Fresh[13]), .ZN(
        Inst_bSbox_AND_M11_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M11_U1_U3 ( .A1(Inst_bSbox_T1), .A2(Inst_bSbox_T15),
        .ZN(Inst_bSbox_AND_M11_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M11_U1_U2 ( .A1(new_AGEMA_signal_2850), .A2(
        new_AGEMA_signal_3003), .ZN(Inst_bSbox_AND_M11_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M11_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M11_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M11_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_T1),
        .CK(clk), .Q(Inst_bSbox_AND_M11_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M11_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M11_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M11_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M11_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M11_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M11_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M11_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2850), .CK(clk), .Q(Inst_bSbox_AND_M11_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M11_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M11_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M11_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M11_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M12_U1_U16 ( .A(Fresh[14]), .B(
        Inst_bSbox_AND_M12_U1_n23), .Z(Inst_bSbox_AND_M12_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M12_U1_U15 ( .A1(new_AGEMA_signal_2853), .A2(
        Inst_bSbox_AND_M12_U1_n22), .ZN(Inst_bSbox_AND_M12_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M12_U1_U14 ( .A(Fresh[14]), .B(
        Inst_bSbox_AND_M12_U1_n21), .Z(Inst_bSbox_AND_M12_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M12_U1_U13 ( .A1(Inst_bSbox_T4), .A2(
        Inst_bSbox_AND_M12_U1_n22), .ZN(Inst_bSbox_AND_M12_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M12_U1_U12 ( .A(Inst_bSbox_AND_M12_U1_n20), .B(
        Inst_bSbox_AND_M12_U1_n19), .ZN(Inst_bSbox_M12) );
  NAND2_X1 Inst_bSbox_AND_M12_U1_U11 ( .A1(Inst_bSbox_AND_M12_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M12_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M12_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M12_U1_U10 ( .A(Inst_bSbox_AND_M12_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M12_U1_z[0]), .Z(Inst_bSbox_AND_M12_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M12_U1_U9 ( .A(Inst_bSbox_AND_M12_U1_n18), .B(
        Inst_bSbox_AND_M12_U1_n17), .ZN(new_AGEMA_signal_3044) );
  NAND2_X1 Inst_bSbox_AND_M12_U1_U8 ( .A1(Inst_bSbox_AND_M12_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M12_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M12_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M12_U1_U7 ( .A(Inst_bSbox_AND_M12_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M12_U1_z[1]), .Z(Inst_bSbox_AND_M12_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M12_U1_U6 ( .A(new_AGEMA_signal_3007), .B(
        Inst_bSbox_AND_M12_U1_n22), .ZN(Inst_bSbox_AND_M12_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M12_U1_U5 ( .A(Inst_bSbox_T27), .B(
        Inst_bSbox_AND_M12_U1_n22), .ZN(Inst_bSbox_AND_M12_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M12_U1_U4 ( .A(Fresh[15]), .ZN(
        Inst_bSbox_AND_M12_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M12_U1_U3 ( .A1(Inst_bSbox_T4), .A2(Inst_bSbox_T27),
        .ZN(Inst_bSbox_AND_M12_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M12_U1_U2 ( .A1(new_AGEMA_signal_2853), .A2(
        new_AGEMA_signal_3007), .ZN(Inst_bSbox_AND_M12_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M12_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M12_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M12_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_T4),
        .CK(clk), .Q(Inst_bSbox_AND_M12_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M12_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M12_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M12_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M12_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M12_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M12_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M12_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2853), .CK(clk), .Q(Inst_bSbox_AND_M12_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M12_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M12_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M12_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M12_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_M13_U1_Ins_0_U1 ( .A(Inst_bSbox_M12), .B(
        Inst_bSbox_M11), .Z(Inst_bSbox_M13) );
  XOR2_X1 Inst_bSbox_XOR_M13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3044), .B(
        new_AGEMA_signal_3043), .Z(new_AGEMA_signal_3124) );
  XOR2_X1 Inst_bSbox_AND_M14_U1_U16 ( .A(Fresh[16]), .B(
        Inst_bSbox_AND_M14_U1_n23), .Z(Inst_bSbox_AND_M14_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M14_U1_U15 ( .A1(new_AGEMA_signal_2851), .A2(
        Inst_bSbox_AND_M14_U1_n22), .ZN(Inst_bSbox_AND_M14_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M14_U1_U14 ( .A(Fresh[16]), .B(
        Inst_bSbox_AND_M14_U1_n21), .Z(Inst_bSbox_AND_M14_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M14_U1_U13 ( .A1(Inst_bSbox_T2), .A2(
        Inst_bSbox_AND_M14_U1_n22), .ZN(Inst_bSbox_AND_M14_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M14_U1_U12 ( .A(Inst_bSbox_AND_M14_U1_n20), .B(
        Inst_bSbox_AND_M14_U1_n19), .ZN(Inst_bSbox_M14) );
  NAND2_X1 Inst_bSbox_AND_M14_U1_U11 ( .A1(Inst_bSbox_AND_M14_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M14_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M14_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M14_U1_U10 ( .A(Inst_bSbox_AND_M14_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M14_U1_z[0]), .Z(Inst_bSbox_AND_M14_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M14_U1_U9 ( .A(Inst_bSbox_AND_M14_U1_n18), .B(
        Inst_bSbox_AND_M14_U1_n17), .ZN(new_AGEMA_signal_3125) );
  NAND2_X1 Inst_bSbox_AND_M14_U1_U8 ( .A1(Inst_bSbox_AND_M14_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M14_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M14_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M14_U1_U7 ( .A(Inst_bSbox_AND_M14_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M14_U1_z[1]), .Z(Inst_bSbox_AND_M14_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M14_U1_U6 ( .A(new_AGEMA_signal_3033), .B(
        Inst_bSbox_AND_M14_U1_n22), .ZN(Inst_bSbox_AND_M14_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M14_U1_U5 ( .A(Inst_bSbox_T10), .B(
        Inst_bSbox_AND_M14_U1_n22), .ZN(Inst_bSbox_AND_M14_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M14_U1_U4 ( .A(Fresh[17]), .ZN(
        Inst_bSbox_AND_M14_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M14_U1_U3 ( .A1(Inst_bSbox_T2), .A2(Inst_bSbox_T10),
        .ZN(Inst_bSbox_AND_M14_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M14_U1_U2 ( .A1(new_AGEMA_signal_2851), .A2(
        new_AGEMA_signal_3033), .ZN(Inst_bSbox_AND_M14_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M14_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M14_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M14_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_T2),
        .CK(clk), .Q(Inst_bSbox_AND_M14_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M14_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M14_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M14_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M14_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M14_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M14_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M14_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2851), .CK(clk), .Q(Inst_bSbox_AND_M14_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M14_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M14_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M14_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M14_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_M15_U1_Ins_0_U1 ( .A(Inst_bSbox_M14), .B(
        Inst_bSbox_M11), .Z(Inst_bSbox_M15) );
  XOR2_X1 Inst_bSbox_XOR_M15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3125), .B(
        new_AGEMA_signal_3043), .Z(new_AGEMA_signal_3263) );
  XOR2_X1 Inst_bSbox_XOR_M16_U1_Ins_0_U1 ( .A(Inst_bSbox_M3), .B(Inst_bSbox_M2), .Z(Inst_bSbox_M16) );
  XOR2_X1 Inst_bSbox_XOR_M16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3120), .B(
        new_AGEMA_signal_3119), .Z(new_AGEMA_signal_3264) );
  XOR2_X1 Inst_bSbox_XOR_M17_U1_Ins_0_U1 ( .A(Inst_bSbox_M5), .B(
        new_AGEMA_signal_3606), .Z(Inst_bSbox_M17) );
  XOR2_X1 Inst_bSbox_XOR_M17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3121), .B(
        new_AGEMA_signal_3607), .Z(new_AGEMA_signal_3265) );
  XOR2_X1 Inst_bSbox_XOR_M18_U1_Ins_0_U1 ( .A(Inst_bSbox_M8), .B(Inst_bSbox_M7), .Z(Inst_bSbox_M18) );
  XOR2_X1 Inst_bSbox_XOR_M18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3122), .B(
        new_AGEMA_signal_3042), .Z(new_AGEMA_signal_3266) );
  XOR2_X1 Inst_bSbox_XOR_M19_U1_Ins_0_U1 ( .A(Inst_bSbox_M10), .B(
        Inst_bSbox_M15), .Z(Inst_bSbox_M19) );
  XOR2_X1 Inst_bSbox_XOR_M19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3262), .B(
        new_AGEMA_signal_3263), .Z(new_AGEMA_signal_3371) );
  XOR2_X1 Inst_bSbox_XOR_M20_U1_Ins_0_U1 ( .A(Inst_bSbox_M16), .B(
        Inst_bSbox_M13), .Z(Inst_bSbox_M20) );
  XOR2_X1 Inst_bSbox_XOR_M20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3264), .B(
        new_AGEMA_signal_3124), .Z(new_AGEMA_signal_3372) );
  XOR2_X1 Inst_bSbox_XOR_M21_U1_Ins_0_U1 ( .A(Inst_bSbox_M17), .B(
        Inst_bSbox_M15), .Z(Inst_bSbox_M21) );
  XOR2_X1 Inst_bSbox_XOR_M21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3265), .B(
        new_AGEMA_signal_3263), .Z(new_AGEMA_signal_3373) );
  XOR2_X1 Inst_bSbox_XOR_M22_U1_Ins_0_U1 ( .A(Inst_bSbox_M18), .B(
        Inst_bSbox_M13), .Z(Inst_bSbox_M22) );
  XOR2_X1 Inst_bSbox_XOR_M22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3266), .B(
        new_AGEMA_signal_3124), .Z(new_AGEMA_signal_3374) );
  XOR2_X1 Inst_bSbox_XOR_M23_U1_Ins_0_U1 ( .A(Inst_bSbox_M19), .B(
        new_AGEMA_signal_3608), .Z(Inst_bSbox_M23) );
  XOR2_X1 Inst_bSbox_XOR_M23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3371), .B(
        new_AGEMA_signal_3609), .Z(new_AGEMA_signal_3383) );
  XOR2_X1 Inst_bSbox_XOR_M24_U1_Ins_0_U1 ( .A(Inst_bSbox_M22), .B(
        Inst_bSbox_M23), .Z(Inst_bSbox_M24) );
  XOR2_X1 Inst_bSbox_XOR_M24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3374), .B(
        new_AGEMA_signal_3383), .Z(new_AGEMA_signal_3387) );
  XOR2_X1 Inst_bSbox_XOR_M27_U1_Ins_0_U1 ( .A(Inst_bSbox_M20), .B(
        Inst_bSbox_M21), .Z(Inst_bSbox_M27) );
  XOR2_X1 Inst_bSbox_XOR_M27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3372), .B(
        new_AGEMA_signal_3373), .Z(new_AGEMA_signal_3385) );
  DFF_X1 new_AGEMA_reg_buffer_1714_s_current_state_reg ( .D(Inst_bSbox_T14),
        .CK(clk), .Q(new_AGEMA_signal_3602) );
  DFF_X1 new_AGEMA_reg_buffer_1715_s_current_state_reg ( .D(
        new_AGEMA_signal_3034), .CK(clk), .Q(new_AGEMA_signal_3603) );
  DFF_X1 new_AGEMA_reg_buffer_1716_s_current_state_reg ( .D(Inst_bSbox_T26),
        .CK(clk), .Q(new_AGEMA_signal_3604) );
  DFF_X1 new_AGEMA_reg_buffer_1717_s_current_state_reg ( .D(
        new_AGEMA_signal_3038), .CK(clk), .Q(new_AGEMA_signal_3605) );
  DFF_X1 new_AGEMA_reg_buffer_1718_s_current_state_reg ( .D(Inst_bSbox_T24),
        .CK(clk), .Q(new_AGEMA_signal_3606) );
  DFF_X1 new_AGEMA_reg_buffer_1719_s_current_state_reg ( .D(
        new_AGEMA_signal_3117), .CK(clk), .Q(new_AGEMA_signal_3607) );
  DFF_X1 new_AGEMA_reg_buffer_1720_s_current_state_reg ( .D(Inst_bSbox_T25),
        .CK(clk), .Q(new_AGEMA_signal_3608) );
  DFF_X1 new_AGEMA_reg_buffer_1721_s_current_state_reg ( .D(
        new_AGEMA_signal_3118), .CK(clk), .Q(new_AGEMA_signal_3609) );
  DFF_X1 new_AGEMA_reg_buffer_1738_s_current_state_reg ( .D(n188), .CK(clk),
        .Q(new_AGEMA_signal_3626) );
  DFF_X1 new_AGEMA_reg_buffer_1742_s_current_state_reg ( .D(
        StateOutXORroundKey[0]), .CK(clk), .Q(new_AGEMA_signal_3630) );
  DFF_X1 new_AGEMA_reg_buffer_1746_s_current_state_reg ( .D(
        new_AGEMA_signal_1984), .CK(clk), .Q(new_AGEMA_signal_3634) );
  DFF_X1 new_AGEMA_reg_buffer_1750_s_current_state_reg ( .D(
        StateOutXORroundKey[1]), .CK(clk), .Q(new_AGEMA_signal_3638) );
  DFF_X1 new_AGEMA_reg_buffer_1754_s_current_state_reg ( .D(
        new_AGEMA_signal_1987), .CK(clk), .Q(new_AGEMA_signal_3642) );
  DFF_X1 new_AGEMA_reg_buffer_1758_s_current_state_reg ( .D(
        StateOutXORroundKey[2]), .CK(clk), .Q(new_AGEMA_signal_3646) );
  DFF_X1 new_AGEMA_reg_buffer_1762_s_current_state_reg ( .D(
        new_AGEMA_signal_1990), .CK(clk), .Q(new_AGEMA_signal_3650) );
  DFF_X1 new_AGEMA_reg_buffer_1766_s_current_state_reg ( .D(
        StateOutXORroundKey[3]), .CK(clk), .Q(new_AGEMA_signal_3654) );
  DFF_X1 new_AGEMA_reg_buffer_1770_s_current_state_reg ( .D(
        new_AGEMA_signal_1993), .CK(clk), .Q(new_AGEMA_signal_3658) );
  DFF_X1 new_AGEMA_reg_buffer_1774_s_current_state_reg ( .D(
        StateOutXORroundKey[4]), .CK(clk), .Q(new_AGEMA_signal_3662) );
  DFF_X1 new_AGEMA_reg_buffer_1778_s_current_state_reg ( .D(
        new_AGEMA_signal_1996), .CK(clk), .Q(new_AGEMA_signal_3666) );
  DFF_X1 new_AGEMA_reg_buffer_1782_s_current_state_reg ( .D(
        StateOutXORroundKey[5]), .CK(clk), .Q(new_AGEMA_signal_3670) );
  DFF_X1 new_AGEMA_reg_buffer_1786_s_current_state_reg ( .D(
        new_AGEMA_signal_1999), .CK(clk), .Q(new_AGEMA_signal_3674) );
  DFF_X1 new_AGEMA_reg_buffer_1790_s_current_state_reg ( .D(
        StateOutXORroundKey[6]), .CK(clk), .Q(new_AGEMA_signal_3678) );
  DFF_X1 new_AGEMA_reg_buffer_1794_s_current_state_reg ( .D(
        new_AGEMA_signal_2002), .CK(clk), .Q(new_AGEMA_signal_3682) );
  DFF_X1 new_AGEMA_reg_buffer_1798_s_current_state_reg ( .D(
        StateOutXORroundKey[7]), .CK(clk), .Q(new_AGEMA_signal_3686) );
  DFF_X1 new_AGEMA_reg_buffer_1802_s_current_state_reg ( .D(
        new_AGEMA_signal_2005), .CK(clk), .Q(new_AGEMA_signal_3690) );
  DFF_X1 new_AGEMA_reg_buffer_1806_s_current_state_reg ( .D(n250), .CK(clk),
        .Q(new_AGEMA_signal_3694) );
  DFF_X1 new_AGEMA_reg_buffer_1810_s_current_state_reg ( .D(ciphertext_s0[8]),
        .CK(clk), .Q(new_AGEMA_signal_3698) );
  DFF_X1 new_AGEMA_reg_buffer_1814_s_current_state_reg ( .D(ciphertext_s1[8]),
        .CK(clk), .Q(new_AGEMA_signal_3702) );
  DFF_X1 new_AGEMA_reg_buffer_1818_s_current_state_reg ( .D(ciphertext_s0[9]),
        .CK(clk), .Q(new_AGEMA_signal_3706) );
  DFF_X1 new_AGEMA_reg_buffer_1822_s_current_state_reg ( .D(ciphertext_s1[9]),
        .CK(clk), .Q(new_AGEMA_signal_3710) );
  DFF_X1 new_AGEMA_reg_buffer_1826_s_current_state_reg ( .D(ciphertext_s0[10]),
        .CK(clk), .Q(new_AGEMA_signal_3714) );
  DFF_X1 new_AGEMA_reg_buffer_1830_s_current_state_reg ( .D(ciphertext_s1[10]),
        .CK(clk), .Q(new_AGEMA_signal_3718) );
  DFF_X1 new_AGEMA_reg_buffer_1834_s_current_state_reg ( .D(ciphertext_s0[11]),
        .CK(clk), .Q(new_AGEMA_signal_3722) );
  DFF_X1 new_AGEMA_reg_buffer_1838_s_current_state_reg ( .D(ciphertext_s1[11]),
        .CK(clk), .Q(new_AGEMA_signal_3726) );
  DFF_X1 new_AGEMA_reg_buffer_1842_s_current_state_reg ( .D(ciphertext_s0[12]),
        .CK(clk), .Q(new_AGEMA_signal_3730) );
  DFF_X1 new_AGEMA_reg_buffer_1846_s_current_state_reg ( .D(ciphertext_s1[12]),
        .CK(clk), .Q(new_AGEMA_signal_3734) );
  DFF_X1 new_AGEMA_reg_buffer_1850_s_current_state_reg ( .D(ciphertext_s0[13]),
        .CK(clk), .Q(new_AGEMA_signal_3738) );
  DFF_X1 new_AGEMA_reg_buffer_1854_s_current_state_reg ( .D(ciphertext_s1[13]),
        .CK(clk), .Q(new_AGEMA_signal_3742) );
  DFF_X1 new_AGEMA_reg_buffer_1858_s_current_state_reg ( .D(ciphertext_s0[14]),
        .CK(clk), .Q(new_AGEMA_signal_3746) );
  DFF_X1 new_AGEMA_reg_buffer_1862_s_current_state_reg ( .D(ciphertext_s1[14]),
        .CK(clk), .Q(new_AGEMA_signal_3750) );
  DFF_X1 new_AGEMA_reg_buffer_1866_s_current_state_reg ( .D(ciphertext_s0[15]),
        .CK(clk), .Q(new_AGEMA_signal_3754) );
  DFF_X1 new_AGEMA_reg_buffer_1870_s_current_state_reg ( .D(ciphertext_s1[15]),
        .CK(clk), .Q(new_AGEMA_signal_3758) );
  DFF_X1 new_AGEMA_reg_buffer_1874_s_current_state_reg ( .D(n199), .CK(clk),
        .Q(new_AGEMA_signal_3762) );
  DFF_X1 new_AGEMA_reg_buffer_1878_s_current_state_reg ( .D(StateInMC[0]),
        .CK(clk), .Q(new_AGEMA_signal_3766) );
  DFF_X1 new_AGEMA_reg_buffer_1882_s_current_state_reg ( .D(
        new_AGEMA_signal_2860), .CK(clk), .Q(new_AGEMA_signal_3770) );
  DFF_X1 new_AGEMA_reg_buffer_1886_s_current_state_reg ( .D(StateInMC[1]),
        .CK(clk), .Q(new_AGEMA_signal_3774) );
  DFF_X1 new_AGEMA_reg_buffer_1890_s_current_state_reg ( .D(
        new_AGEMA_signal_2861), .CK(clk), .Q(new_AGEMA_signal_3778) );
  DFF_X1 new_AGEMA_reg_buffer_1894_s_current_state_reg ( .D(StateInMC[2]),
        .CK(clk), .Q(new_AGEMA_signal_3782) );
  DFF_X1 new_AGEMA_reg_buffer_1898_s_current_state_reg ( .D(
        new_AGEMA_signal_2834), .CK(clk), .Q(new_AGEMA_signal_3786) );
  DFF_X1 new_AGEMA_reg_buffer_1902_s_current_state_reg ( .D(StateInMC[3]),
        .CK(clk), .Q(new_AGEMA_signal_3790) );
  DFF_X1 new_AGEMA_reg_buffer_1906_s_current_state_reg ( .D(
        new_AGEMA_signal_2862), .CK(clk), .Q(new_AGEMA_signal_3794) );
  DFF_X1 new_AGEMA_reg_buffer_1910_s_current_state_reg ( .D(StateInMC[4]),
        .CK(clk), .Q(new_AGEMA_signal_3798) );
  DFF_X1 new_AGEMA_reg_buffer_1914_s_current_state_reg ( .D(
        new_AGEMA_signal_2863), .CK(clk), .Q(new_AGEMA_signal_3802) );
  DFF_X1 new_AGEMA_reg_buffer_1918_s_current_state_reg ( .D(StateInMC[5]),
        .CK(clk), .Q(new_AGEMA_signal_3806) );
  DFF_X1 new_AGEMA_reg_buffer_1922_s_current_state_reg ( .D(
        new_AGEMA_signal_2835), .CK(clk), .Q(new_AGEMA_signal_3810) );
  DFF_X1 new_AGEMA_reg_buffer_1926_s_current_state_reg ( .D(StateInMC[6]),
        .CK(clk), .Q(new_AGEMA_signal_3814) );
  DFF_X1 new_AGEMA_reg_buffer_1930_s_current_state_reg ( .D(
        new_AGEMA_signal_2836), .CK(clk), .Q(new_AGEMA_signal_3818) );
  DFF_X1 new_AGEMA_reg_buffer_1934_s_current_state_reg ( .D(StateInMC[7]),
        .CK(clk), .Q(new_AGEMA_signal_3822) );
  DFF_X1 new_AGEMA_reg_buffer_1938_s_current_state_reg ( .D(
        new_AGEMA_signal_2837), .CK(clk), .Q(new_AGEMA_signal_3826) );
  DFF_X1 new_AGEMA_reg_buffer_1942_s_current_state_reg ( .D(n294), .CK(clk),
        .Q(new_AGEMA_signal_3830) );
  DFF_X1 new_AGEMA_reg_buffer_1946_s_current_state_reg ( .D(plaintext_s0[0]),
        .CK(clk), .Q(new_AGEMA_signal_3834) );
  DFF_X1 new_AGEMA_reg_buffer_1950_s_current_state_reg ( .D(plaintext_s1[0]),
        .CK(clk), .Q(new_AGEMA_signal_3838) );
  DFF_X1 new_AGEMA_reg_buffer_1954_s_current_state_reg ( .D(plaintext_s0[1]),
        .CK(clk), .Q(new_AGEMA_signal_3842) );
  DFF_X1 new_AGEMA_reg_buffer_1958_s_current_state_reg ( .D(plaintext_s1[1]),
        .CK(clk), .Q(new_AGEMA_signal_3846) );
  DFF_X1 new_AGEMA_reg_buffer_1962_s_current_state_reg ( .D(plaintext_s0[2]),
        .CK(clk), .Q(new_AGEMA_signal_3850) );
  DFF_X1 new_AGEMA_reg_buffer_1966_s_current_state_reg ( .D(plaintext_s1[2]),
        .CK(clk), .Q(new_AGEMA_signal_3854) );
  DFF_X1 new_AGEMA_reg_buffer_1970_s_current_state_reg ( .D(plaintext_s0[3]),
        .CK(clk), .Q(new_AGEMA_signal_3858) );
  DFF_X1 new_AGEMA_reg_buffer_1974_s_current_state_reg ( .D(plaintext_s1[3]),
        .CK(clk), .Q(new_AGEMA_signal_3862) );
  DFF_X1 new_AGEMA_reg_buffer_1978_s_current_state_reg ( .D(plaintext_s0[4]),
        .CK(clk), .Q(new_AGEMA_signal_3866) );
  DFF_X1 new_AGEMA_reg_buffer_1982_s_current_state_reg ( .D(plaintext_s1[4]),
        .CK(clk), .Q(new_AGEMA_signal_3870) );
  DFF_X1 new_AGEMA_reg_buffer_1986_s_current_state_reg ( .D(plaintext_s0[5]),
        .CK(clk), .Q(new_AGEMA_signal_3874) );
  DFF_X1 new_AGEMA_reg_buffer_1990_s_current_state_reg ( .D(plaintext_s1[5]),
        .CK(clk), .Q(new_AGEMA_signal_3878) );
  DFF_X1 new_AGEMA_reg_buffer_1994_s_current_state_reg ( .D(plaintext_s0[6]),
        .CK(clk), .Q(new_AGEMA_signal_3882) );
  DFF_X1 new_AGEMA_reg_buffer_1998_s_current_state_reg ( .D(plaintext_s1[6]),
        .CK(clk), .Q(new_AGEMA_signal_3886) );
  DFF_X1 new_AGEMA_reg_buffer_2002_s_current_state_reg ( .D(plaintext_s0[7]),
        .CK(clk), .Q(new_AGEMA_signal_3890) );
  DFF_X1 new_AGEMA_reg_buffer_2006_s_current_state_reg ( .D(plaintext_s1[7]),
        .CK(clk), .Q(new_AGEMA_signal_3894) );
  DFF_X1 new_AGEMA_reg_buffer_2010_s_current_state_reg ( .D(keyStateIn[7]),
        .CK(clk), .Q(new_AGEMA_signal_3898) );
  DFF_X1 new_AGEMA_reg_buffer_2014_s_current_state_reg ( .D(
        new_AGEMA_signal_2004), .CK(clk), .Q(new_AGEMA_signal_3902) );
  DFF_X1 new_AGEMA_reg_buffer_2018_s_current_state_reg ( .D(roundConstant[7]),
        .CK(clk), .Q(new_AGEMA_signal_3906) );
  DFF_X1 new_AGEMA_reg_buffer_2022_s_current_state_reg ( .D(keyStateIn[6]),
        .CK(clk), .Q(new_AGEMA_signal_3910) );
  DFF_X1 new_AGEMA_reg_buffer_2026_s_current_state_reg ( .D(
        new_AGEMA_signal_2001), .CK(clk), .Q(new_AGEMA_signal_3914) );
  DFF_X1 new_AGEMA_reg_buffer_2030_s_current_state_reg ( .D(roundConstant[6]),
        .CK(clk), .Q(new_AGEMA_signal_3918) );
  DFF_X1 new_AGEMA_reg_buffer_2034_s_current_state_reg ( .D(keyStateIn[5]),
        .CK(clk), .Q(new_AGEMA_signal_3922) );
  DFF_X1 new_AGEMA_reg_buffer_2038_s_current_state_reg ( .D(
        new_AGEMA_signal_1998), .CK(clk), .Q(new_AGEMA_signal_3926) );
  DFF_X1 new_AGEMA_reg_buffer_2042_s_current_state_reg ( .D(roundConstant[5]),
        .CK(clk), .Q(new_AGEMA_signal_3930) );
  DFF_X1 new_AGEMA_reg_buffer_2046_s_current_state_reg ( .D(keyStateIn[4]),
        .CK(clk), .Q(new_AGEMA_signal_3934) );
  DFF_X1 new_AGEMA_reg_buffer_2050_s_current_state_reg ( .D(
        new_AGEMA_signal_1995), .CK(clk), .Q(new_AGEMA_signal_3938) );
  DFF_X1 new_AGEMA_reg_buffer_2054_s_current_state_reg ( .D(roundConstant[4]),
        .CK(clk), .Q(new_AGEMA_signal_3942) );
  DFF_X1 new_AGEMA_reg_buffer_2058_s_current_state_reg ( .D(keyStateIn[3]),
        .CK(clk), .Q(new_AGEMA_signal_3946) );
  DFF_X1 new_AGEMA_reg_buffer_2062_s_current_state_reg ( .D(
        new_AGEMA_signal_1992), .CK(clk), .Q(new_AGEMA_signal_3950) );
  DFF_X1 new_AGEMA_reg_buffer_2066_s_current_state_reg ( .D(roundConstant[3]),
        .CK(clk), .Q(new_AGEMA_signal_3954) );
  DFF_X1 new_AGEMA_reg_buffer_2070_s_current_state_reg ( .D(keyStateIn[2]),
        .CK(clk), .Q(new_AGEMA_signal_3958) );
  DFF_X1 new_AGEMA_reg_buffer_2074_s_current_state_reg ( .D(
        new_AGEMA_signal_1989), .CK(clk), .Q(new_AGEMA_signal_3962) );
  DFF_X1 new_AGEMA_reg_buffer_2078_s_current_state_reg ( .D(roundConstant[2]),
        .CK(clk), .Q(new_AGEMA_signal_3966) );
  DFF_X1 new_AGEMA_reg_buffer_2082_s_current_state_reg ( .D(keyStateIn[1]),
        .CK(clk), .Q(new_AGEMA_signal_3970) );
  DFF_X1 new_AGEMA_reg_buffer_2086_s_current_state_reg ( .D(
        new_AGEMA_signal_1986), .CK(clk), .Q(new_AGEMA_signal_3974) );
  DFF_X1 new_AGEMA_reg_buffer_2090_s_current_state_reg ( .D(roundConstant[1]),
        .CK(clk), .Q(new_AGEMA_signal_3978) );
  DFF_X1 new_AGEMA_reg_buffer_2094_s_current_state_reg ( .D(keyStateIn[0]),
        .CK(clk), .Q(new_AGEMA_signal_3982) );
  DFF_X1 new_AGEMA_reg_buffer_2098_s_current_state_reg ( .D(
        new_AGEMA_signal_1983), .CK(clk), .Q(new_AGEMA_signal_3986) );
  DFF_X1 new_AGEMA_reg_buffer_2102_s_current_state_reg ( .D(roundConstant[0]),
        .CK(clk), .Q(new_AGEMA_signal_3990) );
  DFF_X1 new_AGEMA_reg_buffer_2106_s_current_state_reg ( .D(n253), .CK(clk),
        .Q(new_AGEMA_signal_3994) );
  DFF_X1 new_AGEMA_reg_buffer_2110_s_current_state_reg ( .D(
        KeyArray_outS30ser[0]), .CK(clk), .Q(new_AGEMA_signal_3998) );
  DFF_X1 new_AGEMA_reg_buffer_2114_s_current_state_reg ( .D(
        new_AGEMA_signal_2683), .CK(clk), .Q(new_AGEMA_signal_4002) );
  DFF_X1 new_AGEMA_reg_buffer_2118_s_current_state_reg ( .D(n200), .CK(clk),
        .Q(new_AGEMA_signal_4006) );
  DFF_X1 new_AGEMA_reg_buffer_2122_s_current_state_reg ( .D(
        KeyArray_inS30ser[0]), .CK(clk), .Q(new_AGEMA_signal_4010) );
  DFF_X1 new_AGEMA_reg_buffer_2126_s_current_state_reg ( .D(
        new_AGEMA_signal_2708), .CK(clk), .Q(new_AGEMA_signal_4014) );
  DFF_X1 new_AGEMA_reg_buffer_2130_s_current_state_reg ( .D(
        KeyArray_outS30ser[1]), .CK(clk), .Q(new_AGEMA_signal_4018) );
  DFF_X1 new_AGEMA_reg_buffer_2134_s_current_state_reg ( .D(
        new_AGEMA_signal_2686), .CK(clk), .Q(new_AGEMA_signal_4022) );
  DFF_X1 new_AGEMA_reg_buffer_2138_s_current_state_reg ( .D(
        KeyArray_inS30ser[1]), .CK(clk), .Q(new_AGEMA_signal_4026) );
  DFF_X1 new_AGEMA_reg_buffer_2142_s_current_state_reg ( .D(
        new_AGEMA_signal_2711), .CK(clk), .Q(new_AGEMA_signal_4030) );
  DFF_X1 new_AGEMA_reg_buffer_2146_s_current_state_reg ( .D(
        KeyArray_outS30ser[2]), .CK(clk), .Q(new_AGEMA_signal_4034) );
  DFF_X1 new_AGEMA_reg_buffer_2150_s_current_state_reg ( .D(
        new_AGEMA_signal_2689), .CK(clk), .Q(new_AGEMA_signal_4038) );
  DFF_X1 new_AGEMA_reg_buffer_2154_s_current_state_reg ( .D(
        KeyArray_inS30ser[2]), .CK(clk), .Q(new_AGEMA_signal_4042) );
  DFF_X1 new_AGEMA_reg_buffer_2158_s_current_state_reg ( .D(
        new_AGEMA_signal_2714), .CK(clk), .Q(new_AGEMA_signal_4046) );
  DFF_X1 new_AGEMA_reg_buffer_2162_s_current_state_reg ( .D(
        KeyArray_outS30ser[3]), .CK(clk), .Q(new_AGEMA_signal_4050) );
  DFF_X1 new_AGEMA_reg_buffer_2166_s_current_state_reg ( .D(
        new_AGEMA_signal_2692), .CK(clk), .Q(new_AGEMA_signal_4054) );
  DFF_X1 new_AGEMA_reg_buffer_2170_s_current_state_reg ( .D(
        KeyArray_inS30ser[3]), .CK(clk), .Q(new_AGEMA_signal_4058) );
  DFF_X1 new_AGEMA_reg_buffer_2174_s_current_state_reg ( .D(
        new_AGEMA_signal_2717), .CK(clk), .Q(new_AGEMA_signal_4062) );
  DFF_X1 new_AGEMA_reg_buffer_2178_s_current_state_reg ( .D(
        KeyArray_outS30ser[4]), .CK(clk), .Q(new_AGEMA_signal_4066) );
  DFF_X1 new_AGEMA_reg_buffer_2182_s_current_state_reg ( .D(
        new_AGEMA_signal_2695), .CK(clk), .Q(new_AGEMA_signal_4070) );
  DFF_X1 new_AGEMA_reg_buffer_2186_s_current_state_reg ( .D(
        KeyArray_inS30ser[4]), .CK(clk), .Q(new_AGEMA_signal_4074) );
  DFF_X1 new_AGEMA_reg_buffer_2190_s_current_state_reg ( .D(
        new_AGEMA_signal_2720), .CK(clk), .Q(new_AGEMA_signal_4078) );
  DFF_X1 new_AGEMA_reg_buffer_2194_s_current_state_reg ( .D(
        KeyArray_outS30ser[5]), .CK(clk), .Q(new_AGEMA_signal_4082) );
  DFF_X1 new_AGEMA_reg_buffer_2198_s_current_state_reg ( .D(
        new_AGEMA_signal_2698), .CK(clk), .Q(new_AGEMA_signal_4086) );
  DFF_X1 new_AGEMA_reg_buffer_2202_s_current_state_reg ( .D(
        KeyArray_inS30ser[5]), .CK(clk), .Q(new_AGEMA_signal_4090) );
  DFF_X1 new_AGEMA_reg_buffer_2206_s_current_state_reg ( .D(
        new_AGEMA_signal_2723), .CK(clk), .Q(new_AGEMA_signal_4094) );
  DFF_X1 new_AGEMA_reg_buffer_2210_s_current_state_reg ( .D(
        KeyArray_outS30ser[6]), .CK(clk), .Q(new_AGEMA_signal_4098) );
  DFF_X1 new_AGEMA_reg_buffer_2214_s_current_state_reg ( .D(
        new_AGEMA_signal_2701), .CK(clk), .Q(new_AGEMA_signal_4102) );
  DFF_X1 new_AGEMA_reg_buffer_2218_s_current_state_reg ( .D(
        KeyArray_inS30ser[6]), .CK(clk), .Q(new_AGEMA_signal_4106) );
  DFF_X1 new_AGEMA_reg_buffer_2222_s_current_state_reg ( .D(
        new_AGEMA_signal_2726), .CK(clk), .Q(new_AGEMA_signal_4110) );
  DFF_X1 new_AGEMA_reg_buffer_2226_s_current_state_reg ( .D(
        KeyArray_outS30ser[7]), .CK(clk), .Q(new_AGEMA_signal_4114) );
  DFF_X1 new_AGEMA_reg_buffer_2230_s_current_state_reg ( .D(
        new_AGEMA_signal_2704), .CK(clk), .Q(new_AGEMA_signal_4118) );
  DFF_X1 new_AGEMA_reg_buffer_2234_s_current_state_reg ( .D(
        KeyArray_inS30ser[7]), .CK(clk), .Q(new_AGEMA_signal_4122) );
  DFF_X1 new_AGEMA_reg_buffer_2238_s_current_state_reg ( .D(
        new_AGEMA_signal_2729), .CK(clk), .Q(new_AGEMA_signal_4126) );
  DFF_X1 new_AGEMA_reg_buffer_2242_s_current_state_reg ( .D(Inst_bSbox_T6),
        .CK(clk), .Q(new_AGEMA_signal_4130) );
  DFF_X1 new_AGEMA_reg_buffer_2245_s_current_state_reg ( .D(
        new_AGEMA_signal_3000), .CK(clk), .Q(new_AGEMA_signal_4133) );
  DFF_X1 new_AGEMA_reg_buffer_2248_s_current_state_reg ( .D(Inst_bSbox_T8),
        .CK(clk), .Q(new_AGEMA_signal_4136) );
  DFF_X1 new_AGEMA_reg_buffer_2251_s_current_state_reg ( .D(
        new_AGEMA_signal_3032), .CK(clk), .Q(new_AGEMA_signal_4139) );
  DFF_X1 new_AGEMA_reg_buffer_2254_s_current_state_reg ( .D(SboxIn[0]), .CK(
        clk), .Q(new_AGEMA_signal_4142) );
  DFF_X1 new_AGEMA_reg_buffer_2257_s_current_state_reg ( .D(
        new_AGEMA_signal_2826), .CK(clk), .Q(new_AGEMA_signal_4145) );
  DFF_X1 new_AGEMA_reg_buffer_2260_s_current_state_reg ( .D(Inst_bSbox_T16),
        .CK(clk), .Q(new_AGEMA_signal_4148) );
  DFF_X1 new_AGEMA_reg_buffer_2263_s_current_state_reg ( .D(
        new_AGEMA_signal_3004), .CK(clk), .Q(new_AGEMA_signal_4151) );
  DFF_X1 new_AGEMA_reg_buffer_2266_s_current_state_reg ( .D(Inst_bSbox_T9),
        .CK(clk), .Q(new_AGEMA_signal_4154) );
  DFF_X1 new_AGEMA_reg_buffer_2269_s_current_state_reg ( .D(
        new_AGEMA_signal_3001), .CK(clk), .Q(new_AGEMA_signal_4157) );
  DFF_X1 new_AGEMA_reg_buffer_2272_s_current_state_reg ( .D(Inst_bSbox_T17),
        .CK(clk), .Q(new_AGEMA_signal_4160) );
  DFF_X1 new_AGEMA_reg_buffer_2275_s_current_state_reg ( .D(
        new_AGEMA_signal_3035), .CK(clk), .Q(new_AGEMA_signal_4163) );
  DFF_X1 new_AGEMA_reg_buffer_2278_s_current_state_reg ( .D(Inst_bSbox_T15),
        .CK(clk), .Q(new_AGEMA_signal_4166) );
  DFF_X1 new_AGEMA_reg_buffer_2281_s_current_state_reg ( .D(
        new_AGEMA_signal_3003), .CK(clk), .Q(new_AGEMA_signal_4169) );
  DFF_X1 new_AGEMA_reg_buffer_2284_s_current_state_reg ( .D(Inst_bSbox_T27),
        .CK(clk), .Q(new_AGEMA_signal_4172) );
  DFF_X1 new_AGEMA_reg_buffer_2287_s_current_state_reg ( .D(
        new_AGEMA_signal_3007), .CK(clk), .Q(new_AGEMA_signal_4175) );
  DFF_X1 new_AGEMA_reg_buffer_2290_s_current_state_reg ( .D(Inst_bSbox_T10),
        .CK(clk), .Q(new_AGEMA_signal_4178) );
  DFF_X1 new_AGEMA_reg_buffer_2293_s_current_state_reg ( .D(
        new_AGEMA_signal_3033), .CK(clk), .Q(new_AGEMA_signal_4181) );
  DFF_X1 new_AGEMA_reg_buffer_2296_s_current_state_reg ( .D(Inst_bSbox_T13),
        .CK(clk), .Q(new_AGEMA_signal_4184) );
  DFF_X1 new_AGEMA_reg_buffer_2299_s_current_state_reg ( .D(
        new_AGEMA_signal_3002), .CK(clk), .Q(new_AGEMA_signal_4187) );
  DFF_X1 new_AGEMA_reg_buffer_2302_s_current_state_reg ( .D(Inst_bSbox_T23),
        .CK(clk), .Q(new_AGEMA_signal_4190) );
  DFF_X1 new_AGEMA_reg_buffer_2305_s_current_state_reg ( .D(
        new_AGEMA_signal_3037), .CK(clk), .Q(new_AGEMA_signal_4193) );
  DFF_X1 new_AGEMA_reg_buffer_2308_s_current_state_reg ( .D(Inst_bSbox_T19),
        .CK(clk), .Q(new_AGEMA_signal_4196) );
  DFF_X1 new_AGEMA_reg_buffer_2311_s_current_state_reg ( .D(
        new_AGEMA_signal_3005), .CK(clk), .Q(new_AGEMA_signal_4199) );
  DFF_X1 new_AGEMA_reg_buffer_2314_s_current_state_reg ( .D(Inst_bSbox_T3),
        .CK(clk), .Q(new_AGEMA_signal_4202) );
  DFF_X1 new_AGEMA_reg_buffer_2317_s_current_state_reg ( .D(
        new_AGEMA_signal_2852), .CK(clk), .Q(new_AGEMA_signal_4205) );
  DFF_X1 new_AGEMA_reg_buffer_2320_s_current_state_reg ( .D(Inst_bSbox_T22),
        .CK(clk), .Q(new_AGEMA_signal_4208) );
  DFF_X1 new_AGEMA_reg_buffer_2323_s_current_state_reg ( .D(
        new_AGEMA_signal_3006), .CK(clk), .Q(new_AGEMA_signal_4211) );
  DFF_X1 new_AGEMA_reg_buffer_2326_s_current_state_reg ( .D(Inst_bSbox_T20),
        .CK(clk), .Q(new_AGEMA_signal_4214) );
  DFF_X1 new_AGEMA_reg_buffer_2329_s_current_state_reg ( .D(
        new_AGEMA_signal_3036), .CK(clk), .Q(new_AGEMA_signal_4217) );
  DFF_X1 new_AGEMA_reg_buffer_2332_s_current_state_reg ( .D(Inst_bSbox_T1),
        .CK(clk), .Q(new_AGEMA_signal_4220) );
  DFF_X1 new_AGEMA_reg_buffer_2335_s_current_state_reg ( .D(
        new_AGEMA_signal_2850), .CK(clk), .Q(new_AGEMA_signal_4223) );
  DFF_X1 new_AGEMA_reg_buffer_2338_s_current_state_reg ( .D(Inst_bSbox_T4),
        .CK(clk), .Q(new_AGEMA_signal_4226) );
  DFF_X1 new_AGEMA_reg_buffer_2341_s_current_state_reg ( .D(
        new_AGEMA_signal_2853), .CK(clk), .Q(new_AGEMA_signal_4229) );
  DFF_X1 new_AGEMA_reg_buffer_2344_s_current_state_reg ( .D(Inst_bSbox_T2),
        .CK(clk), .Q(new_AGEMA_signal_4232) );
  DFF_X1 new_AGEMA_reg_buffer_2347_s_current_state_reg ( .D(
        new_AGEMA_signal_2851), .CK(clk), .Q(new_AGEMA_signal_4235) );
  DFF_X1 new_AGEMA_reg_buffer_2350_s_current_state_reg ( .D(ctrl_seq6_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4238) );
  DFF_X1 new_AGEMA_reg_buffer_2354_s_current_state_reg ( .D(ctrl_seq6_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4242) );
  DFF_X1 new_AGEMA_reg_buffer_2358_s_current_state_reg ( .D(ctrl_seq6_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4246) );
  DFF_X1 new_AGEMA_reg_buffer_2362_s_current_state_reg ( .D(ctrl_seq6_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4250) );
  DFF_X1 new_AGEMA_reg_buffer_2366_s_current_state_reg ( .D(ctrl_seq6_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4254) );
  DFF_X1 new_AGEMA_reg_buffer_2370_s_current_state_reg ( .D(ctrl_seq4_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4258) );
  DFF_X1 new_AGEMA_reg_buffer_2374_s_current_state_reg ( .D(ctrl_seq4_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4262) );
  DFF_X1 new_AGEMA_reg_buffer_2378_s_current_state_reg ( .D(ctrl_N14), .CK(clk), .Q(new_AGEMA_signal_4266) );
  DFF_X1 new_AGEMA_reg_buffer_2382_s_current_state_reg ( .D(n250), .CK(clk),
        .Q(new_AGEMA_signal_4270) );
  DFF_X1 new_AGEMA_reg_buffer_2386_s_current_state_reg ( .D(
        stateArray_S00reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4274)
         );
  DFF_X1 new_AGEMA_reg_buffer_2390_s_current_state_reg ( .D(
        new_AGEMA_signal_3126), .CK(clk), .Q(new_AGEMA_signal_4278) );
  DFF_X1 new_AGEMA_reg_buffer_2394_s_current_state_reg ( .D(
        stateArray_S00reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4282)
         );
  DFF_X1 new_AGEMA_reg_buffer_2398_s_current_state_reg ( .D(
        new_AGEMA_signal_3127), .CK(clk), .Q(new_AGEMA_signal_4286) );
  DFF_X1 new_AGEMA_reg_buffer_2402_s_current_state_reg ( .D(
        stateArray_S00reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4290)
         );
  DFF_X1 new_AGEMA_reg_buffer_2406_s_current_state_reg ( .D(
        new_AGEMA_signal_3128), .CK(clk), .Q(new_AGEMA_signal_4294) );
  DFF_X1 new_AGEMA_reg_buffer_2410_s_current_state_reg ( .D(
        stateArray_S00reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4298)
         );
  DFF_X1 new_AGEMA_reg_buffer_2414_s_current_state_reg ( .D(
        new_AGEMA_signal_3129), .CK(clk), .Q(new_AGEMA_signal_4302) );
  DFF_X1 new_AGEMA_reg_buffer_2418_s_current_state_reg ( .D(
        stateArray_S00reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4306)
         );
  DFF_X1 new_AGEMA_reg_buffer_2422_s_current_state_reg ( .D(
        new_AGEMA_signal_3130), .CK(clk), .Q(new_AGEMA_signal_4310) );
  DFF_X1 new_AGEMA_reg_buffer_2426_s_current_state_reg ( .D(
        stateArray_S00reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4314)
         );
  DFF_X1 new_AGEMA_reg_buffer_2430_s_current_state_reg ( .D(
        new_AGEMA_signal_3131), .CK(clk), .Q(new_AGEMA_signal_4318) );
  DFF_X1 new_AGEMA_reg_buffer_2434_s_current_state_reg ( .D(
        stateArray_S00reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4322)
         );
  DFF_X1 new_AGEMA_reg_buffer_2438_s_current_state_reg ( .D(
        new_AGEMA_signal_3132), .CK(clk), .Q(new_AGEMA_signal_4326) );
  DFF_X1 new_AGEMA_reg_buffer_2442_s_current_state_reg ( .D(
        stateArray_S00reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4330)
         );
  DFF_X1 new_AGEMA_reg_buffer_2446_s_current_state_reg ( .D(
        new_AGEMA_signal_3133), .CK(clk), .Q(new_AGEMA_signal_4334) );
  DFF_X1 new_AGEMA_reg_buffer_2450_s_current_state_reg ( .D(
        stateArray_S01reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4338)
         );
  DFF_X1 new_AGEMA_reg_buffer_2454_s_current_state_reg ( .D(
        new_AGEMA_signal_3134), .CK(clk), .Q(new_AGEMA_signal_4342) );
  DFF_X1 new_AGEMA_reg_buffer_2458_s_current_state_reg ( .D(
        stateArray_S01reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4346)
         );
  DFF_X1 new_AGEMA_reg_buffer_2462_s_current_state_reg ( .D(
        new_AGEMA_signal_3135), .CK(clk), .Q(new_AGEMA_signal_4350) );
  DFF_X1 new_AGEMA_reg_buffer_2466_s_current_state_reg ( .D(
        stateArray_S01reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4354)
         );
  DFF_X1 new_AGEMA_reg_buffer_2470_s_current_state_reg ( .D(
        new_AGEMA_signal_3136), .CK(clk), .Q(new_AGEMA_signal_4358) );
  DFF_X1 new_AGEMA_reg_buffer_2474_s_current_state_reg ( .D(
        stateArray_S01reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4362)
         );
  DFF_X1 new_AGEMA_reg_buffer_2478_s_current_state_reg ( .D(
        new_AGEMA_signal_3137), .CK(clk), .Q(new_AGEMA_signal_4366) );
  DFF_X1 new_AGEMA_reg_buffer_2482_s_current_state_reg ( .D(
        stateArray_S01reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4370)
         );
  DFF_X1 new_AGEMA_reg_buffer_2486_s_current_state_reg ( .D(
        new_AGEMA_signal_3138), .CK(clk), .Q(new_AGEMA_signal_4374) );
  DFF_X1 new_AGEMA_reg_buffer_2490_s_current_state_reg ( .D(
        stateArray_S01reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4378)
         );
  DFF_X1 new_AGEMA_reg_buffer_2494_s_current_state_reg ( .D(
        new_AGEMA_signal_3139), .CK(clk), .Q(new_AGEMA_signal_4382) );
  DFF_X1 new_AGEMA_reg_buffer_2498_s_current_state_reg ( .D(
        stateArray_S01reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4386)
         );
  DFF_X1 new_AGEMA_reg_buffer_2502_s_current_state_reg ( .D(
        new_AGEMA_signal_3140), .CK(clk), .Q(new_AGEMA_signal_4390) );
  DFF_X1 new_AGEMA_reg_buffer_2506_s_current_state_reg ( .D(
        stateArray_S01reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4394)
         );
  DFF_X1 new_AGEMA_reg_buffer_2510_s_current_state_reg ( .D(
        new_AGEMA_signal_3141), .CK(clk), .Q(new_AGEMA_signal_4398) );
  DFF_X1 new_AGEMA_reg_buffer_2514_s_current_state_reg ( .D(
        stateArray_S02reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4402)
         );
  DFF_X1 new_AGEMA_reg_buffer_2518_s_current_state_reg ( .D(
        new_AGEMA_signal_3142), .CK(clk), .Q(new_AGEMA_signal_4406) );
  DFF_X1 new_AGEMA_reg_buffer_2522_s_current_state_reg ( .D(
        stateArray_S02reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4410)
         );
  DFF_X1 new_AGEMA_reg_buffer_2526_s_current_state_reg ( .D(
        new_AGEMA_signal_3143), .CK(clk), .Q(new_AGEMA_signal_4414) );
  DFF_X1 new_AGEMA_reg_buffer_2530_s_current_state_reg ( .D(
        stateArray_S02reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4418)
         );
  DFF_X1 new_AGEMA_reg_buffer_2534_s_current_state_reg ( .D(
        new_AGEMA_signal_3144), .CK(clk), .Q(new_AGEMA_signal_4422) );
  DFF_X1 new_AGEMA_reg_buffer_2538_s_current_state_reg ( .D(
        stateArray_S02reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4426)
         );
  DFF_X1 new_AGEMA_reg_buffer_2542_s_current_state_reg ( .D(
        new_AGEMA_signal_3145), .CK(clk), .Q(new_AGEMA_signal_4430) );
  DFF_X1 new_AGEMA_reg_buffer_2546_s_current_state_reg ( .D(
        stateArray_S02reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4434)
         );
  DFF_X1 new_AGEMA_reg_buffer_2550_s_current_state_reg ( .D(
        new_AGEMA_signal_3146), .CK(clk), .Q(new_AGEMA_signal_4438) );
  DFF_X1 new_AGEMA_reg_buffer_2554_s_current_state_reg ( .D(
        stateArray_S02reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4442)
         );
  DFF_X1 new_AGEMA_reg_buffer_2558_s_current_state_reg ( .D(
        new_AGEMA_signal_3147), .CK(clk), .Q(new_AGEMA_signal_4446) );
  DFF_X1 new_AGEMA_reg_buffer_2562_s_current_state_reg ( .D(
        stateArray_S02reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4450)
         );
  DFF_X1 new_AGEMA_reg_buffer_2566_s_current_state_reg ( .D(
        new_AGEMA_signal_3148), .CK(clk), .Q(new_AGEMA_signal_4454) );
  DFF_X1 new_AGEMA_reg_buffer_2570_s_current_state_reg ( .D(
        stateArray_S02reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4458)
         );
  DFF_X1 new_AGEMA_reg_buffer_2574_s_current_state_reg ( .D(
        new_AGEMA_signal_3149), .CK(clk), .Q(new_AGEMA_signal_4462) );
  DFF_X1 new_AGEMA_reg_buffer_2578_s_current_state_reg ( .D(
        stateArray_S03reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4466)
         );
  DFF_X1 new_AGEMA_reg_buffer_2582_s_current_state_reg ( .D(
        new_AGEMA_signal_3150), .CK(clk), .Q(new_AGEMA_signal_4470) );
  DFF_X1 new_AGEMA_reg_buffer_2586_s_current_state_reg ( .D(
        stateArray_S03reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4474)
         );
  DFF_X1 new_AGEMA_reg_buffer_2590_s_current_state_reg ( .D(
        new_AGEMA_signal_3151), .CK(clk), .Q(new_AGEMA_signal_4478) );
  DFF_X1 new_AGEMA_reg_buffer_2594_s_current_state_reg ( .D(
        stateArray_S03reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4482)
         );
  DFF_X1 new_AGEMA_reg_buffer_2598_s_current_state_reg ( .D(
        new_AGEMA_signal_3152), .CK(clk), .Q(new_AGEMA_signal_4486) );
  DFF_X1 new_AGEMA_reg_buffer_2602_s_current_state_reg ( .D(
        stateArray_S03reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4490)
         );
  DFF_X1 new_AGEMA_reg_buffer_2606_s_current_state_reg ( .D(
        new_AGEMA_signal_3153), .CK(clk), .Q(new_AGEMA_signal_4494) );
  DFF_X1 new_AGEMA_reg_buffer_2610_s_current_state_reg ( .D(
        stateArray_S03reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4498)
         );
  DFF_X1 new_AGEMA_reg_buffer_2614_s_current_state_reg ( .D(
        new_AGEMA_signal_3154), .CK(clk), .Q(new_AGEMA_signal_4502) );
  DFF_X1 new_AGEMA_reg_buffer_2618_s_current_state_reg ( .D(
        stateArray_S03reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4506)
         );
  DFF_X1 new_AGEMA_reg_buffer_2622_s_current_state_reg ( .D(
        new_AGEMA_signal_3155), .CK(clk), .Q(new_AGEMA_signal_4510) );
  DFF_X1 new_AGEMA_reg_buffer_2626_s_current_state_reg ( .D(
        stateArray_S03reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4514)
         );
  DFF_X1 new_AGEMA_reg_buffer_2630_s_current_state_reg ( .D(
        new_AGEMA_signal_3156), .CK(clk), .Q(new_AGEMA_signal_4518) );
  DFF_X1 new_AGEMA_reg_buffer_2634_s_current_state_reg ( .D(
        stateArray_S03reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4522)
         );
  DFF_X1 new_AGEMA_reg_buffer_2638_s_current_state_reg ( .D(
        new_AGEMA_signal_3157), .CK(clk), .Q(new_AGEMA_signal_4526) );
  DFF_X1 new_AGEMA_reg_buffer_2642_s_current_state_reg ( .D(
        stateArray_S10reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4530)
         );
  DFF_X1 new_AGEMA_reg_buffer_2646_s_current_state_reg ( .D(
        new_AGEMA_signal_3158), .CK(clk), .Q(new_AGEMA_signal_4534) );
  DFF_X1 new_AGEMA_reg_buffer_2650_s_current_state_reg ( .D(
        stateArray_S10reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4538)
         );
  DFF_X1 new_AGEMA_reg_buffer_2654_s_current_state_reg ( .D(
        new_AGEMA_signal_3159), .CK(clk), .Q(new_AGEMA_signal_4542) );
  DFF_X1 new_AGEMA_reg_buffer_2658_s_current_state_reg ( .D(
        stateArray_S10reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4546)
         );
  DFF_X1 new_AGEMA_reg_buffer_2662_s_current_state_reg ( .D(
        new_AGEMA_signal_3160), .CK(clk), .Q(new_AGEMA_signal_4550) );
  DFF_X1 new_AGEMA_reg_buffer_2666_s_current_state_reg ( .D(
        stateArray_S10reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4554)
         );
  DFF_X1 new_AGEMA_reg_buffer_2670_s_current_state_reg ( .D(
        new_AGEMA_signal_3161), .CK(clk), .Q(new_AGEMA_signal_4558) );
  DFF_X1 new_AGEMA_reg_buffer_2674_s_current_state_reg ( .D(
        stateArray_S10reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4562)
         );
  DFF_X1 new_AGEMA_reg_buffer_2678_s_current_state_reg ( .D(
        new_AGEMA_signal_3162), .CK(clk), .Q(new_AGEMA_signal_4566) );
  DFF_X1 new_AGEMA_reg_buffer_2682_s_current_state_reg ( .D(
        stateArray_S10reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4570)
         );
  DFF_X1 new_AGEMA_reg_buffer_2686_s_current_state_reg ( .D(
        new_AGEMA_signal_3163), .CK(clk), .Q(new_AGEMA_signal_4574) );
  DFF_X1 new_AGEMA_reg_buffer_2690_s_current_state_reg ( .D(
        stateArray_S10reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4578)
         );
  DFF_X1 new_AGEMA_reg_buffer_2694_s_current_state_reg ( .D(
        new_AGEMA_signal_3164), .CK(clk), .Q(new_AGEMA_signal_4582) );
  DFF_X1 new_AGEMA_reg_buffer_2698_s_current_state_reg ( .D(
        stateArray_S10reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4586)
         );
  DFF_X1 new_AGEMA_reg_buffer_2702_s_current_state_reg ( .D(
        new_AGEMA_signal_3165), .CK(clk), .Q(new_AGEMA_signal_4590) );
  DFF_X1 new_AGEMA_reg_buffer_2706_s_current_state_reg ( .D(
        stateArray_S11reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4594)
         );
  DFF_X1 new_AGEMA_reg_buffer_2710_s_current_state_reg ( .D(
        new_AGEMA_signal_3166), .CK(clk), .Q(new_AGEMA_signal_4598) );
  DFF_X1 new_AGEMA_reg_buffer_2714_s_current_state_reg ( .D(
        stateArray_S11reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4602)
         );
  DFF_X1 new_AGEMA_reg_buffer_2718_s_current_state_reg ( .D(
        new_AGEMA_signal_3167), .CK(clk), .Q(new_AGEMA_signal_4606) );
  DFF_X1 new_AGEMA_reg_buffer_2722_s_current_state_reg ( .D(
        stateArray_S11reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4610)
         );
  DFF_X1 new_AGEMA_reg_buffer_2726_s_current_state_reg ( .D(
        new_AGEMA_signal_3168), .CK(clk), .Q(new_AGEMA_signal_4614) );
  DFF_X1 new_AGEMA_reg_buffer_2730_s_current_state_reg ( .D(
        stateArray_S11reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4618)
         );
  DFF_X1 new_AGEMA_reg_buffer_2734_s_current_state_reg ( .D(
        new_AGEMA_signal_3169), .CK(clk), .Q(new_AGEMA_signal_4622) );
  DFF_X1 new_AGEMA_reg_buffer_2738_s_current_state_reg ( .D(
        stateArray_S11reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4626)
         );
  DFF_X1 new_AGEMA_reg_buffer_2742_s_current_state_reg ( .D(
        new_AGEMA_signal_3170), .CK(clk), .Q(new_AGEMA_signal_4630) );
  DFF_X1 new_AGEMA_reg_buffer_2746_s_current_state_reg ( .D(
        stateArray_S11reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4634)
         );
  DFF_X1 new_AGEMA_reg_buffer_2750_s_current_state_reg ( .D(
        new_AGEMA_signal_3171), .CK(clk), .Q(new_AGEMA_signal_4638) );
  DFF_X1 new_AGEMA_reg_buffer_2754_s_current_state_reg ( .D(
        stateArray_S11reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4642)
         );
  DFF_X1 new_AGEMA_reg_buffer_2758_s_current_state_reg ( .D(
        new_AGEMA_signal_3172), .CK(clk), .Q(new_AGEMA_signal_4646) );
  DFF_X1 new_AGEMA_reg_buffer_2762_s_current_state_reg ( .D(
        stateArray_S11reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4650)
         );
  DFF_X1 new_AGEMA_reg_buffer_2766_s_current_state_reg ( .D(
        new_AGEMA_signal_3173), .CK(clk), .Q(new_AGEMA_signal_4654) );
  DFF_X1 new_AGEMA_reg_buffer_2770_s_current_state_reg ( .D(
        stateArray_S12reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4658)
         );
  DFF_X1 new_AGEMA_reg_buffer_2774_s_current_state_reg ( .D(
        new_AGEMA_signal_3174), .CK(clk), .Q(new_AGEMA_signal_4662) );
  DFF_X1 new_AGEMA_reg_buffer_2778_s_current_state_reg ( .D(
        stateArray_S12reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4666)
         );
  DFF_X1 new_AGEMA_reg_buffer_2782_s_current_state_reg ( .D(
        new_AGEMA_signal_3175), .CK(clk), .Q(new_AGEMA_signal_4670) );
  DFF_X1 new_AGEMA_reg_buffer_2786_s_current_state_reg ( .D(
        stateArray_S12reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4674)
         );
  DFF_X1 new_AGEMA_reg_buffer_2790_s_current_state_reg ( .D(
        new_AGEMA_signal_3176), .CK(clk), .Q(new_AGEMA_signal_4678) );
  DFF_X1 new_AGEMA_reg_buffer_2794_s_current_state_reg ( .D(
        stateArray_S12reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4682)
         );
  DFF_X1 new_AGEMA_reg_buffer_2798_s_current_state_reg ( .D(
        new_AGEMA_signal_3177), .CK(clk), .Q(new_AGEMA_signal_4686) );
  DFF_X1 new_AGEMA_reg_buffer_2802_s_current_state_reg ( .D(
        stateArray_S12reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4690)
         );
  DFF_X1 new_AGEMA_reg_buffer_2806_s_current_state_reg ( .D(
        new_AGEMA_signal_3178), .CK(clk), .Q(new_AGEMA_signal_4694) );
  DFF_X1 new_AGEMA_reg_buffer_2810_s_current_state_reg ( .D(
        stateArray_S12reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4698)
         );
  DFF_X1 new_AGEMA_reg_buffer_2814_s_current_state_reg ( .D(
        new_AGEMA_signal_3179), .CK(clk), .Q(new_AGEMA_signal_4702) );
  DFF_X1 new_AGEMA_reg_buffer_2818_s_current_state_reg ( .D(
        stateArray_S12reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4706)
         );
  DFF_X1 new_AGEMA_reg_buffer_2822_s_current_state_reg ( .D(
        new_AGEMA_signal_3180), .CK(clk), .Q(new_AGEMA_signal_4710) );
  DFF_X1 new_AGEMA_reg_buffer_2826_s_current_state_reg ( .D(
        stateArray_S12reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4714)
         );
  DFF_X1 new_AGEMA_reg_buffer_2830_s_current_state_reg ( .D(
        new_AGEMA_signal_3181), .CK(clk), .Q(new_AGEMA_signal_4718) );
  DFF_X1 new_AGEMA_reg_buffer_2834_s_current_state_reg ( .D(
        stateArray_S13reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4722)
         );
  DFF_X1 new_AGEMA_reg_buffer_2838_s_current_state_reg ( .D(
        new_AGEMA_signal_3182), .CK(clk), .Q(new_AGEMA_signal_4726) );
  DFF_X1 new_AGEMA_reg_buffer_2842_s_current_state_reg ( .D(
        stateArray_S13reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4730)
         );
  DFF_X1 new_AGEMA_reg_buffer_2846_s_current_state_reg ( .D(
        new_AGEMA_signal_3183), .CK(clk), .Q(new_AGEMA_signal_4734) );
  DFF_X1 new_AGEMA_reg_buffer_2850_s_current_state_reg ( .D(
        stateArray_S13reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4738)
         );
  DFF_X1 new_AGEMA_reg_buffer_2854_s_current_state_reg ( .D(
        new_AGEMA_signal_3184), .CK(clk), .Q(new_AGEMA_signal_4742) );
  DFF_X1 new_AGEMA_reg_buffer_2858_s_current_state_reg ( .D(
        stateArray_S13reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4746)
         );
  DFF_X1 new_AGEMA_reg_buffer_2862_s_current_state_reg ( .D(
        new_AGEMA_signal_3185), .CK(clk), .Q(new_AGEMA_signal_4750) );
  DFF_X1 new_AGEMA_reg_buffer_2866_s_current_state_reg ( .D(
        stateArray_S13reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4754)
         );
  DFF_X1 new_AGEMA_reg_buffer_2870_s_current_state_reg ( .D(
        new_AGEMA_signal_3186), .CK(clk), .Q(new_AGEMA_signal_4758) );
  DFF_X1 new_AGEMA_reg_buffer_2874_s_current_state_reg ( .D(
        stateArray_S13reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4762)
         );
  DFF_X1 new_AGEMA_reg_buffer_2878_s_current_state_reg ( .D(
        new_AGEMA_signal_3187), .CK(clk), .Q(new_AGEMA_signal_4766) );
  DFF_X1 new_AGEMA_reg_buffer_2882_s_current_state_reg ( .D(
        stateArray_S13reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4770)
         );
  DFF_X1 new_AGEMA_reg_buffer_2886_s_current_state_reg ( .D(
        new_AGEMA_signal_3188), .CK(clk), .Q(new_AGEMA_signal_4774) );
  DFF_X1 new_AGEMA_reg_buffer_2890_s_current_state_reg ( .D(
        stateArray_S13reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4778)
         );
  DFF_X1 new_AGEMA_reg_buffer_2894_s_current_state_reg ( .D(
        new_AGEMA_signal_3189), .CK(clk), .Q(new_AGEMA_signal_4782) );
  DFF_X1 new_AGEMA_reg_buffer_2898_s_current_state_reg ( .D(
        stateArray_S20reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4786)
         );
  DFF_X1 new_AGEMA_reg_buffer_2902_s_current_state_reg ( .D(
        new_AGEMA_signal_3190), .CK(clk), .Q(new_AGEMA_signal_4790) );
  DFF_X1 new_AGEMA_reg_buffer_2906_s_current_state_reg ( .D(
        stateArray_S20reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4794)
         );
  DFF_X1 new_AGEMA_reg_buffer_2910_s_current_state_reg ( .D(
        new_AGEMA_signal_3191), .CK(clk), .Q(new_AGEMA_signal_4798) );
  DFF_X1 new_AGEMA_reg_buffer_2914_s_current_state_reg ( .D(
        stateArray_S20reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4802)
         );
  DFF_X1 new_AGEMA_reg_buffer_2918_s_current_state_reg ( .D(
        new_AGEMA_signal_3192), .CK(clk), .Q(new_AGEMA_signal_4806) );
  DFF_X1 new_AGEMA_reg_buffer_2922_s_current_state_reg ( .D(
        stateArray_S20reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4810)
         );
  DFF_X1 new_AGEMA_reg_buffer_2926_s_current_state_reg ( .D(
        new_AGEMA_signal_3193), .CK(clk), .Q(new_AGEMA_signal_4814) );
  DFF_X1 new_AGEMA_reg_buffer_2930_s_current_state_reg ( .D(
        stateArray_S20reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4818)
         );
  DFF_X1 new_AGEMA_reg_buffer_2934_s_current_state_reg ( .D(
        new_AGEMA_signal_3194), .CK(clk), .Q(new_AGEMA_signal_4822) );
  DFF_X1 new_AGEMA_reg_buffer_2938_s_current_state_reg ( .D(
        stateArray_S20reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4826)
         );
  DFF_X1 new_AGEMA_reg_buffer_2942_s_current_state_reg ( .D(
        new_AGEMA_signal_3195), .CK(clk), .Q(new_AGEMA_signal_4830) );
  DFF_X1 new_AGEMA_reg_buffer_2946_s_current_state_reg ( .D(
        stateArray_S20reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4834)
         );
  DFF_X1 new_AGEMA_reg_buffer_2950_s_current_state_reg ( .D(
        new_AGEMA_signal_3196), .CK(clk), .Q(new_AGEMA_signal_4838) );
  DFF_X1 new_AGEMA_reg_buffer_2954_s_current_state_reg ( .D(
        stateArray_S20reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4842)
         );
  DFF_X1 new_AGEMA_reg_buffer_2958_s_current_state_reg ( .D(
        new_AGEMA_signal_3197), .CK(clk), .Q(new_AGEMA_signal_4846) );
  DFF_X1 new_AGEMA_reg_buffer_2962_s_current_state_reg ( .D(
        stateArray_S21reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4850)
         );
  DFF_X1 new_AGEMA_reg_buffer_2966_s_current_state_reg ( .D(
        new_AGEMA_signal_3198), .CK(clk), .Q(new_AGEMA_signal_4854) );
  DFF_X1 new_AGEMA_reg_buffer_2970_s_current_state_reg ( .D(
        stateArray_S21reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4858)
         );
  DFF_X1 new_AGEMA_reg_buffer_2974_s_current_state_reg ( .D(
        new_AGEMA_signal_3199), .CK(clk), .Q(new_AGEMA_signal_4862) );
  DFF_X1 new_AGEMA_reg_buffer_2978_s_current_state_reg ( .D(
        stateArray_S21reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4866)
         );
  DFF_X1 new_AGEMA_reg_buffer_2982_s_current_state_reg ( .D(
        new_AGEMA_signal_3200), .CK(clk), .Q(new_AGEMA_signal_4870) );
  DFF_X1 new_AGEMA_reg_buffer_2986_s_current_state_reg ( .D(
        stateArray_S21reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4874)
         );
  DFF_X1 new_AGEMA_reg_buffer_2990_s_current_state_reg ( .D(
        new_AGEMA_signal_3201), .CK(clk), .Q(new_AGEMA_signal_4878) );
  DFF_X1 new_AGEMA_reg_buffer_2994_s_current_state_reg ( .D(
        stateArray_S21reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4882)
         );
  DFF_X1 new_AGEMA_reg_buffer_2998_s_current_state_reg ( .D(
        new_AGEMA_signal_3202), .CK(clk), .Q(new_AGEMA_signal_4886) );
  DFF_X1 new_AGEMA_reg_buffer_3002_s_current_state_reg ( .D(
        stateArray_S21reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4890)
         );
  DFF_X1 new_AGEMA_reg_buffer_3006_s_current_state_reg ( .D(
        new_AGEMA_signal_3203), .CK(clk), .Q(new_AGEMA_signal_4894) );
  DFF_X1 new_AGEMA_reg_buffer_3010_s_current_state_reg ( .D(
        stateArray_S21reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4898)
         );
  DFF_X1 new_AGEMA_reg_buffer_3014_s_current_state_reg ( .D(
        new_AGEMA_signal_3204), .CK(clk), .Q(new_AGEMA_signal_4902) );
  DFF_X1 new_AGEMA_reg_buffer_3018_s_current_state_reg ( .D(
        stateArray_S21reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4906)
         );
  DFF_X1 new_AGEMA_reg_buffer_3022_s_current_state_reg ( .D(
        new_AGEMA_signal_3205), .CK(clk), .Q(new_AGEMA_signal_4910) );
  DFF_X1 new_AGEMA_reg_buffer_3026_s_current_state_reg ( .D(
        stateArray_S22reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4914)
         );
  DFF_X1 new_AGEMA_reg_buffer_3030_s_current_state_reg ( .D(
        new_AGEMA_signal_3206), .CK(clk), .Q(new_AGEMA_signal_4918) );
  DFF_X1 new_AGEMA_reg_buffer_3034_s_current_state_reg ( .D(
        stateArray_S22reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4922)
         );
  DFF_X1 new_AGEMA_reg_buffer_3038_s_current_state_reg ( .D(
        new_AGEMA_signal_3207), .CK(clk), .Q(new_AGEMA_signal_4926) );
  DFF_X1 new_AGEMA_reg_buffer_3042_s_current_state_reg ( .D(
        stateArray_S22reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4930)
         );
  DFF_X1 new_AGEMA_reg_buffer_3046_s_current_state_reg ( .D(
        new_AGEMA_signal_3208), .CK(clk), .Q(new_AGEMA_signal_4934) );
  DFF_X1 new_AGEMA_reg_buffer_3050_s_current_state_reg ( .D(
        stateArray_S22reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_4938)
         );
  DFF_X1 new_AGEMA_reg_buffer_3054_s_current_state_reg ( .D(
        new_AGEMA_signal_3209), .CK(clk), .Q(new_AGEMA_signal_4942) );
  DFF_X1 new_AGEMA_reg_buffer_3058_s_current_state_reg ( .D(
        stateArray_S22reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_4946)
         );
  DFF_X1 new_AGEMA_reg_buffer_3062_s_current_state_reg ( .D(
        new_AGEMA_signal_3210), .CK(clk), .Q(new_AGEMA_signal_4950) );
  DFF_X1 new_AGEMA_reg_buffer_3066_s_current_state_reg ( .D(
        stateArray_S22reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_4954)
         );
  DFF_X1 new_AGEMA_reg_buffer_3070_s_current_state_reg ( .D(
        new_AGEMA_signal_3211), .CK(clk), .Q(new_AGEMA_signal_4958) );
  DFF_X1 new_AGEMA_reg_buffer_3074_s_current_state_reg ( .D(
        stateArray_S22reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_4962)
         );
  DFF_X1 new_AGEMA_reg_buffer_3078_s_current_state_reg ( .D(
        new_AGEMA_signal_3212), .CK(clk), .Q(new_AGEMA_signal_4966) );
  DFF_X1 new_AGEMA_reg_buffer_3082_s_current_state_reg ( .D(
        stateArray_S22reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_4970)
         );
  DFF_X1 new_AGEMA_reg_buffer_3086_s_current_state_reg ( .D(
        new_AGEMA_signal_3213), .CK(clk), .Q(new_AGEMA_signal_4974) );
  DFF_X1 new_AGEMA_reg_buffer_3090_s_current_state_reg ( .D(
        stateArray_S23reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_4978)
         );
  DFF_X1 new_AGEMA_reg_buffer_3094_s_current_state_reg ( .D(
        new_AGEMA_signal_3214), .CK(clk), .Q(new_AGEMA_signal_4982) );
  DFF_X1 new_AGEMA_reg_buffer_3098_s_current_state_reg ( .D(
        stateArray_S23reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_4986)
         );
  DFF_X1 new_AGEMA_reg_buffer_3102_s_current_state_reg ( .D(
        new_AGEMA_signal_3215), .CK(clk), .Q(new_AGEMA_signal_4990) );
  DFF_X1 new_AGEMA_reg_buffer_3106_s_current_state_reg ( .D(
        stateArray_S23reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_4994)
         );
  DFF_X1 new_AGEMA_reg_buffer_3110_s_current_state_reg ( .D(
        new_AGEMA_signal_3216), .CK(clk), .Q(new_AGEMA_signal_4998) );
  DFF_X1 new_AGEMA_reg_buffer_3114_s_current_state_reg ( .D(
        stateArray_S23reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_5002)
         );
  DFF_X1 new_AGEMA_reg_buffer_3118_s_current_state_reg ( .D(
        new_AGEMA_signal_3217), .CK(clk), .Q(new_AGEMA_signal_5006) );
  DFF_X1 new_AGEMA_reg_buffer_3122_s_current_state_reg ( .D(
        stateArray_S23reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_5010)
         );
  DFF_X1 new_AGEMA_reg_buffer_3126_s_current_state_reg ( .D(
        new_AGEMA_signal_3218), .CK(clk), .Q(new_AGEMA_signal_5014) );
  DFF_X1 new_AGEMA_reg_buffer_3130_s_current_state_reg ( .D(
        stateArray_S23reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_5018)
         );
  DFF_X1 new_AGEMA_reg_buffer_3134_s_current_state_reg ( .D(
        new_AGEMA_signal_3219), .CK(clk), .Q(new_AGEMA_signal_5022) );
  DFF_X1 new_AGEMA_reg_buffer_3138_s_current_state_reg ( .D(
        stateArray_S23reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_5026)
         );
  DFF_X1 new_AGEMA_reg_buffer_3142_s_current_state_reg ( .D(
        new_AGEMA_signal_3220), .CK(clk), .Q(new_AGEMA_signal_5030) );
  DFF_X1 new_AGEMA_reg_buffer_3146_s_current_state_reg ( .D(
        stateArray_S23reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_5034)
         );
  DFF_X1 new_AGEMA_reg_buffer_3150_s_current_state_reg ( .D(
        new_AGEMA_signal_3221), .CK(clk), .Q(new_AGEMA_signal_5038) );
  DFF_X1 new_AGEMA_reg_buffer_3154_s_current_state_reg ( .D(
        stateArray_S30reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_5042)
         );
  DFF_X1 new_AGEMA_reg_buffer_3158_s_current_state_reg ( .D(
        new_AGEMA_signal_3222), .CK(clk), .Q(new_AGEMA_signal_5046) );
  DFF_X1 new_AGEMA_reg_buffer_3162_s_current_state_reg ( .D(
        stateArray_S30reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_5050)
         );
  DFF_X1 new_AGEMA_reg_buffer_3166_s_current_state_reg ( .D(
        new_AGEMA_signal_3223), .CK(clk), .Q(new_AGEMA_signal_5054) );
  DFF_X1 new_AGEMA_reg_buffer_3170_s_current_state_reg ( .D(
        stateArray_S30reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_5058)
         );
  DFF_X1 new_AGEMA_reg_buffer_3174_s_current_state_reg ( .D(
        new_AGEMA_signal_3224), .CK(clk), .Q(new_AGEMA_signal_5062) );
  DFF_X1 new_AGEMA_reg_buffer_3178_s_current_state_reg ( .D(
        stateArray_S30reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_5066)
         );
  DFF_X1 new_AGEMA_reg_buffer_3182_s_current_state_reg ( .D(
        new_AGEMA_signal_3225), .CK(clk), .Q(new_AGEMA_signal_5070) );
  DFF_X1 new_AGEMA_reg_buffer_3186_s_current_state_reg ( .D(
        stateArray_S30reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_5074)
         );
  DFF_X1 new_AGEMA_reg_buffer_3190_s_current_state_reg ( .D(
        new_AGEMA_signal_3226), .CK(clk), .Q(new_AGEMA_signal_5078) );
  DFF_X1 new_AGEMA_reg_buffer_3194_s_current_state_reg ( .D(
        stateArray_S30reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_5082)
         );
  DFF_X1 new_AGEMA_reg_buffer_3198_s_current_state_reg ( .D(
        new_AGEMA_signal_3227), .CK(clk), .Q(new_AGEMA_signal_5086) );
  DFF_X1 new_AGEMA_reg_buffer_3202_s_current_state_reg ( .D(
        stateArray_S30reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_5090)
         );
  DFF_X1 new_AGEMA_reg_buffer_3206_s_current_state_reg ( .D(
        new_AGEMA_signal_3228), .CK(clk), .Q(new_AGEMA_signal_5094) );
  DFF_X1 new_AGEMA_reg_buffer_3210_s_current_state_reg ( .D(
        stateArray_S30reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_5098)
         );
  DFF_X1 new_AGEMA_reg_buffer_3214_s_current_state_reg ( .D(
        new_AGEMA_signal_3229), .CK(clk), .Q(new_AGEMA_signal_5102) );
  DFF_X1 new_AGEMA_reg_buffer_3218_s_current_state_reg ( .D(
        stateArray_S31reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_5106)
         );
  DFF_X1 new_AGEMA_reg_buffer_3222_s_current_state_reg ( .D(
        new_AGEMA_signal_3230), .CK(clk), .Q(new_AGEMA_signal_5110) );
  DFF_X1 new_AGEMA_reg_buffer_3226_s_current_state_reg ( .D(
        stateArray_S31reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_5114)
         );
  DFF_X1 new_AGEMA_reg_buffer_3230_s_current_state_reg ( .D(
        new_AGEMA_signal_3231), .CK(clk), .Q(new_AGEMA_signal_5118) );
  DFF_X1 new_AGEMA_reg_buffer_3234_s_current_state_reg ( .D(
        stateArray_S31reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_5122)
         );
  DFF_X1 new_AGEMA_reg_buffer_3238_s_current_state_reg ( .D(
        new_AGEMA_signal_3232), .CK(clk), .Q(new_AGEMA_signal_5126) );
  DFF_X1 new_AGEMA_reg_buffer_3242_s_current_state_reg ( .D(
        stateArray_S31reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_5130)
         );
  DFF_X1 new_AGEMA_reg_buffer_3246_s_current_state_reg ( .D(
        new_AGEMA_signal_3233), .CK(clk), .Q(new_AGEMA_signal_5134) );
  DFF_X1 new_AGEMA_reg_buffer_3250_s_current_state_reg ( .D(
        stateArray_S31reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_5138)
         );
  DFF_X1 new_AGEMA_reg_buffer_3254_s_current_state_reg ( .D(
        new_AGEMA_signal_3234), .CK(clk), .Q(new_AGEMA_signal_5142) );
  DFF_X1 new_AGEMA_reg_buffer_3258_s_current_state_reg ( .D(
        stateArray_S31reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_5146)
         );
  DFF_X1 new_AGEMA_reg_buffer_3262_s_current_state_reg ( .D(
        new_AGEMA_signal_3235), .CK(clk), .Q(new_AGEMA_signal_5150) );
  DFF_X1 new_AGEMA_reg_buffer_3266_s_current_state_reg ( .D(
        stateArray_S31reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_5154)
         );
  DFF_X1 new_AGEMA_reg_buffer_3270_s_current_state_reg ( .D(
        new_AGEMA_signal_3236), .CK(clk), .Q(new_AGEMA_signal_5158) );
  DFF_X1 new_AGEMA_reg_buffer_3274_s_current_state_reg ( .D(
        stateArray_S31reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_5162)
         );
  DFF_X1 new_AGEMA_reg_buffer_3278_s_current_state_reg ( .D(
        new_AGEMA_signal_3237), .CK(clk), .Q(new_AGEMA_signal_5166) );
  DFF_X1 new_AGEMA_reg_buffer_3282_s_current_state_reg ( .D(
        stateArray_S32reg_gff_1_SFF_0_QD), .CK(clk), .Q(new_AGEMA_signal_5170)
         );
  DFF_X1 new_AGEMA_reg_buffer_3286_s_current_state_reg ( .D(
        new_AGEMA_signal_3238), .CK(clk), .Q(new_AGEMA_signal_5174) );
  DFF_X1 new_AGEMA_reg_buffer_3290_s_current_state_reg ( .D(
        stateArray_S32reg_gff_1_SFF_1_QD), .CK(clk), .Q(new_AGEMA_signal_5178)
         );
  DFF_X1 new_AGEMA_reg_buffer_3294_s_current_state_reg ( .D(
        new_AGEMA_signal_3239), .CK(clk), .Q(new_AGEMA_signal_5182) );
  DFF_X1 new_AGEMA_reg_buffer_3298_s_current_state_reg ( .D(
        stateArray_S32reg_gff_1_SFF_2_QD), .CK(clk), .Q(new_AGEMA_signal_5186)
         );
  DFF_X1 new_AGEMA_reg_buffer_3302_s_current_state_reg ( .D(
        new_AGEMA_signal_3240), .CK(clk), .Q(new_AGEMA_signal_5190) );
  DFF_X1 new_AGEMA_reg_buffer_3306_s_current_state_reg ( .D(
        stateArray_S32reg_gff_1_SFF_3_QD), .CK(clk), .Q(new_AGEMA_signal_5194)
         );
  DFF_X1 new_AGEMA_reg_buffer_3310_s_current_state_reg ( .D(
        new_AGEMA_signal_3241), .CK(clk), .Q(new_AGEMA_signal_5198) );
  DFF_X1 new_AGEMA_reg_buffer_3314_s_current_state_reg ( .D(
        stateArray_S32reg_gff_1_SFF_4_QD), .CK(clk), .Q(new_AGEMA_signal_5202)
         );
  DFF_X1 new_AGEMA_reg_buffer_3318_s_current_state_reg ( .D(
        new_AGEMA_signal_3242), .CK(clk), .Q(new_AGEMA_signal_5206) );
  DFF_X1 new_AGEMA_reg_buffer_3322_s_current_state_reg ( .D(
        stateArray_S32reg_gff_1_SFF_5_QD), .CK(clk), .Q(new_AGEMA_signal_5210)
         );
  DFF_X1 new_AGEMA_reg_buffer_3326_s_current_state_reg ( .D(
        new_AGEMA_signal_3243), .CK(clk), .Q(new_AGEMA_signal_5214) );
  DFF_X1 new_AGEMA_reg_buffer_3330_s_current_state_reg ( .D(
        stateArray_S32reg_gff_1_SFF_6_QD), .CK(clk), .Q(new_AGEMA_signal_5218)
         );
  DFF_X1 new_AGEMA_reg_buffer_3334_s_current_state_reg ( .D(
        new_AGEMA_signal_3244), .CK(clk), .Q(new_AGEMA_signal_5222) );
  DFF_X1 new_AGEMA_reg_buffer_3338_s_current_state_reg ( .D(
        stateArray_S32reg_gff_1_SFF_7_QD), .CK(clk), .Q(new_AGEMA_signal_5226)
         );
  DFF_X1 new_AGEMA_reg_buffer_3342_s_current_state_reg ( .D(
        new_AGEMA_signal_3245), .CK(clk), .Q(new_AGEMA_signal_5230) );
  DFF_X1 new_AGEMA_reg_buffer_3346_s_current_state_reg ( .D(
        KeyArray_S00reg_gff_1_SFF_0_n5), .CK(clk), .Q(new_AGEMA_signal_5234)
         );
  DFF_X1 new_AGEMA_reg_buffer_3350_s_current_state_reg ( .D(
        new_AGEMA_signal_3375), .CK(clk), .Q(new_AGEMA_signal_5238) );
  DFF_X1 new_AGEMA_reg_buffer_3354_s_current_state_reg ( .D(
        KeyArray_S00reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_5242)
         );
  DFF_X1 new_AGEMA_reg_buffer_3358_s_current_state_reg ( .D(
        new_AGEMA_signal_3376), .CK(clk), .Q(new_AGEMA_signal_5246) );
  DFF_X1 new_AGEMA_reg_buffer_3362_s_current_state_reg ( .D(
        KeyArray_S00reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_5250)
         );
  DFF_X1 new_AGEMA_reg_buffer_3366_s_current_state_reg ( .D(
        new_AGEMA_signal_3377), .CK(clk), .Q(new_AGEMA_signal_5254) );
  DFF_X1 new_AGEMA_reg_buffer_3370_s_current_state_reg ( .D(
        KeyArray_S00reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_5258)
         );
  DFF_X1 new_AGEMA_reg_buffer_3374_s_current_state_reg ( .D(
        new_AGEMA_signal_3378), .CK(clk), .Q(new_AGEMA_signal_5262) );
  DFF_X1 new_AGEMA_reg_buffer_3378_s_current_state_reg ( .D(
        KeyArray_S00reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_5266)
         );
  DFF_X1 new_AGEMA_reg_buffer_3382_s_current_state_reg ( .D(
        new_AGEMA_signal_3379), .CK(clk), .Q(new_AGEMA_signal_5270) );
  DFF_X1 new_AGEMA_reg_buffer_3386_s_current_state_reg ( .D(
        KeyArray_S00reg_gff_1_SFF_5_n6), .CK(clk), .Q(new_AGEMA_signal_5274)
         );
  DFF_X1 new_AGEMA_reg_buffer_3390_s_current_state_reg ( .D(
        new_AGEMA_signal_3380), .CK(clk), .Q(new_AGEMA_signal_5278) );
  DFF_X1 new_AGEMA_reg_buffer_3394_s_current_state_reg ( .D(
        KeyArray_S00reg_gff_1_SFF_6_n6), .CK(clk), .Q(new_AGEMA_signal_5282)
         );
  DFF_X1 new_AGEMA_reg_buffer_3398_s_current_state_reg ( .D(
        new_AGEMA_signal_3381), .CK(clk), .Q(new_AGEMA_signal_5286) );
  DFF_X1 new_AGEMA_reg_buffer_3402_s_current_state_reg ( .D(
        KeyArray_S00reg_gff_1_SFF_7_n6), .CK(clk), .Q(new_AGEMA_signal_5290)
         );
  DFF_X1 new_AGEMA_reg_buffer_3406_s_current_state_reg ( .D(
        new_AGEMA_signal_3382), .CK(clk), .Q(new_AGEMA_signal_5294) );
  DFF_X1 new_AGEMA_reg_buffer_3410_s_current_state_reg ( .D(
        KeyArray_S01reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_5298)
         );
  DFF_X1 new_AGEMA_reg_buffer_3414_s_current_state_reg ( .D(
        new_AGEMA_signal_3275), .CK(clk), .Q(new_AGEMA_signal_5302) );
  DFF_X1 new_AGEMA_reg_buffer_3418_s_current_state_reg ( .D(
        KeyArray_S01reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_5306)
         );
  DFF_X1 new_AGEMA_reg_buffer_3422_s_current_state_reg ( .D(
        new_AGEMA_signal_3276), .CK(clk), .Q(new_AGEMA_signal_5310) );
  DFF_X1 new_AGEMA_reg_buffer_3426_s_current_state_reg ( .D(
        KeyArray_S01reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_5314)
         );
  DFF_X1 new_AGEMA_reg_buffer_3430_s_current_state_reg ( .D(
        new_AGEMA_signal_3277), .CK(clk), .Q(new_AGEMA_signal_5318) );
  DFF_X1 new_AGEMA_reg_buffer_3434_s_current_state_reg ( .D(
        KeyArray_S01reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_5322)
         );
  DFF_X1 new_AGEMA_reg_buffer_3438_s_current_state_reg ( .D(
        new_AGEMA_signal_3278), .CK(clk), .Q(new_AGEMA_signal_5326) );
  DFF_X1 new_AGEMA_reg_buffer_3442_s_current_state_reg ( .D(
        KeyArray_S01reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_5330)
         );
  DFF_X1 new_AGEMA_reg_buffer_3446_s_current_state_reg ( .D(
        new_AGEMA_signal_3279), .CK(clk), .Q(new_AGEMA_signal_5334) );
  DFF_X1 new_AGEMA_reg_buffer_3450_s_current_state_reg ( .D(
        KeyArray_S01reg_gff_1_SFF_5_n6), .CK(clk), .Q(new_AGEMA_signal_5338)
         );
  DFF_X1 new_AGEMA_reg_buffer_3454_s_current_state_reg ( .D(
        new_AGEMA_signal_3280), .CK(clk), .Q(new_AGEMA_signal_5342) );
  DFF_X1 new_AGEMA_reg_buffer_3458_s_current_state_reg ( .D(
        KeyArray_S01reg_gff_1_SFF_6_n6), .CK(clk), .Q(new_AGEMA_signal_5346)
         );
  DFF_X1 new_AGEMA_reg_buffer_3462_s_current_state_reg ( .D(
        new_AGEMA_signal_3281), .CK(clk), .Q(new_AGEMA_signal_5350) );
  DFF_X1 new_AGEMA_reg_buffer_3466_s_current_state_reg ( .D(
        KeyArray_S01reg_gff_1_SFF_7_n6), .CK(clk), .Q(new_AGEMA_signal_5354)
         );
  DFF_X1 new_AGEMA_reg_buffer_3470_s_current_state_reg ( .D(
        new_AGEMA_signal_3282), .CK(clk), .Q(new_AGEMA_signal_5358) );
  DFF_X1 new_AGEMA_reg_buffer_3474_s_current_state_reg ( .D(
        KeyArray_S02reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_5362)
         );
  DFF_X1 new_AGEMA_reg_buffer_3478_s_current_state_reg ( .D(
        new_AGEMA_signal_3283), .CK(clk), .Q(new_AGEMA_signal_5366) );
  DFF_X1 new_AGEMA_reg_buffer_3482_s_current_state_reg ( .D(
        KeyArray_S02reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_5370)
         );
  DFF_X1 new_AGEMA_reg_buffer_3486_s_current_state_reg ( .D(
        new_AGEMA_signal_3284), .CK(clk), .Q(new_AGEMA_signal_5374) );
  DFF_X1 new_AGEMA_reg_buffer_3490_s_current_state_reg ( .D(
        KeyArray_S02reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_5378)
         );
  DFF_X1 new_AGEMA_reg_buffer_3494_s_current_state_reg ( .D(
        new_AGEMA_signal_3285), .CK(clk), .Q(new_AGEMA_signal_5382) );
  DFF_X1 new_AGEMA_reg_buffer_3498_s_current_state_reg ( .D(
        KeyArray_S02reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_5386)
         );
  DFF_X1 new_AGEMA_reg_buffer_3502_s_current_state_reg ( .D(
        new_AGEMA_signal_3286), .CK(clk), .Q(new_AGEMA_signal_5390) );
  DFF_X1 new_AGEMA_reg_buffer_3506_s_current_state_reg ( .D(
        KeyArray_S02reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_5394)
         );
  DFF_X1 new_AGEMA_reg_buffer_3510_s_current_state_reg ( .D(
        new_AGEMA_signal_3287), .CK(clk), .Q(new_AGEMA_signal_5398) );
  DFF_X1 new_AGEMA_reg_buffer_3514_s_current_state_reg ( .D(
        KeyArray_S02reg_gff_1_SFF_5_n6), .CK(clk), .Q(new_AGEMA_signal_5402)
         );
  DFF_X1 new_AGEMA_reg_buffer_3518_s_current_state_reg ( .D(
        new_AGEMA_signal_3288), .CK(clk), .Q(new_AGEMA_signal_5406) );
  DFF_X1 new_AGEMA_reg_buffer_3522_s_current_state_reg ( .D(
        KeyArray_S02reg_gff_1_SFF_6_n6), .CK(clk), .Q(new_AGEMA_signal_5410)
         );
  DFF_X1 new_AGEMA_reg_buffer_3526_s_current_state_reg ( .D(
        new_AGEMA_signal_3289), .CK(clk), .Q(new_AGEMA_signal_5414) );
  DFF_X1 new_AGEMA_reg_buffer_3530_s_current_state_reg ( .D(
        KeyArray_S02reg_gff_1_SFF_7_n6), .CK(clk), .Q(new_AGEMA_signal_5418)
         );
  DFF_X1 new_AGEMA_reg_buffer_3534_s_current_state_reg ( .D(
        new_AGEMA_signal_3290), .CK(clk), .Q(new_AGEMA_signal_5422) );
  DFF_X1 new_AGEMA_reg_buffer_3538_s_current_state_reg ( .D(
        KeyArray_S03reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_5426)
         );
  DFF_X1 new_AGEMA_reg_buffer_3542_s_current_state_reg ( .D(
        new_AGEMA_signal_3291), .CK(clk), .Q(new_AGEMA_signal_5430) );
  DFF_X1 new_AGEMA_reg_buffer_3546_s_current_state_reg ( .D(
        KeyArray_S03reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_5434)
         );
  DFF_X1 new_AGEMA_reg_buffer_3550_s_current_state_reg ( .D(
        new_AGEMA_signal_3292), .CK(clk), .Q(new_AGEMA_signal_5438) );
  DFF_X1 new_AGEMA_reg_buffer_3554_s_current_state_reg ( .D(
        KeyArray_S03reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_5442)
         );
  DFF_X1 new_AGEMA_reg_buffer_3558_s_current_state_reg ( .D(
        new_AGEMA_signal_3293), .CK(clk), .Q(new_AGEMA_signal_5446) );
  DFF_X1 new_AGEMA_reg_buffer_3562_s_current_state_reg ( .D(
        KeyArray_S03reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_5450)
         );
  DFF_X1 new_AGEMA_reg_buffer_3566_s_current_state_reg ( .D(
        new_AGEMA_signal_3294), .CK(clk), .Q(new_AGEMA_signal_5454) );
  DFF_X1 new_AGEMA_reg_buffer_3570_s_current_state_reg ( .D(
        KeyArray_S03reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_5458)
         );
  DFF_X1 new_AGEMA_reg_buffer_3574_s_current_state_reg ( .D(
        new_AGEMA_signal_3295), .CK(clk), .Q(new_AGEMA_signal_5462) );
  DFF_X1 new_AGEMA_reg_buffer_3578_s_current_state_reg ( .D(
        KeyArray_S03reg_gff_1_SFF_5_n5), .CK(clk), .Q(new_AGEMA_signal_5466)
         );
  DFF_X1 new_AGEMA_reg_buffer_3582_s_current_state_reg ( .D(
        new_AGEMA_signal_3296), .CK(clk), .Q(new_AGEMA_signal_5470) );
  DFF_X1 new_AGEMA_reg_buffer_3586_s_current_state_reg ( .D(
        KeyArray_S03reg_gff_1_SFF_6_n5), .CK(clk), .Q(new_AGEMA_signal_5474)
         );
  DFF_X1 new_AGEMA_reg_buffer_3590_s_current_state_reg ( .D(
        new_AGEMA_signal_3297), .CK(clk), .Q(new_AGEMA_signal_5478) );
  DFF_X1 new_AGEMA_reg_buffer_3594_s_current_state_reg ( .D(
        KeyArray_S03reg_gff_1_SFF_7_n5), .CK(clk), .Q(new_AGEMA_signal_5482)
         );
  DFF_X1 new_AGEMA_reg_buffer_3598_s_current_state_reg ( .D(
        new_AGEMA_signal_3298), .CK(clk), .Q(new_AGEMA_signal_5486) );
  DFF_X1 new_AGEMA_reg_buffer_3602_s_current_state_reg ( .D(
        KeyArray_S10reg_gff_1_SFF_0_n5), .CK(clk), .Q(new_AGEMA_signal_5490)
         );
  DFF_X1 new_AGEMA_reg_buffer_3606_s_current_state_reg ( .D(
        new_AGEMA_signal_3299), .CK(clk), .Q(new_AGEMA_signal_5494) );
  DFF_X1 new_AGEMA_reg_buffer_3610_s_current_state_reg ( .D(
        KeyArray_S10reg_gff_1_SFF_1_n5), .CK(clk), .Q(new_AGEMA_signal_5498)
         );
  DFF_X1 new_AGEMA_reg_buffer_3614_s_current_state_reg ( .D(
        new_AGEMA_signal_3300), .CK(clk), .Q(new_AGEMA_signal_5502) );
  DFF_X1 new_AGEMA_reg_buffer_3618_s_current_state_reg ( .D(
        KeyArray_S10reg_gff_1_SFF_2_n5), .CK(clk), .Q(new_AGEMA_signal_5506)
         );
  DFF_X1 new_AGEMA_reg_buffer_3622_s_current_state_reg ( .D(
        new_AGEMA_signal_3301), .CK(clk), .Q(new_AGEMA_signal_5510) );
  DFF_X1 new_AGEMA_reg_buffer_3626_s_current_state_reg ( .D(
        KeyArray_S10reg_gff_1_SFF_3_n5), .CK(clk), .Q(new_AGEMA_signal_5514)
         );
  DFF_X1 new_AGEMA_reg_buffer_3630_s_current_state_reg ( .D(
        new_AGEMA_signal_3302), .CK(clk), .Q(new_AGEMA_signal_5518) );
  DFF_X1 new_AGEMA_reg_buffer_3634_s_current_state_reg ( .D(
        KeyArray_S10reg_gff_1_SFF_4_n5), .CK(clk), .Q(new_AGEMA_signal_5522)
         );
  DFF_X1 new_AGEMA_reg_buffer_3638_s_current_state_reg ( .D(
        new_AGEMA_signal_3303), .CK(clk), .Q(new_AGEMA_signal_5526) );
  DFF_X1 new_AGEMA_reg_buffer_3642_s_current_state_reg ( .D(
        KeyArray_S10reg_gff_1_SFF_5_n5), .CK(clk), .Q(new_AGEMA_signal_5530)
         );
  DFF_X1 new_AGEMA_reg_buffer_3646_s_current_state_reg ( .D(
        new_AGEMA_signal_3304), .CK(clk), .Q(new_AGEMA_signal_5534) );
  DFF_X1 new_AGEMA_reg_buffer_3650_s_current_state_reg ( .D(
        KeyArray_S10reg_gff_1_SFF_6_n5), .CK(clk), .Q(new_AGEMA_signal_5538)
         );
  DFF_X1 new_AGEMA_reg_buffer_3654_s_current_state_reg ( .D(
        new_AGEMA_signal_3305), .CK(clk), .Q(new_AGEMA_signal_5542) );
  DFF_X1 new_AGEMA_reg_buffer_3658_s_current_state_reg ( .D(
        KeyArray_S10reg_gff_1_SFF_7_n5), .CK(clk), .Q(new_AGEMA_signal_5546)
         );
  DFF_X1 new_AGEMA_reg_buffer_3662_s_current_state_reg ( .D(
        new_AGEMA_signal_3306), .CK(clk), .Q(new_AGEMA_signal_5550) );
  DFF_X1 new_AGEMA_reg_buffer_3666_s_current_state_reg ( .D(
        KeyArray_S11reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_5554)
         );
  DFF_X1 new_AGEMA_reg_buffer_3670_s_current_state_reg ( .D(
        new_AGEMA_signal_3307), .CK(clk), .Q(new_AGEMA_signal_5558) );
  DFF_X1 new_AGEMA_reg_buffer_3674_s_current_state_reg ( .D(
        KeyArray_S11reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_5562)
         );
  DFF_X1 new_AGEMA_reg_buffer_3678_s_current_state_reg ( .D(
        new_AGEMA_signal_3308), .CK(clk), .Q(new_AGEMA_signal_5566) );
  DFF_X1 new_AGEMA_reg_buffer_3682_s_current_state_reg ( .D(
        KeyArray_S11reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_5570)
         );
  DFF_X1 new_AGEMA_reg_buffer_3686_s_current_state_reg ( .D(
        new_AGEMA_signal_3309), .CK(clk), .Q(new_AGEMA_signal_5574) );
  DFF_X1 new_AGEMA_reg_buffer_3690_s_current_state_reg ( .D(
        KeyArray_S11reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_5578)
         );
  DFF_X1 new_AGEMA_reg_buffer_3694_s_current_state_reg ( .D(
        new_AGEMA_signal_3310), .CK(clk), .Q(new_AGEMA_signal_5582) );
  DFF_X1 new_AGEMA_reg_buffer_3698_s_current_state_reg ( .D(
        KeyArray_S11reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_5586)
         );
  DFF_X1 new_AGEMA_reg_buffer_3702_s_current_state_reg ( .D(
        new_AGEMA_signal_3311), .CK(clk), .Q(new_AGEMA_signal_5590) );
  DFF_X1 new_AGEMA_reg_buffer_3706_s_current_state_reg ( .D(
        KeyArray_S11reg_gff_1_SFF_5_n6), .CK(clk), .Q(new_AGEMA_signal_5594)
         );
  DFF_X1 new_AGEMA_reg_buffer_3710_s_current_state_reg ( .D(
        new_AGEMA_signal_3312), .CK(clk), .Q(new_AGEMA_signal_5598) );
  DFF_X1 new_AGEMA_reg_buffer_3714_s_current_state_reg ( .D(
        KeyArray_S11reg_gff_1_SFF_6_n6), .CK(clk), .Q(new_AGEMA_signal_5602)
         );
  DFF_X1 new_AGEMA_reg_buffer_3718_s_current_state_reg ( .D(
        new_AGEMA_signal_3313), .CK(clk), .Q(new_AGEMA_signal_5606) );
  DFF_X1 new_AGEMA_reg_buffer_3722_s_current_state_reg ( .D(
        KeyArray_S11reg_gff_1_SFF_7_n6), .CK(clk), .Q(new_AGEMA_signal_5610)
         );
  DFF_X1 new_AGEMA_reg_buffer_3726_s_current_state_reg ( .D(
        new_AGEMA_signal_3314), .CK(clk), .Q(new_AGEMA_signal_5614) );
  DFF_X1 new_AGEMA_reg_buffer_3730_s_current_state_reg ( .D(
        KeyArray_S12reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_5618)
         );
  DFF_X1 new_AGEMA_reg_buffer_3734_s_current_state_reg ( .D(
        new_AGEMA_signal_3093), .CK(clk), .Q(new_AGEMA_signal_5622) );
  DFF_X1 new_AGEMA_reg_buffer_3738_s_current_state_reg ( .D(
        KeyArray_S12reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_5626)
         );
  DFF_X1 new_AGEMA_reg_buffer_3742_s_current_state_reg ( .D(
        new_AGEMA_signal_3094), .CK(clk), .Q(new_AGEMA_signal_5630) );
  DFF_X1 new_AGEMA_reg_buffer_3746_s_current_state_reg ( .D(
        KeyArray_S12reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_5634)
         );
  DFF_X1 new_AGEMA_reg_buffer_3750_s_current_state_reg ( .D(
        new_AGEMA_signal_3095), .CK(clk), .Q(new_AGEMA_signal_5638) );
  DFF_X1 new_AGEMA_reg_buffer_3754_s_current_state_reg ( .D(
        KeyArray_S12reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_5642)
         );
  DFF_X1 new_AGEMA_reg_buffer_3758_s_current_state_reg ( .D(
        new_AGEMA_signal_3096), .CK(clk), .Q(new_AGEMA_signal_5646) );
  DFF_X1 new_AGEMA_reg_buffer_3762_s_current_state_reg ( .D(
        KeyArray_S12reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_5650)
         );
  DFF_X1 new_AGEMA_reg_buffer_3766_s_current_state_reg ( .D(
        new_AGEMA_signal_3097), .CK(clk), .Q(new_AGEMA_signal_5654) );
  DFF_X1 new_AGEMA_reg_buffer_3770_s_current_state_reg ( .D(
        KeyArray_S12reg_gff_1_SFF_5_n6), .CK(clk), .Q(new_AGEMA_signal_5658)
         );
  DFF_X1 new_AGEMA_reg_buffer_3774_s_current_state_reg ( .D(
        new_AGEMA_signal_3098), .CK(clk), .Q(new_AGEMA_signal_5662) );
  DFF_X1 new_AGEMA_reg_buffer_3778_s_current_state_reg ( .D(
        KeyArray_S12reg_gff_1_SFF_6_n6), .CK(clk), .Q(new_AGEMA_signal_5666)
         );
  DFF_X1 new_AGEMA_reg_buffer_3782_s_current_state_reg ( .D(
        new_AGEMA_signal_3099), .CK(clk), .Q(new_AGEMA_signal_5670) );
  DFF_X1 new_AGEMA_reg_buffer_3786_s_current_state_reg ( .D(
        KeyArray_S12reg_gff_1_SFF_7_n6), .CK(clk), .Q(new_AGEMA_signal_5674)
         );
  DFF_X1 new_AGEMA_reg_buffer_3790_s_current_state_reg ( .D(
        new_AGEMA_signal_3100), .CK(clk), .Q(new_AGEMA_signal_5678) );
  DFF_X1 new_AGEMA_reg_buffer_3794_s_current_state_reg ( .D(
        KeyArray_S13reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_5682)
         );
  DFF_X1 new_AGEMA_reg_buffer_3798_s_current_state_reg ( .D(
        new_AGEMA_signal_3101), .CK(clk), .Q(new_AGEMA_signal_5686) );
  DFF_X1 new_AGEMA_reg_buffer_3802_s_current_state_reg ( .D(
        KeyArray_S13reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_5690)
         );
  DFF_X1 new_AGEMA_reg_buffer_3806_s_current_state_reg ( .D(
        new_AGEMA_signal_3102), .CK(clk), .Q(new_AGEMA_signal_5694) );
  DFF_X1 new_AGEMA_reg_buffer_3810_s_current_state_reg ( .D(
        KeyArray_S13reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_5698)
         );
  DFF_X1 new_AGEMA_reg_buffer_3814_s_current_state_reg ( .D(
        new_AGEMA_signal_3103), .CK(clk), .Q(new_AGEMA_signal_5702) );
  DFF_X1 new_AGEMA_reg_buffer_3818_s_current_state_reg ( .D(
        KeyArray_S13reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_5706)
         );
  DFF_X1 new_AGEMA_reg_buffer_3822_s_current_state_reg ( .D(
        new_AGEMA_signal_3104), .CK(clk), .Q(new_AGEMA_signal_5710) );
  DFF_X1 new_AGEMA_reg_buffer_3826_s_current_state_reg ( .D(
        KeyArray_S13reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_5714)
         );
  DFF_X1 new_AGEMA_reg_buffer_3830_s_current_state_reg ( .D(
        new_AGEMA_signal_3105), .CK(clk), .Q(new_AGEMA_signal_5718) );
  DFF_X1 new_AGEMA_reg_buffer_3834_s_current_state_reg ( .D(
        KeyArray_S13reg_gff_1_SFF_5_n5), .CK(clk), .Q(new_AGEMA_signal_5722)
         );
  DFF_X1 new_AGEMA_reg_buffer_3838_s_current_state_reg ( .D(
        new_AGEMA_signal_3106), .CK(clk), .Q(new_AGEMA_signal_5726) );
  DFF_X1 new_AGEMA_reg_buffer_3842_s_current_state_reg ( .D(
        KeyArray_S13reg_gff_1_SFF_6_n5), .CK(clk), .Q(new_AGEMA_signal_5730)
         );
  DFF_X1 new_AGEMA_reg_buffer_3846_s_current_state_reg ( .D(
        new_AGEMA_signal_3107), .CK(clk), .Q(new_AGEMA_signal_5734) );
  DFF_X1 new_AGEMA_reg_buffer_3850_s_current_state_reg ( .D(
        KeyArray_S13reg_gff_1_SFF_7_n5), .CK(clk), .Q(new_AGEMA_signal_5738)
         );
  DFF_X1 new_AGEMA_reg_buffer_3854_s_current_state_reg ( .D(
        new_AGEMA_signal_3108), .CK(clk), .Q(new_AGEMA_signal_5742) );
  DFF_X1 new_AGEMA_reg_buffer_3858_s_current_state_reg ( .D(
        KeyArray_S20reg_gff_1_SFF_0_n5), .CK(clk), .Q(new_AGEMA_signal_5746)
         );
  DFF_X1 new_AGEMA_reg_buffer_3862_s_current_state_reg ( .D(
        new_AGEMA_signal_3315), .CK(clk), .Q(new_AGEMA_signal_5750) );
  DFF_X1 new_AGEMA_reg_buffer_3866_s_current_state_reg ( .D(
        KeyArray_S20reg_gff_1_SFF_1_n5), .CK(clk), .Q(new_AGEMA_signal_5754)
         );
  DFF_X1 new_AGEMA_reg_buffer_3870_s_current_state_reg ( .D(
        new_AGEMA_signal_3316), .CK(clk), .Q(new_AGEMA_signal_5758) );
  DFF_X1 new_AGEMA_reg_buffer_3874_s_current_state_reg ( .D(
        KeyArray_S20reg_gff_1_SFF_2_n5), .CK(clk), .Q(new_AGEMA_signal_5762)
         );
  DFF_X1 new_AGEMA_reg_buffer_3878_s_current_state_reg ( .D(
        new_AGEMA_signal_3317), .CK(clk), .Q(new_AGEMA_signal_5766) );
  DFF_X1 new_AGEMA_reg_buffer_3882_s_current_state_reg ( .D(
        KeyArray_S20reg_gff_1_SFF_3_n5), .CK(clk), .Q(new_AGEMA_signal_5770)
         );
  DFF_X1 new_AGEMA_reg_buffer_3886_s_current_state_reg ( .D(
        new_AGEMA_signal_3318), .CK(clk), .Q(new_AGEMA_signal_5774) );
  DFF_X1 new_AGEMA_reg_buffer_3890_s_current_state_reg ( .D(
        KeyArray_S20reg_gff_1_SFF_4_n5), .CK(clk), .Q(new_AGEMA_signal_5778)
         );
  DFF_X1 new_AGEMA_reg_buffer_3894_s_current_state_reg ( .D(
        new_AGEMA_signal_3319), .CK(clk), .Q(new_AGEMA_signal_5782) );
  DFF_X1 new_AGEMA_reg_buffer_3898_s_current_state_reg ( .D(
        KeyArray_S20reg_gff_1_SFF_5_n5), .CK(clk), .Q(new_AGEMA_signal_5786)
         );
  DFF_X1 new_AGEMA_reg_buffer_3902_s_current_state_reg ( .D(
        new_AGEMA_signal_3320), .CK(clk), .Q(new_AGEMA_signal_5790) );
  DFF_X1 new_AGEMA_reg_buffer_3906_s_current_state_reg ( .D(
        KeyArray_S20reg_gff_1_SFF_6_n5), .CK(clk), .Q(new_AGEMA_signal_5794)
         );
  DFF_X1 new_AGEMA_reg_buffer_3910_s_current_state_reg ( .D(
        new_AGEMA_signal_3321), .CK(clk), .Q(new_AGEMA_signal_5798) );
  DFF_X1 new_AGEMA_reg_buffer_3914_s_current_state_reg ( .D(
        KeyArray_S20reg_gff_1_SFF_7_n5), .CK(clk), .Q(new_AGEMA_signal_5802)
         );
  DFF_X1 new_AGEMA_reg_buffer_3918_s_current_state_reg ( .D(
        new_AGEMA_signal_3322), .CK(clk), .Q(new_AGEMA_signal_5806) );
  DFF_X1 new_AGEMA_reg_buffer_3922_s_current_state_reg ( .D(
        KeyArray_S21reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_5810)
         );
  DFF_X1 new_AGEMA_reg_buffer_3926_s_current_state_reg ( .D(
        new_AGEMA_signal_3323), .CK(clk), .Q(new_AGEMA_signal_5814) );
  DFF_X1 new_AGEMA_reg_buffer_3930_s_current_state_reg ( .D(
        KeyArray_S21reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_5818)
         );
  DFF_X1 new_AGEMA_reg_buffer_3934_s_current_state_reg ( .D(
        new_AGEMA_signal_3324), .CK(clk), .Q(new_AGEMA_signal_5822) );
  DFF_X1 new_AGEMA_reg_buffer_3938_s_current_state_reg ( .D(
        KeyArray_S21reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_5826)
         );
  DFF_X1 new_AGEMA_reg_buffer_3942_s_current_state_reg ( .D(
        new_AGEMA_signal_3325), .CK(clk), .Q(new_AGEMA_signal_5830) );
  DFF_X1 new_AGEMA_reg_buffer_3946_s_current_state_reg ( .D(
        KeyArray_S21reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_5834)
         );
  DFF_X1 new_AGEMA_reg_buffer_3950_s_current_state_reg ( .D(
        new_AGEMA_signal_3326), .CK(clk), .Q(new_AGEMA_signal_5838) );
  DFF_X1 new_AGEMA_reg_buffer_3954_s_current_state_reg ( .D(
        KeyArray_S21reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_5842)
         );
  DFF_X1 new_AGEMA_reg_buffer_3958_s_current_state_reg ( .D(
        new_AGEMA_signal_3327), .CK(clk), .Q(new_AGEMA_signal_5846) );
  DFF_X1 new_AGEMA_reg_buffer_3962_s_current_state_reg ( .D(
        KeyArray_S21reg_gff_1_SFF_5_n6), .CK(clk), .Q(new_AGEMA_signal_5850)
         );
  DFF_X1 new_AGEMA_reg_buffer_3966_s_current_state_reg ( .D(
        new_AGEMA_signal_3328), .CK(clk), .Q(new_AGEMA_signal_5854) );
  DFF_X1 new_AGEMA_reg_buffer_3970_s_current_state_reg ( .D(
        KeyArray_S21reg_gff_1_SFF_6_n6), .CK(clk), .Q(new_AGEMA_signal_5858)
         );
  DFF_X1 new_AGEMA_reg_buffer_3974_s_current_state_reg ( .D(
        new_AGEMA_signal_3329), .CK(clk), .Q(new_AGEMA_signal_5862) );
  DFF_X1 new_AGEMA_reg_buffer_3978_s_current_state_reg ( .D(
        KeyArray_S21reg_gff_1_SFF_7_n6), .CK(clk), .Q(new_AGEMA_signal_5866)
         );
  DFF_X1 new_AGEMA_reg_buffer_3982_s_current_state_reg ( .D(
        new_AGEMA_signal_3330), .CK(clk), .Q(new_AGEMA_signal_5870) );
  DFF_X1 new_AGEMA_reg_buffer_3986_s_current_state_reg ( .D(
        KeyArray_S22reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_5874)
         );
  DFF_X1 new_AGEMA_reg_buffer_3990_s_current_state_reg ( .D(
        new_AGEMA_signal_3331), .CK(clk), .Q(new_AGEMA_signal_5878) );
  DFF_X1 new_AGEMA_reg_buffer_3994_s_current_state_reg ( .D(
        KeyArray_S22reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_5882)
         );
  DFF_X1 new_AGEMA_reg_buffer_3998_s_current_state_reg ( .D(
        new_AGEMA_signal_3332), .CK(clk), .Q(new_AGEMA_signal_5886) );
  DFF_X1 new_AGEMA_reg_buffer_4002_s_current_state_reg ( .D(
        KeyArray_S22reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_5890)
         );
  DFF_X1 new_AGEMA_reg_buffer_4006_s_current_state_reg ( .D(
        new_AGEMA_signal_3333), .CK(clk), .Q(new_AGEMA_signal_5894) );
  DFF_X1 new_AGEMA_reg_buffer_4010_s_current_state_reg ( .D(
        KeyArray_S22reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_5898)
         );
  DFF_X1 new_AGEMA_reg_buffer_4014_s_current_state_reg ( .D(
        new_AGEMA_signal_3334), .CK(clk), .Q(new_AGEMA_signal_5902) );
  DFF_X1 new_AGEMA_reg_buffer_4018_s_current_state_reg ( .D(
        KeyArray_S22reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_5906)
         );
  DFF_X1 new_AGEMA_reg_buffer_4022_s_current_state_reg ( .D(
        new_AGEMA_signal_3335), .CK(clk), .Q(new_AGEMA_signal_5910) );
  DFF_X1 new_AGEMA_reg_buffer_4026_s_current_state_reg ( .D(
        KeyArray_S22reg_gff_1_SFF_5_n6), .CK(clk), .Q(new_AGEMA_signal_5914)
         );
  DFF_X1 new_AGEMA_reg_buffer_4030_s_current_state_reg ( .D(
        new_AGEMA_signal_3336), .CK(clk), .Q(new_AGEMA_signal_5918) );
  DFF_X1 new_AGEMA_reg_buffer_4034_s_current_state_reg ( .D(
        KeyArray_S22reg_gff_1_SFF_6_n6), .CK(clk), .Q(new_AGEMA_signal_5922)
         );
  DFF_X1 new_AGEMA_reg_buffer_4038_s_current_state_reg ( .D(
        new_AGEMA_signal_3337), .CK(clk), .Q(new_AGEMA_signal_5926) );
  DFF_X1 new_AGEMA_reg_buffer_4042_s_current_state_reg ( .D(
        KeyArray_S22reg_gff_1_SFF_7_n6), .CK(clk), .Q(new_AGEMA_signal_5930)
         );
  DFF_X1 new_AGEMA_reg_buffer_4046_s_current_state_reg ( .D(
        new_AGEMA_signal_3338), .CK(clk), .Q(new_AGEMA_signal_5934) );
  DFF_X1 new_AGEMA_reg_buffer_4050_s_current_state_reg ( .D(
        KeyArray_S23reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_5938)
         );
  DFF_X1 new_AGEMA_reg_buffer_4054_s_current_state_reg ( .D(
        new_AGEMA_signal_3339), .CK(clk), .Q(new_AGEMA_signal_5942) );
  DFF_X1 new_AGEMA_reg_buffer_4058_s_current_state_reg ( .D(
        KeyArray_S23reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_5946)
         );
  DFF_X1 new_AGEMA_reg_buffer_4062_s_current_state_reg ( .D(
        new_AGEMA_signal_3340), .CK(clk), .Q(new_AGEMA_signal_5950) );
  DFF_X1 new_AGEMA_reg_buffer_4066_s_current_state_reg ( .D(
        KeyArray_S23reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_5954)
         );
  DFF_X1 new_AGEMA_reg_buffer_4070_s_current_state_reg ( .D(
        new_AGEMA_signal_3341), .CK(clk), .Q(new_AGEMA_signal_5958) );
  DFF_X1 new_AGEMA_reg_buffer_4074_s_current_state_reg ( .D(
        KeyArray_S23reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_5962)
         );
  DFF_X1 new_AGEMA_reg_buffer_4078_s_current_state_reg ( .D(
        new_AGEMA_signal_3342), .CK(clk), .Q(new_AGEMA_signal_5966) );
  DFF_X1 new_AGEMA_reg_buffer_4082_s_current_state_reg ( .D(
        KeyArray_S23reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_5970)
         );
  DFF_X1 new_AGEMA_reg_buffer_4086_s_current_state_reg ( .D(
        new_AGEMA_signal_3343), .CK(clk), .Q(new_AGEMA_signal_5974) );
  DFF_X1 new_AGEMA_reg_buffer_4090_s_current_state_reg ( .D(
        KeyArray_S23reg_gff_1_SFF_5_n5), .CK(clk), .Q(new_AGEMA_signal_5978)
         );
  DFF_X1 new_AGEMA_reg_buffer_4094_s_current_state_reg ( .D(
        new_AGEMA_signal_3344), .CK(clk), .Q(new_AGEMA_signal_5982) );
  DFF_X1 new_AGEMA_reg_buffer_4098_s_current_state_reg ( .D(
        KeyArray_S23reg_gff_1_SFF_6_n5), .CK(clk), .Q(new_AGEMA_signal_5986)
         );
  DFF_X1 new_AGEMA_reg_buffer_4102_s_current_state_reg ( .D(
        new_AGEMA_signal_3345), .CK(clk), .Q(new_AGEMA_signal_5990) );
  DFF_X1 new_AGEMA_reg_buffer_4106_s_current_state_reg ( .D(
        KeyArray_S23reg_gff_1_SFF_7_n5), .CK(clk), .Q(new_AGEMA_signal_5994)
         );
  DFF_X1 new_AGEMA_reg_buffer_4110_s_current_state_reg ( .D(
        new_AGEMA_signal_3346), .CK(clk), .Q(new_AGEMA_signal_5998) );
  DFF_X1 new_AGEMA_reg_buffer_4114_s_current_state_reg ( .D(
        KeyArray_S31reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_6002)
         );
  DFF_X1 new_AGEMA_reg_buffer_4118_s_current_state_reg ( .D(
        new_AGEMA_signal_3347), .CK(clk), .Q(new_AGEMA_signal_6006) );
  DFF_X1 new_AGEMA_reg_buffer_4122_s_current_state_reg ( .D(
        KeyArray_S31reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_6010)
         );
  DFF_X1 new_AGEMA_reg_buffer_4126_s_current_state_reg ( .D(
        new_AGEMA_signal_3348), .CK(clk), .Q(new_AGEMA_signal_6014) );
  DFF_X1 new_AGEMA_reg_buffer_4130_s_current_state_reg ( .D(
        KeyArray_S31reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_6018)
         );
  DFF_X1 new_AGEMA_reg_buffer_4134_s_current_state_reg ( .D(
        new_AGEMA_signal_3349), .CK(clk), .Q(new_AGEMA_signal_6022) );
  DFF_X1 new_AGEMA_reg_buffer_4138_s_current_state_reg ( .D(
        KeyArray_S31reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_6026)
         );
  DFF_X1 new_AGEMA_reg_buffer_4142_s_current_state_reg ( .D(
        new_AGEMA_signal_3350), .CK(clk), .Q(new_AGEMA_signal_6030) );
  DFF_X1 new_AGEMA_reg_buffer_4146_s_current_state_reg ( .D(
        KeyArray_S31reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_6034)
         );
  DFF_X1 new_AGEMA_reg_buffer_4150_s_current_state_reg ( .D(
        new_AGEMA_signal_3351), .CK(clk), .Q(new_AGEMA_signal_6038) );
  DFF_X1 new_AGEMA_reg_buffer_4154_s_current_state_reg ( .D(
        KeyArray_S31reg_gff_1_SFF_5_n6), .CK(clk), .Q(new_AGEMA_signal_6042)
         );
  DFF_X1 new_AGEMA_reg_buffer_4158_s_current_state_reg ( .D(
        new_AGEMA_signal_3352), .CK(clk), .Q(new_AGEMA_signal_6046) );
  DFF_X1 new_AGEMA_reg_buffer_4162_s_current_state_reg ( .D(
        KeyArray_S31reg_gff_1_SFF_6_n6), .CK(clk), .Q(new_AGEMA_signal_6050)
         );
  DFF_X1 new_AGEMA_reg_buffer_4166_s_current_state_reg ( .D(
        new_AGEMA_signal_3353), .CK(clk), .Q(new_AGEMA_signal_6054) );
  DFF_X1 new_AGEMA_reg_buffer_4170_s_current_state_reg ( .D(
        KeyArray_S31reg_gff_1_SFF_7_n6), .CK(clk), .Q(new_AGEMA_signal_6058)
         );
  DFF_X1 new_AGEMA_reg_buffer_4174_s_current_state_reg ( .D(
        new_AGEMA_signal_3354), .CK(clk), .Q(new_AGEMA_signal_6062) );
  DFF_X1 new_AGEMA_reg_buffer_4178_s_current_state_reg ( .D(
        KeyArray_S32reg_gff_1_SFF_0_n6), .CK(clk), .Q(new_AGEMA_signal_6066)
         );
  DFF_X1 new_AGEMA_reg_buffer_4182_s_current_state_reg ( .D(
        new_AGEMA_signal_3355), .CK(clk), .Q(new_AGEMA_signal_6070) );
  DFF_X1 new_AGEMA_reg_buffer_4186_s_current_state_reg ( .D(
        KeyArray_S32reg_gff_1_SFF_1_n6), .CK(clk), .Q(new_AGEMA_signal_6074)
         );
  DFF_X1 new_AGEMA_reg_buffer_4190_s_current_state_reg ( .D(
        new_AGEMA_signal_3356), .CK(clk), .Q(new_AGEMA_signal_6078) );
  DFF_X1 new_AGEMA_reg_buffer_4194_s_current_state_reg ( .D(
        KeyArray_S32reg_gff_1_SFF_2_n6), .CK(clk), .Q(new_AGEMA_signal_6082)
         );
  DFF_X1 new_AGEMA_reg_buffer_4198_s_current_state_reg ( .D(
        new_AGEMA_signal_3357), .CK(clk), .Q(new_AGEMA_signal_6086) );
  DFF_X1 new_AGEMA_reg_buffer_4202_s_current_state_reg ( .D(
        KeyArray_S32reg_gff_1_SFF_3_n6), .CK(clk), .Q(new_AGEMA_signal_6090)
         );
  DFF_X1 new_AGEMA_reg_buffer_4206_s_current_state_reg ( .D(
        new_AGEMA_signal_3358), .CK(clk), .Q(new_AGEMA_signal_6094) );
  DFF_X1 new_AGEMA_reg_buffer_4210_s_current_state_reg ( .D(
        KeyArray_S32reg_gff_1_SFF_4_n6), .CK(clk), .Q(new_AGEMA_signal_6098)
         );
  DFF_X1 new_AGEMA_reg_buffer_4214_s_current_state_reg ( .D(
        new_AGEMA_signal_3359), .CK(clk), .Q(new_AGEMA_signal_6102) );
  DFF_X1 new_AGEMA_reg_buffer_4218_s_current_state_reg ( .D(
        KeyArray_S32reg_gff_1_SFF_5_n6), .CK(clk), .Q(new_AGEMA_signal_6106)
         );
  DFF_X1 new_AGEMA_reg_buffer_4222_s_current_state_reg ( .D(
        new_AGEMA_signal_3360), .CK(clk), .Q(new_AGEMA_signal_6110) );
  DFF_X1 new_AGEMA_reg_buffer_4226_s_current_state_reg ( .D(
        KeyArray_S32reg_gff_1_SFF_6_n5), .CK(clk), .Q(new_AGEMA_signal_6114)
         );
  DFF_X1 new_AGEMA_reg_buffer_4230_s_current_state_reg ( .D(
        new_AGEMA_signal_3361), .CK(clk), .Q(new_AGEMA_signal_6118) );
  DFF_X1 new_AGEMA_reg_buffer_4234_s_current_state_reg ( .D(
        KeyArray_S32reg_gff_1_SFF_7_n5), .CK(clk), .Q(new_AGEMA_signal_6122)
         );
  DFF_X1 new_AGEMA_reg_buffer_4238_s_current_state_reg ( .D(
        new_AGEMA_signal_3362), .CK(clk), .Q(new_AGEMA_signal_6126) );
  DFF_X1 new_AGEMA_reg_buffer_4242_s_current_state_reg ( .D(
        KeyArray_S33reg_gff_1_SFF_0_n5), .CK(clk), .Q(new_AGEMA_signal_6130)
         );
  DFF_X1 new_AGEMA_reg_buffer_4246_s_current_state_reg ( .D(
        new_AGEMA_signal_3363), .CK(clk), .Q(new_AGEMA_signal_6134) );
  DFF_X1 new_AGEMA_reg_buffer_4250_s_current_state_reg ( .D(
        KeyArray_S33reg_gff_1_SFF_1_n5), .CK(clk), .Q(new_AGEMA_signal_6138)
         );
  DFF_X1 new_AGEMA_reg_buffer_4254_s_current_state_reg ( .D(
        new_AGEMA_signal_3364), .CK(clk), .Q(new_AGEMA_signal_6142) );
  DFF_X1 new_AGEMA_reg_buffer_4258_s_current_state_reg ( .D(
        KeyArray_S33reg_gff_1_SFF_2_n5), .CK(clk), .Q(new_AGEMA_signal_6146)
         );
  DFF_X1 new_AGEMA_reg_buffer_4262_s_current_state_reg ( .D(
        new_AGEMA_signal_3365), .CK(clk), .Q(new_AGEMA_signal_6150) );
  DFF_X1 new_AGEMA_reg_buffer_4266_s_current_state_reg ( .D(
        KeyArray_S33reg_gff_1_SFF_3_n5), .CK(clk), .Q(new_AGEMA_signal_6154)
         );
  DFF_X1 new_AGEMA_reg_buffer_4270_s_current_state_reg ( .D(
        new_AGEMA_signal_3366), .CK(clk), .Q(new_AGEMA_signal_6158) );
  DFF_X1 new_AGEMA_reg_buffer_4274_s_current_state_reg ( .D(
        KeyArray_S33reg_gff_1_SFF_4_n5), .CK(clk), .Q(new_AGEMA_signal_6162)
         );
  DFF_X1 new_AGEMA_reg_buffer_4278_s_current_state_reg ( .D(
        new_AGEMA_signal_3367), .CK(clk), .Q(new_AGEMA_signal_6166) );
  DFF_X1 new_AGEMA_reg_buffer_4282_s_current_state_reg ( .D(
        KeyArray_S33reg_gff_1_SFF_5_n5), .CK(clk), .Q(new_AGEMA_signal_6170)
         );
  DFF_X1 new_AGEMA_reg_buffer_4286_s_current_state_reg ( .D(
        new_AGEMA_signal_3368), .CK(clk), .Q(new_AGEMA_signal_6174) );
  DFF_X1 new_AGEMA_reg_buffer_4290_s_current_state_reg ( .D(
        KeyArray_S33reg_gff_1_SFF_6_n5), .CK(clk), .Q(new_AGEMA_signal_6178)
         );
  DFF_X1 new_AGEMA_reg_buffer_4294_s_current_state_reg ( .D(
        new_AGEMA_signal_3369), .CK(clk), .Q(new_AGEMA_signal_6182) );
  DFF_X1 new_AGEMA_reg_buffer_4298_s_current_state_reg ( .D(
        KeyArray_S33reg_gff_1_SFF_7_n5), .CK(clk), .Q(new_AGEMA_signal_6186)
         );
  DFF_X1 new_AGEMA_reg_buffer_4302_s_current_state_reg ( .D(
        new_AGEMA_signal_3370), .CK(clk), .Q(new_AGEMA_signal_6190) );
  DFF_X1 new_AGEMA_reg_buffer_4306_s_current_state_reg ( .D(calcRCon_n51),
        .CK(clk), .Q(new_AGEMA_signal_6194) );
  DFF_X1 new_AGEMA_reg_buffer_4310_s_current_state_reg ( .D(calcRCon_n50),
        .CK(clk), .Q(new_AGEMA_signal_6198) );
  DFF_X1 new_AGEMA_reg_buffer_4314_s_current_state_reg ( .D(calcRCon_n49),
        .CK(clk), .Q(new_AGEMA_signal_6202) );
  DFF_X1 new_AGEMA_reg_buffer_4318_s_current_state_reg ( .D(calcRCon_n48),
        .CK(clk), .Q(new_AGEMA_signal_6206) );
  DFF_X1 new_AGEMA_reg_buffer_4322_s_current_state_reg ( .D(calcRCon_n47),
        .CK(clk), .Q(new_AGEMA_signal_6210) );
  DFF_X1 new_AGEMA_reg_buffer_4326_s_current_state_reg ( .D(calcRCon_n46),
        .CK(clk), .Q(new_AGEMA_signal_6214) );
  DFF_X1 new_AGEMA_reg_buffer_4330_s_current_state_reg ( .D(calcRCon_n45),
        .CK(clk), .Q(new_AGEMA_signal_6218) );
  DFF_X1 new_AGEMA_reg_buffer_4334_s_current_state_reg ( .D(calcRCon_n44),
        .CK(clk), .Q(new_AGEMA_signal_6222) );
  DFF_X1 new_AGEMA_reg_buffer_4338_s_current_state_reg ( .D(n189), .CK(clk),
        .Q(new_AGEMA_signal_6226) );
  XOR2_X1 Inst_bSbox_AND_M25_U1_U16 ( .A(Fresh[18]), .B(
        Inst_bSbox_AND_M25_U1_n23), .Z(Inst_bSbox_AND_M25_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M25_U1_U15 ( .A1(new_AGEMA_signal_3374), .A2(
        Inst_bSbox_AND_M25_U1_n22), .ZN(Inst_bSbox_AND_M25_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M25_U1_U14 ( .A(Fresh[18]), .B(
        Inst_bSbox_AND_M25_U1_n21), .Z(Inst_bSbox_AND_M25_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M25_U1_U13 ( .A1(Inst_bSbox_M22), .A2(
        Inst_bSbox_AND_M25_U1_n22), .ZN(Inst_bSbox_AND_M25_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M25_U1_U12 ( .A(Inst_bSbox_AND_M25_U1_n20), .B(
        Inst_bSbox_AND_M25_U1_n19), .ZN(Inst_bSbox_M25) );
  NAND2_X1 Inst_bSbox_AND_M25_U1_U11 ( .A1(Inst_bSbox_AND_M25_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M25_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M25_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M25_U1_U10 ( .A(Inst_bSbox_AND_M25_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M25_U1_z[0]), .Z(Inst_bSbox_AND_M25_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M25_U1_U9 ( .A(Inst_bSbox_AND_M25_U1_n18), .B(
        Inst_bSbox_AND_M25_U1_n17), .ZN(new_AGEMA_signal_3384) );
  NAND2_X1 Inst_bSbox_AND_M25_U1_U8 ( .A1(Inst_bSbox_AND_M25_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M25_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M25_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M25_U1_U7 ( .A(Inst_bSbox_AND_M25_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M25_U1_z[1]), .Z(Inst_bSbox_AND_M25_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M25_U1_U6 ( .A(new_AGEMA_signal_3372), .B(
        Inst_bSbox_AND_M25_U1_n22), .ZN(Inst_bSbox_AND_M25_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M25_U1_U5 ( .A(Inst_bSbox_M20), .B(
        Inst_bSbox_AND_M25_U1_n22), .ZN(Inst_bSbox_AND_M25_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M25_U1_U4 ( .A(Fresh[19]), .ZN(
        Inst_bSbox_AND_M25_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M25_U1_U3 ( .A1(new_AGEMA_signal_3374), .A2(
        new_AGEMA_signal_3372), .ZN(Inst_bSbox_AND_M25_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M25_U1_U2 ( .A1(Inst_bSbox_M22), .A2(Inst_bSbox_M20),
        .ZN(Inst_bSbox_AND_M25_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M25_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M25_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M25_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M22),
        .CK(clk), .Q(Inst_bSbox_AND_M25_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M25_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M25_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M25_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M25_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M25_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M25_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M25_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3374), .CK(clk), .Q(Inst_bSbox_AND_M25_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M25_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M25_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M25_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M25_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_M26_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3610), .B(
        Inst_bSbox_M25), .Z(Inst_bSbox_M26) );
  XOR2_X1 Inst_bSbox_XOR_M26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3611), .B(
        new_AGEMA_signal_3384), .Z(new_AGEMA_signal_3388) );
  XOR2_X1 Inst_bSbox_XOR_M28_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3612), .B(
        Inst_bSbox_M25), .Z(Inst_bSbox_M28) );
  XOR2_X1 Inst_bSbox_XOR_M28_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3613), .B(
        new_AGEMA_signal_3384), .Z(new_AGEMA_signal_3389) );
  XOR2_X1 Inst_bSbox_AND_M31_U1_U16 ( .A(Fresh[20]), .B(
        Inst_bSbox_AND_M31_U1_n23), .Z(Inst_bSbox_AND_M31_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M31_U1_U15 ( .A1(new_AGEMA_signal_3372), .A2(
        Inst_bSbox_AND_M31_U1_n22), .ZN(Inst_bSbox_AND_M31_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M31_U1_U14 ( .A(Fresh[20]), .B(
        Inst_bSbox_AND_M31_U1_n21), .Z(Inst_bSbox_AND_M31_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M31_U1_U13 ( .A1(Inst_bSbox_M20), .A2(
        Inst_bSbox_AND_M31_U1_n22), .ZN(Inst_bSbox_AND_M31_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M31_U1_U12 ( .A(Inst_bSbox_AND_M31_U1_n20), .B(
        Inst_bSbox_AND_M31_U1_n19), .ZN(Inst_bSbox_M31) );
  NAND2_X1 Inst_bSbox_AND_M31_U1_U11 ( .A1(Inst_bSbox_AND_M31_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M31_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M31_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M31_U1_U10 ( .A(Inst_bSbox_AND_M31_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M31_U1_z[0]), .Z(Inst_bSbox_AND_M31_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M31_U1_U9 ( .A(Inst_bSbox_AND_M31_U1_n18), .B(
        Inst_bSbox_AND_M31_U1_n17), .ZN(new_AGEMA_signal_3390) );
  NAND2_X1 Inst_bSbox_AND_M31_U1_U8 ( .A1(Inst_bSbox_AND_M31_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M31_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M31_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M31_U1_U7 ( .A(Inst_bSbox_AND_M31_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M31_U1_z[1]), .Z(Inst_bSbox_AND_M31_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M31_U1_U6 ( .A(new_AGEMA_signal_3383), .B(
        Inst_bSbox_AND_M31_U1_n22), .ZN(Inst_bSbox_AND_M31_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M31_U1_U5 ( .A(Inst_bSbox_M23), .B(
        Inst_bSbox_AND_M31_U1_n22), .ZN(Inst_bSbox_AND_M31_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M31_U1_U4 ( .A(Fresh[21]), .ZN(
        Inst_bSbox_AND_M31_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M31_U1_U3 ( .A1(Inst_bSbox_M20), .A2(Inst_bSbox_M23),
        .ZN(Inst_bSbox_AND_M31_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M31_U1_U2 ( .A1(new_AGEMA_signal_3372), .A2(
        new_AGEMA_signal_3383), .ZN(Inst_bSbox_AND_M31_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M31_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M31_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M31_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M20),
        .CK(clk), .Q(Inst_bSbox_AND_M31_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M31_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M31_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M31_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M31_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M31_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M31_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M31_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3372), .CK(clk), .Q(Inst_bSbox_AND_M31_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M31_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M31_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M31_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M31_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_M33_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3614), .B(
        Inst_bSbox_M25), .Z(Inst_bSbox_M33) );
  XOR2_X1 Inst_bSbox_XOR_M33_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3615), .B(
        new_AGEMA_signal_3384), .Z(new_AGEMA_signal_3391) );
  XOR2_X1 Inst_bSbox_AND_M34_U1_U16 ( .A(Fresh[22]), .B(
        Inst_bSbox_AND_M34_U1_n23), .Z(Inst_bSbox_AND_M34_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M34_U1_U15 ( .A1(new_AGEMA_signal_3373), .A2(
        Inst_bSbox_AND_M34_U1_n22), .ZN(Inst_bSbox_AND_M34_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M34_U1_U14 ( .A(Fresh[22]), .B(
        Inst_bSbox_AND_M34_U1_n21), .Z(Inst_bSbox_AND_M34_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M34_U1_U13 ( .A1(Inst_bSbox_M21), .A2(
        Inst_bSbox_AND_M34_U1_n22), .ZN(Inst_bSbox_AND_M34_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M34_U1_U12 ( .A(Inst_bSbox_AND_M34_U1_n20), .B(
        Inst_bSbox_AND_M34_U1_n19), .ZN(Inst_bSbox_M34) );
  NAND2_X1 Inst_bSbox_AND_M34_U1_U11 ( .A1(Inst_bSbox_AND_M34_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M34_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M34_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M34_U1_U10 ( .A(Inst_bSbox_AND_M34_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M34_U1_z[0]), .Z(Inst_bSbox_AND_M34_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M34_U1_U9 ( .A(Inst_bSbox_AND_M34_U1_n18), .B(
        Inst_bSbox_AND_M34_U1_n17), .ZN(new_AGEMA_signal_3386) );
  NAND2_X1 Inst_bSbox_AND_M34_U1_U8 ( .A1(Inst_bSbox_AND_M34_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M34_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M34_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M34_U1_U7 ( .A(Inst_bSbox_AND_M34_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M34_U1_z[1]), .Z(Inst_bSbox_AND_M34_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M34_U1_U6 ( .A(new_AGEMA_signal_3374), .B(
        Inst_bSbox_AND_M34_U1_n22), .ZN(Inst_bSbox_AND_M34_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M34_U1_U5 ( .A(Inst_bSbox_M22), .B(
        Inst_bSbox_AND_M34_U1_n22), .ZN(Inst_bSbox_AND_M34_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M34_U1_U4 ( .A(Fresh[23]), .ZN(
        Inst_bSbox_AND_M34_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M34_U1_U3 ( .A1(new_AGEMA_signal_3373), .A2(
        new_AGEMA_signal_3374), .ZN(Inst_bSbox_AND_M34_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M34_U1_U2 ( .A1(Inst_bSbox_M21), .A2(Inst_bSbox_M22),
        .ZN(Inst_bSbox_AND_M34_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M34_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M34_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M34_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M21),
        .CK(clk), .Q(Inst_bSbox_AND_M34_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M34_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M34_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M34_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M34_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M34_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M34_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M34_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3373), .CK(clk), .Q(Inst_bSbox_AND_M34_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M34_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M34_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M34_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M34_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_M36_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3616), .B(
        Inst_bSbox_M25), .Z(Inst_bSbox_M36) );
  XOR2_X1 Inst_bSbox_XOR_M36_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3617), .B(
        new_AGEMA_signal_3384), .Z(new_AGEMA_signal_3396) );
  DFF_X1 new_AGEMA_reg_buffer_1722_s_current_state_reg ( .D(Inst_bSbox_M21),
        .CK(clk), .Q(new_AGEMA_signal_3610) );
  DFF_X1 new_AGEMA_reg_buffer_1723_s_current_state_reg ( .D(
        new_AGEMA_signal_3373), .CK(clk), .Q(new_AGEMA_signal_3611) );
  DFF_X1 new_AGEMA_reg_buffer_1724_s_current_state_reg ( .D(Inst_bSbox_M23),
        .CK(clk), .Q(new_AGEMA_signal_3612) );
  DFF_X1 new_AGEMA_reg_buffer_1725_s_current_state_reg ( .D(
        new_AGEMA_signal_3383), .CK(clk), .Q(new_AGEMA_signal_3613) );
  DFF_X1 new_AGEMA_reg_buffer_1726_s_current_state_reg ( .D(Inst_bSbox_M27),
        .CK(clk), .Q(new_AGEMA_signal_3614) );
  DFF_X1 new_AGEMA_reg_buffer_1727_s_current_state_reg ( .D(
        new_AGEMA_signal_3385), .CK(clk), .Q(new_AGEMA_signal_3615) );
  DFF_X1 new_AGEMA_reg_buffer_1728_s_current_state_reg ( .D(Inst_bSbox_M24),
        .CK(clk), .Q(new_AGEMA_signal_3616) );
  DFF_X1 new_AGEMA_reg_buffer_1729_s_current_state_reg ( .D(
        new_AGEMA_signal_3387), .CK(clk), .Q(new_AGEMA_signal_3617) );
  DFF_X1 new_AGEMA_reg_buffer_1739_s_current_state_reg ( .D(
        new_AGEMA_signal_3626), .CK(clk), .Q(new_AGEMA_signal_3627) );
  DFF_X1 new_AGEMA_reg_buffer_1743_s_current_state_reg ( .D(
        new_AGEMA_signal_3630), .CK(clk), .Q(new_AGEMA_signal_3631) );
  DFF_X1 new_AGEMA_reg_buffer_1747_s_current_state_reg ( .D(
        new_AGEMA_signal_3634), .CK(clk), .Q(new_AGEMA_signal_3635) );
  DFF_X1 new_AGEMA_reg_buffer_1751_s_current_state_reg ( .D(
        new_AGEMA_signal_3638), .CK(clk), .Q(new_AGEMA_signal_3639) );
  DFF_X1 new_AGEMA_reg_buffer_1755_s_current_state_reg ( .D(
        new_AGEMA_signal_3642), .CK(clk), .Q(new_AGEMA_signal_3643) );
  DFF_X1 new_AGEMA_reg_buffer_1759_s_current_state_reg ( .D(
        new_AGEMA_signal_3646), .CK(clk), .Q(new_AGEMA_signal_3647) );
  DFF_X1 new_AGEMA_reg_buffer_1763_s_current_state_reg ( .D(
        new_AGEMA_signal_3650), .CK(clk), .Q(new_AGEMA_signal_3651) );
  DFF_X1 new_AGEMA_reg_buffer_1767_s_current_state_reg ( .D(
        new_AGEMA_signal_3654), .CK(clk), .Q(new_AGEMA_signal_3655) );
  DFF_X1 new_AGEMA_reg_buffer_1771_s_current_state_reg ( .D(
        new_AGEMA_signal_3658), .CK(clk), .Q(new_AGEMA_signal_3659) );
  DFF_X1 new_AGEMA_reg_buffer_1775_s_current_state_reg ( .D(
        new_AGEMA_signal_3662), .CK(clk), .Q(new_AGEMA_signal_3663) );
  DFF_X1 new_AGEMA_reg_buffer_1779_s_current_state_reg ( .D(
        new_AGEMA_signal_3666), .CK(clk), .Q(new_AGEMA_signal_3667) );
  DFF_X1 new_AGEMA_reg_buffer_1783_s_current_state_reg ( .D(
        new_AGEMA_signal_3670), .CK(clk), .Q(new_AGEMA_signal_3671) );
  DFF_X1 new_AGEMA_reg_buffer_1787_s_current_state_reg ( .D(
        new_AGEMA_signal_3674), .CK(clk), .Q(new_AGEMA_signal_3675) );
  DFF_X1 new_AGEMA_reg_buffer_1791_s_current_state_reg ( .D(
        new_AGEMA_signal_3678), .CK(clk), .Q(new_AGEMA_signal_3679) );
  DFF_X1 new_AGEMA_reg_buffer_1795_s_current_state_reg ( .D(
        new_AGEMA_signal_3682), .CK(clk), .Q(new_AGEMA_signal_3683) );
  DFF_X1 new_AGEMA_reg_buffer_1799_s_current_state_reg ( .D(
        new_AGEMA_signal_3686), .CK(clk), .Q(new_AGEMA_signal_3687) );
  DFF_X1 new_AGEMA_reg_buffer_1803_s_current_state_reg ( .D(
        new_AGEMA_signal_3690), .CK(clk), .Q(new_AGEMA_signal_3691) );
  DFF_X1 new_AGEMA_reg_buffer_1807_s_current_state_reg ( .D(
        new_AGEMA_signal_3694), .CK(clk), .Q(new_AGEMA_signal_3695) );
  DFF_X1 new_AGEMA_reg_buffer_1811_s_current_state_reg ( .D(
        new_AGEMA_signal_3698), .CK(clk), .Q(new_AGEMA_signal_3699) );
  DFF_X1 new_AGEMA_reg_buffer_1815_s_current_state_reg ( .D(
        new_AGEMA_signal_3702), .CK(clk), .Q(new_AGEMA_signal_3703) );
  DFF_X1 new_AGEMA_reg_buffer_1819_s_current_state_reg ( .D(
        new_AGEMA_signal_3706), .CK(clk), .Q(new_AGEMA_signal_3707) );
  DFF_X1 new_AGEMA_reg_buffer_1823_s_current_state_reg ( .D(
        new_AGEMA_signal_3710), .CK(clk), .Q(new_AGEMA_signal_3711) );
  DFF_X1 new_AGEMA_reg_buffer_1827_s_current_state_reg ( .D(
        new_AGEMA_signal_3714), .CK(clk), .Q(new_AGEMA_signal_3715) );
  DFF_X1 new_AGEMA_reg_buffer_1831_s_current_state_reg ( .D(
        new_AGEMA_signal_3718), .CK(clk), .Q(new_AGEMA_signal_3719) );
  DFF_X1 new_AGEMA_reg_buffer_1835_s_current_state_reg ( .D(
        new_AGEMA_signal_3722), .CK(clk), .Q(new_AGEMA_signal_3723) );
  DFF_X1 new_AGEMA_reg_buffer_1839_s_current_state_reg ( .D(
        new_AGEMA_signal_3726), .CK(clk), .Q(new_AGEMA_signal_3727) );
  DFF_X1 new_AGEMA_reg_buffer_1843_s_current_state_reg ( .D(
        new_AGEMA_signal_3730), .CK(clk), .Q(new_AGEMA_signal_3731) );
  DFF_X1 new_AGEMA_reg_buffer_1847_s_current_state_reg ( .D(
        new_AGEMA_signal_3734), .CK(clk), .Q(new_AGEMA_signal_3735) );
  DFF_X1 new_AGEMA_reg_buffer_1851_s_current_state_reg ( .D(
        new_AGEMA_signal_3738), .CK(clk), .Q(new_AGEMA_signal_3739) );
  DFF_X1 new_AGEMA_reg_buffer_1855_s_current_state_reg ( .D(
        new_AGEMA_signal_3742), .CK(clk), .Q(new_AGEMA_signal_3743) );
  DFF_X1 new_AGEMA_reg_buffer_1859_s_current_state_reg ( .D(
        new_AGEMA_signal_3746), .CK(clk), .Q(new_AGEMA_signal_3747) );
  DFF_X1 new_AGEMA_reg_buffer_1863_s_current_state_reg ( .D(
        new_AGEMA_signal_3750), .CK(clk), .Q(new_AGEMA_signal_3751) );
  DFF_X1 new_AGEMA_reg_buffer_1867_s_current_state_reg ( .D(
        new_AGEMA_signal_3754), .CK(clk), .Q(new_AGEMA_signal_3755) );
  DFF_X1 new_AGEMA_reg_buffer_1871_s_current_state_reg ( .D(
        new_AGEMA_signal_3758), .CK(clk), .Q(new_AGEMA_signal_3759) );
  DFF_X1 new_AGEMA_reg_buffer_1875_s_current_state_reg ( .D(
        new_AGEMA_signal_3762), .CK(clk), .Q(new_AGEMA_signal_3763) );
  DFF_X1 new_AGEMA_reg_buffer_1879_s_current_state_reg ( .D(
        new_AGEMA_signal_3766), .CK(clk), .Q(new_AGEMA_signal_3767) );
  DFF_X1 new_AGEMA_reg_buffer_1883_s_current_state_reg ( .D(
        new_AGEMA_signal_3770), .CK(clk), .Q(new_AGEMA_signal_3771) );
  DFF_X1 new_AGEMA_reg_buffer_1887_s_current_state_reg ( .D(
        new_AGEMA_signal_3774), .CK(clk), .Q(new_AGEMA_signal_3775) );
  DFF_X1 new_AGEMA_reg_buffer_1891_s_current_state_reg ( .D(
        new_AGEMA_signal_3778), .CK(clk), .Q(new_AGEMA_signal_3779) );
  DFF_X1 new_AGEMA_reg_buffer_1895_s_current_state_reg ( .D(
        new_AGEMA_signal_3782), .CK(clk), .Q(new_AGEMA_signal_3783) );
  DFF_X1 new_AGEMA_reg_buffer_1899_s_current_state_reg ( .D(
        new_AGEMA_signal_3786), .CK(clk), .Q(new_AGEMA_signal_3787) );
  DFF_X1 new_AGEMA_reg_buffer_1903_s_current_state_reg ( .D(
        new_AGEMA_signal_3790), .CK(clk), .Q(new_AGEMA_signal_3791) );
  DFF_X1 new_AGEMA_reg_buffer_1907_s_current_state_reg ( .D(
        new_AGEMA_signal_3794), .CK(clk), .Q(new_AGEMA_signal_3795) );
  DFF_X1 new_AGEMA_reg_buffer_1911_s_current_state_reg ( .D(
        new_AGEMA_signal_3798), .CK(clk), .Q(new_AGEMA_signal_3799) );
  DFF_X1 new_AGEMA_reg_buffer_1915_s_current_state_reg ( .D(
        new_AGEMA_signal_3802), .CK(clk), .Q(new_AGEMA_signal_3803) );
  DFF_X1 new_AGEMA_reg_buffer_1919_s_current_state_reg ( .D(
        new_AGEMA_signal_3806), .CK(clk), .Q(new_AGEMA_signal_3807) );
  DFF_X1 new_AGEMA_reg_buffer_1923_s_current_state_reg ( .D(
        new_AGEMA_signal_3810), .CK(clk), .Q(new_AGEMA_signal_3811) );
  DFF_X1 new_AGEMA_reg_buffer_1927_s_current_state_reg ( .D(
        new_AGEMA_signal_3814), .CK(clk), .Q(new_AGEMA_signal_3815) );
  DFF_X1 new_AGEMA_reg_buffer_1931_s_current_state_reg ( .D(
        new_AGEMA_signal_3818), .CK(clk), .Q(new_AGEMA_signal_3819) );
  DFF_X1 new_AGEMA_reg_buffer_1935_s_current_state_reg ( .D(
        new_AGEMA_signal_3822), .CK(clk), .Q(new_AGEMA_signal_3823) );
  DFF_X1 new_AGEMA_reg_buffer_1939_s_current_state_reg ( .D(
        new_AGEMA_signal_3826), .CK(clk), .Q(new_AGEMA_signal_3827) );
  DFF_X1 new_AGEMA_reg_buffer_1943_s_current_state_reg ( .D(
        new_AGEMA_signal_3830), .CK(clk), .Q(new_AGEMA_signal_3831) );
  DFF_X1 new_AGEMA_reg_buffer_1947_s_current_state_reg ( .D(
        new_AGEMA_signal_3834), .CK(clk), .Q(new_AGEMA_signal_3835) );
  DFF_X1 new_AGEMA_reg_buffer_1951_s_current_state_reg ( .D(
        new_AGEMA_signal_3838), .CK(clk), .Q(new_AGEMA_signal_3839) );
  DFF_X1 new_AGEMA_reg_buffer_1955_s_current_state_reg ( .D(
        new_AGEMA_signal_3842), .CK(clk), .Q(new_AGEMA_signal_3843) );
  DFF_X1 new_AGEMA_reg_buffer_1959_s_current_state_reg ( .D(
        new_AGEMA_signal_3846), .CK(clk), .Q(new_AGEMA_signal_3847) );
  DFF_X1 new_AGEMA_reg_buffer_1963_s_current_state_reg ( .D(
        new_AGEMA_signal_3850), .CK(clk), .Q(new_AGEMA_signal_3851) );
  DFF_X1 new_AGEMA_reg_buffer_1967_s_current_state_reg ( .D(
        new_AGEMA_signal_3854), .CK(clk), .Q(new_AGEMA_signal_3855) );
  DFF_X1 new_AGEMA_reg_buffer_1971_s_current_state_reg ( .D(
        new_AGEMA_signal_3858), .CK(clk), .Q(new_AGEMA_signal_3859) );
  DFF_X1 new_AGEMA_reg_buffer_1975_s_current_state_reg ( .D(
        new_AGEMA_signal_3862), .CK(clk), .Q(new_AGEMA_signal_3863) );
  DFF_X1 new_AGEMA_reg_buffer_1979_s_current_state_reg ( .D(
        new_AGEMA_signal_3866), .CK(clk), .Q(new_AGEMA_signal_3867) );
  DFF_X1 new_AGEMA_reg_buffer_1983_s_current_state_reg ( .D(
        new_AGEMA_signal_3870), .CK(clk), .Q(new_AGEMA_signal_3871) );
  DFF_X1 new_AGEMA_reg_buffer_1987_s_current_state_reg ( .D(
        new_AGEMA_signal_3874), .CK(clk), .Q(new_AGEMA_signal_3875) );
  DFF_X1 new_AGEMA_reg_buffer_1991_s_current_state_reg ( .D(
        new_AGEMA_signal_3878), .CK(clk), .Q(new_AGEMA_signal_3879) );
  DFF_X1 new_AGEMA_reg_buffer_1995_s_current_state_reg ( .D(
        new_AGEMA_signal_3882), .CK(clk), .Q(new_AGEMA_signal_3883) );
  DFF_X1 new_AGEMA_reg_buffer_1999_s_current_state_reg ( .D(
        new_AGEMA_signal_3886), .CK(clk), .Q(new_AGEMA_signal_3887) );
  DFF_X1 new_AGEMA_reg_buffer_2003_s_current_state_reg ( .D(
        new_AGEMA_signal_3890), .CK(clk), .Q(new_AGEMA_signal_3891) );
  DFF_X1 new_AGEMA_reg_buffer_2007_s_current_state_reg ( .D(
        new_AGEMA_signal_3894), .CK(clk), .Q(new_AGEMA_signal_3895) );
  DFF_X1 new_AGEMA_reg_buffer_2011_s_current_state_reg ( .D(
        new_AGEMA_signal_3898), .CK(clk), .Q(new_AGEMA_signal_3899) );
  DFF_X1 new_AGEMA_reg_buffer_2015_s_current_state_reg ( .D(
        new_AGEMA_signal_3902), .CK(clk), .Q(new_AGEMA_signal_3903) );
  DFF_X1 new_AGEMA_reg_buffer_2019_s_current_state_reg ( .D(
        new_AGEMA_signal_3906), .CK(clk), .Q(new_AGEMA_signal_3907) );
  DFF_X1 new_AGEMA_reg_buffer_2023_s_current_state_reg ( .D(
        new_AGEMA_signal_3910), .CK(clk), .Q(new_AGEMA_signal_3911) );
  DFF_X1 new_AGEMA_reg_buffer_2027_s_current_state_reg ( .D(
        new_AGEMA_signal_3914), .CK(clk), .Q(new_AGEMA_signal_3915) );
  DFF_X1 new_AGEMA_reg_buffer_2031_s_current_state_reg ( .D(
        new_AGEMA_signal_3918), .CK(clk), .Q(new_AGEMA_signal_3919) );
  DFF_X1 new_AGEMA_reg_buffer_2035_s_current_state_reg ( .D(
        new_AGEMA_signal_3922), .CK(clk), .Q(new_AGEMA_signal_3923) );
  DFF_X1 new_AGEMA_reg_buffer_2039_s_current_state_reg ( .D(
        new_AGEMA_signal_3926), .CK(clk), .Q(new_AGEMA_signal_3927) );
  DFF_X1 new_AGEMA_reg_buffer_2043_s_current_state_reg ( .D(
        new_AGEMA_signal_3930), .CK(clk), .Q(new_AGEMA_signal_3931) );
  DFF_X1 new_AGEMA_reg_buffer_2047_s_current_state_reg ( .D(
        new_AGEMA_signal_3934), .CK(clk), .Q(new_AGEMA_signal_3935) );
  DFF_X1 new_AGEMA_reg_buffer_2051_s_current_state_reg ( .D(
        new_AGEMA_signal_3938), .CK(clk), .Q(new_AGEMA_signal_3939) );
  DFF_X1 new_AGEMA_reg_buffer_2055_s_current_state_reg ( .D(
        new_AGEMA_signal_3942), .CK(clk), .Q(new_AGEMA_signal_3943) );
  DFF_X1 new_AGEMA_reg_buffer_2059_s_current_state_reg ( .D(
        new_AGEMA_signal_3946), .CK(clk), .Q(new_AGEMA_signal_3947) );
  DFF_X1 new_AGEMA_reg_buffer_2063_s_current_state_reg ( .D(
        new_AGEMA_signal_3950), .CK(clk), .Q(new_AGEMA_signal_3951) );
  DFF_X1 new_AGEMA_reg_buffer_2067_s_current_state_reg ( .D(
        new_AGEMA_signal_3954), .CK(clk), .Q(new_AGEMA_signal_3955) );
  DFF_X1 new_AGEMA_reg_buffer_2071_s_current_state_reg ( .D(
        new_AGEMA_signal_3958), .CK(clk), .Q(new_AGEMA_signal_3959) );
  DFF_X1 new_AGEMA_reg_buffer_2075_s_current_state_reg ( .D(
        new_AGEMA_signal_3962), .CK(clk), .Q(new_AGEMA_signal_3963) );
  DFF_X1 new_AGEMA_reg_buffer_2079_s_current_state_reg ( .D(
        new_AGEMA_signal_3966), .CK(clk), .Q(new_AGEMA_signal_3967) );
  DFF_X1 new_AGEMA_reg_buffer_2083_s_current_state_reg ( .D(
        new_AGEMA_signal_3970), .CK(clk), .Q(new_AGEMA_signal_3971) );
  DFF_X1 new_AGEMA_reg_buffer_2087_s_current_state_reg ( .D(
        new_AGEMA_signal_3974), .CK(clk), .Q(new_AGEMA_signal_3975) );
  DFF_X1 new_AGEMA_reg_buffer_2091_s_current_state_reg ( .D(
        new_AGEMA_signal_3978), .CK(clk), .Q(new_AGEMA_signal_3979) );
  DFF_X1 new_AGEMA_reg_buffer_2095_s_current_state_reg ( .D(
        new_AGEMA_signal_3982), .CK(clk), .Q(new_AGEMA_signal_3983) );
  DFF_X1 new_AGEMA_reg_buffer_2099_s_current_state_reg ( .D(
        new_AGEMA_signal_3986), .CK(clk), .Q(new_AGEMA_signal_3987) );
  DFF_X1 new_AGEMA_reg_buffer_2103_s_current_state_reg ( .D(
        new_AGEMA_signal_3990), .CK(clk), .Q(new_AGEMA_signal_3991) );
  DFF_X1 new_AGEMA_reg_buffer_2107_s_current_state_reg ( .D(
        new_AGEMA_signal_3994), .CK(clk), .Q(new_AGEMA_signal_3995) );
  DFF_X1 new_AGEMA_reg_buffer_2111_s_current_state_reg ( .D(
        new_AGEMA_signal_3998), .CK(clk), .Q(new_AGEMA_signal_3999) );
  DFF_X1 new_AGEMA_reg_buffer_2115_s_current_state_reg ( .D(
        new_AGEMA_signal_4002), .CK(clk), .Q(new_AGEMA_signal_4003) );
  DFF_X1 new_AGEMA_reg_buffer_2119_s_current_state_reg ( .D(
        new_AGEMA_signal_4006), .CK(clk), .Q(new_AGEMA_signal_4007) );
  DFF_X1 new_AGEMA_reg_buffer_2123_s_current_state_reg ( .D(
        new_AGEMA_signal_4010), .CK(clk), .Q(new_AGEMA_signal_4011) );
  DFF_X1 new_AGEMA_reg_buffer_2127_s_current_state_reg ( .D(
        new_AGEMA_signal_4014), .CK(clk), .Q(new_AGEMA_signal_4015) );
  DFF_X1 new_AGEMA_reg_buffer_2131_s_current_state_reg ( .D(
        new_AGEMA_signal_4018), .CK(clk), .Q(new_AGEMA_signal_4019) );
  DFF_X1 new_AGEMA_reg_buffer_2135_s_current_state_reg ( .D(
        new_AGEMA_signal_4022), .CK(clk), .Q(new_AGEMA_signal_4023) );
  DFF_X1 new_AGEMA_reg_buffer_2139_s_current_state_reg ( .D(
        new_AGEMA_signal_4026), .CK(clk), .Q(new_AGEMA_signal_4027) );
  DFF_X1 new_AGEMA_reg_buffer_2143_s_current_state_reg ( .D(
        new_AGEMA_signal_4030), .CK(clk), .Q(new_AGEMA_signal_4031) );
  DFF_X1 new_AGEMA_reg_buffer_2147_s_current_state_reg ( .D(
        new_AGEMA_signal_4034), .CK(clk), .Q(new_AGEMA_signal_4035) );
  DFF_X1 new_AGEMA_reg_buffer_2151_s_current_state_reg ( .D(
        new_AGEMA_signal_4038), .CK(clk), .Q(new_AGEMA_signal_4039) );
  DFF_X1 new_AGEMA_reg_buffer_2155_s_current_state_reg ( .D(
        new_AGEMA_signal_4042), .CK(clk), .Q(new_AGEMA_signal_4043) );
  DFF_X1 new_AGEMA_reg_buffer_2159_s_current_state_reg ( .D(
        new_AGEMA_signal_4046), .CK(clk), .Q(new_AGEMA_signal_4047) );
  DFF_X1 new_AGEMA_reg_buffer_2163_s_current_state_reg ( .D(
        new_AGEMA_signal_4050), .CK(clk), .Q(new_AGEMA_signal_4051) );
  DFF_X1 new_AGEMA_reg_buffer_2167_s_current_state_reg ( .D(
        new_AGEMA_signal_4054), .CK(clk), .Q(new_AGEMA_signal_4055) );
  DFF_X1 new_AGEMA_reg_buffer_2171_s_current_state_reg ( .D(
        new_AGEMA_signal_4058), .CK(clk), .Q(new_AGEMA_signal_4059) );
  DFF_X1 new_AGEMA_reg_buffer_2175_s_current_state_reg ( .D(
        new_AGEMA_signal_4062), .CK(clk), .Q(new_AGEMA_signal_4063) );
  DFF_X1 new_AGEMA_reg_buffer_2179_s_current_state_reg ( .D(
        new_AGEMA_signal_4066), .CK(clk), .Q(new_AGEMA_signal_4067) );
  DFF_X1 new_AGEMA_reg_buffer_2183_s_current_state_reg ( .D(
        new_AGEMA_signal_4070), .CK(clk), .Q(new_AGEMA_signal_4071) );
  DFF_X1 new_AGEMA_reg_buffer_2187_s_current_state_reg ( .D(
        new_AGEMA_signal_4074), .CK(clk), .Q(new_AGEMA_signal_4075) );
  DFF_X1 new_AGEMA_reg_buffer_2191_s_current_state_reg ( .D(
        new_AGEMA_signal_4078), .CK(clk), .Q(new_AGEMA_signal_4079) );
  DFF_X1 new_AGEMA_reg_buffer_2195_s_current_state_reg ( .D(
        new_AGEMA_signal_4082), .CK(clk), .Q(new_AGEMA_signal_4083) );
  DFF_X1 new_AGEMA_reg_buffer_2199_s_current_state_reg ( .D(
        new_AGEMA_signal_4086), .CK(clk), .Q(new_AGEMA_signal_4087) );
  DFF_X1 new_AGEMA_reg_buffer_2203_s_current_state_reg ( .D(
        new_AGEMA_signal_4090), .CK(clk), .Q(new_AGEMA_signal_4091) );
  DFF_X1 new_AGEMA_reg_buffer_2207_s_current_state_reg ( .D(
        new_AGEMA_signal_4094), .CK(clk), .Q(new_AGEMA_signal_4095) );
  DFF_X1 new_AGEMA_reg_buffer_2211_s_current_state_reg ( .D(
        new_AGEMA_signal_4098), .CK(clk), .Q(new_AGEMA_signal_4099) );
  DFF_X1 new_AGEMA_reg_buffer_2215_s_current_state_reg ( .D(
        new_AGEMA_signal_4102), .CK(clk), .Q(new_AGEMA_signal_4103) );
  DFF_X1 new_AGEMA_reg_buffer_2219_s_current_state_reg ( .D(
        new_AGEMA_signal_4106), .CK(clk), .Q(new_AGEMA_signal_4107) );
  DFF_X1 new_AGEMA_reg_buffer_2223_s_current_state_reg ( .D(
        new_AGEMA_signal_4110), .CK(clk), .Q(new_AGEMA_signal_4111) );
  DFF_X1 new_AGEMA_reg_buffer_2227_s_current_state_reg ( .D(
        new_AGEMA_signal_4114), .CK(clk), .Q(new_AGEMA_signal_4115) );
  DFF_X1 new_AGEMA_reg_buffer_2231_s_current_state_reg ( .D(
        new_AGEMA_signal_4118), .CK(clk), .Q(new_AGEMA_signal_4119) );
  DFF_X1 new_AGEMA_reg_buffer_2235_s_current_state_reg ( .D(
        new_AGEMA_signal_4122), .CK(clk), .Q(new_AGEMA_signal_4123) );
  DFF_X1 new_AGEMA_reg_buffer_2239_s_current_state_reg ( .D(
        new_AGEMA_signal_4126), .CK(clk), .Q(new_AGEMA_signal_4127) );
  DFF_X1 new_AGEMA_reg_buffer_2243_s_current_state_reg ( .D(
        new_AGEMA_signal_4130), .CK(clk), .Q(new_AGEMA_signal_4131) );
  DFF_X1 new_AGEMA_reg_buffer_2246_s_current_state_reg ( .D(
        new_AGEMA_signal_4133), .CK(clk), .Q(new_AGEMA_signal_4134) );
  DFF_X1 new_AGEMA_reg_buffer_2249_s_current_state_reg ( .D(
        new_AGEMA_signal_4136), .CK(clk), .Q(new_AGEMA_signal_4137) );
  DFF_X1 new_AGEMA_reg_buffer_2252_s_current_state_reg ( .D(
        new_AGEMA_signal_4139), .CK(clk), .Q(new_AGEMA_signal_4140) );
  DFF_X1 new_AGEMA_reg_buffer_2255_s_current_state_reg ( .D(
        new_AGEMA_signal_4142), .CK(clk), .Q(new_AGEMA_signal_4143) );
  DFF_X1 new_AGEMA_reg_buffer_2258_s_current_state_reg ( .D(
        new_AGEMA_signal_4145), .CK(clk), .Q(new_AGEMA_signal_4146) );
  DFF_X1 new_AGEMA_reg_buffer_2261_s_current_state_reg ( .D(
        new_AGEMA_signal_4148), .CK(clk), .Q(new_AGEMA_signal_4149) );
  DFF_X1 new_AGEMA_reg_buffer_2264_s_current_state_reg ( .D(
        new_AGEMA_signal_4151), .CK(clk), .Q(new_AGEMA_signal_4152) );
  DFF_X1 new_AGEMA_reg_buffer_2267_s_current_state_reg ( .D(
        new_AGEMA_signal_4154), .CK(clk), .Q(new_AGEMA_signal_4155) );
  DFF_X1 new_AGEMA_reg_buffer_2270_s_current_state_reg ( .D(
        new_AGEMA_signal_4157), .CK(clk), .Q(new_AGEMA_signal_4158) );
  DFF_X1 new_AGEMA_reg_buffer_2273_s_current_state_reg ( .D(
        new_AGEMA_signal_4160), .CK(clk), .Q(new_AGEMA_signal_4161) );
  DFF_X1 new_AGEMA_reg_buffer_2276_s_current_state_reg ( .D(
        new_AGEMA_signal_4163), .CK(clk), .Q(new_AGEMA_signal_4164) );
  DFF_X1 new_AGEMA_reg_buffer_2279_s_current_state_reg ( .D(
        new_AGEMA_signal_4166), .CK(clk), .Q(new_AGEMA_signal_4167) );
  DFF_X1 new_AGEMA_reg_buffer_2282_s_current_state_reg ( .D(
        new_AGEMA_signal_4169), .CK(clk), .Q(new_AGEMA_signal_4170) );
  DFF_X1 new_AGEMA_reg_buffer_2285_s_current_state_reg ( .D(
        new_AGEMA_signal_4172), .CK(clk), .Q(new_AGEMA_signal_4173) );
  DFF_X1 new_AGEMA_reg_buffer_2288_s_current_state_reg ( .D(
        new_AGEMA_signal_4175), .CK(clk), .Q(new_AGEMA_signal_4176) );
  DFF_X1 new_AGEMA_reg_buffer_2291_s_current_state_reg ( .D(
        new_AGEMA_signal_4178), .CK(clk), .Q(new_AGEMA_signal_4179) );
  DFF_X1 new_AGEMA_reg_buffer_2294_s_current_state_reg ( .D(
        new_AGEMA_signal_4181), .CK(clk), .Q(new_AGEMA_signal_4182) );
  DFF_X1 new_AGEMA_reg_buffer_2297_s_current_state_reg ( .D(
        new_AGEMA_signal_4184), .CK(clk), .Q(new_AGEMA_signal_4185) );
  DFF_X1 new_AGEMA_reg_buffer_2300_s_current_state_reg ( .D(
        new_AGEMA_signal_4187), .CK(clk), .Q(new_AGEMA_signal_4188) );
  DFF_X1 new_AGEMA_reg_buffer_2303_s_current_state_reg ( .D(
        new_AGEMA_signal_4190), .CK(clk), .Q(new_AGEMA_signal_4191) );
  DFF_X1 new_AGEMA_reg_buffer_2306_s_current_state_reg ( .D(
        new_AGEMA_signal_4193), .CK(clk), .Q(new_AGEMA_signal_4194) );
  DFF_X1 new_AGEMA_reg_buffer_2309_s_current_state_reg ( .D(
        new_AGEMA_signal_4196), .CK(clk), .Q(new_AGEMA_signal_4197) );
  DFF_X1 new_AGEMA_reg_buffer_2312_s_current_state_reg ( .D(
        new_AGEMA_signal_4199), .CK(clk), .Q(new_AGEMA_signal_4200) );
  DFF_X1 new_AGEMA_reg_buffer_2315_s_current_state_reg ( .D(
        new_AGEMA_signal_4202), .CK(clk), .Q(new_AGEMA_signal_4203) );
  DFF_X1 new_AGEMA_reg_buffer_2318_s_current_state_reg ( .D(
        new_AGEMA_signal_4205), .CK(clk), .Q(new_AGEMA_signal_4206) );
  DFF_X1 new_AGEMA_reg_buffer_2321_s_current_state_reg ( .D(
        new_AGEMA_signal_4208), .CK(clk), .Q(new_AGEMA_signal_4209) );
  DFF_X1 new_AGEMA_reg_buffer_2324_s_current_state_reg ( .D(
        new_AGEMA_signal_4211), .CK(clk), .Q(new_AGEMA_signal_4212) );
  DFF_X1 new_AGEMA_reg_buffer_2327_s_current_state_reg ( .D(
        new_AGEMA_signal_4214), .CK(clk), .Q(new_AGEMA_signal_4215) );
  DFF_X1 new_AGEMA_reg_buffer_2330_s_current_state_reg ( .D(
        new_AGEMA_signal_4217), .CK(clk), .Q(new_AGEMA_signal_4218) );
  DFF_X1 new_AGEMA_reg_buffer_2333_s_current_state_reg ( .D(
        new_AGEMA_signal_4220), .CK(clk), .Q(new_AGEMA_signal_4221) );
  DFF_X1 new_AGEMA_reg_buffer_2336_s_current_state_reg ( .D(
        new_AGEMA_signal_4223), .CK(clk), .Q(new_AGEMA_signal_4224) );
  DFF_X1 new_AGEMA_reg_buffer_2339_s_current_state_reg ( .D(
        new_AGEMA_signal_4226), .CK(clk), .Q(new_AGEMA_signal_4227) );
  DFF_X1 new_AGEMA_reg_buffer_2342_s_current_state_reg ( .D(
        new_AGEMA_signal_4229), .CK(clk), .Q(new_AGEMA_signal_4230) );
  DFF_X1 new_AGEMA_reg_buffer_2345_s_current_state_reg ( .D(
        new_AGEMA_signal_4232), .CK(clk), .Q(new_AGEMA_signal_4233) );
  DFF_X1 new_AGEMA_reg_buffer_2348_s_current_state_reg ( .D(
        new_AGEMA_signal_4235), .CK(clk), .Q(new_AGEMA_signal_4236) );
  DFF_X1 new_AGEMA_reg_buffer_2351_s_current_state_reg ( .D(
        new_AGEMA_signal_4238), .CK(clk), .Q(new_AGEMA_signal_4239) );
  DFF_X1 new_AGEMA_reg_buffer_2355_s_current_state_reg ( .D(
        new_AGEMA_signal_4242), .CK(clk), .Q(new_AGEMA_signal_4243) );
  DFF_X1 new_AGEMA_reg_buffer_2359_s_current_state_reg ( .D(
        new_AGEMA_signal_4246), .CK(clk), .Q(new_AGEMA_signal_4247) );
  DFF_X1 new_AGEMA_reg_buffer_2363_s_current_state_reg ( .D(
        new_AGEMA_signal_4250), .CK(clk), .Q(new_AGEMA_signal_4251) );
  DFF_X1 new_AGEMA_reg_buffer_2367_s_current_state_reg ( .D(
        new_AGEMA_signal_4254), .CK(clk), .Q(new_AGEMA_signal_4255) );
  DFF_X1 new_AGEMA_reg_buffer_2371_s_current_state_reg ( .D(
        new_AGEMA_signal_4258), .CK(clk), .Q(new_AGEMA_signal_4259) );
  DFF_X1 new_AGEMA_reg_buffer_2375_s_current_state_reg ( .D(
        new_AGEMA_signal_4262), .CK(clk), .Q(new_AGEMA_signal_4263) );
  DFF_X1 new_AGEMA_reg_buffer_2379_s_current_state_reg ( .D(
        new_AGEMA_signal_4266), .CK(clk), .Q(new_AGEMA_signal_4267) );
  DFF_X1 new_AGEMA_reg_buffer_2383_s_current_state_reg ( .D(
        new_AGEMA_signal_4270), .CK(clk), .Q(new_AGEMA_signal_4271) );
  DFF_X1 new_AGEMA_reg_buffer_2387_s_current_state_reg ( .D(
        new_AGEMA_signal_4274), .CK(clk), .Q(new_AGEMA_signal_4275) );
  DFF_X1 new_AGEMA_reg_buffer_2391_s_current_state_reg ( .D(
        new_AGEMA_signal_4278), .CK(clk), .Q(new_AGEMA_signal_4279) );
  DFF_X1 new_AGEMA_reg_buffer_2395_s_current_state_reg ( .D(
        new_AGEMA_signal_4282), .CK(clk), .Q(new_AGEMA_signal_4283) );
  DFF_X1 new_AGEMA_reg_buffer_2399_s_current_state_reg ( .D(
        new_AGEMA_signal_4286), .CK(clk), .Q(new_AGEMA_signal_4287) );
  DFF_X1 new_AGEMA_reg_buffer_2403_s_current_state_reg ( .D(
        new_AGEMA_signal_4290), .CK(clk), .Q(new_AGEMA_signal_4291) );
  DFF_X1 new_AGEMA_reg_buffer_2407_s_current_state_reg ( .D(
        new_AGEMA_signal_4294), .CK(clk), .Q(new_AGEMA_signal_4295) );
  DFF_X1 new_AGEMA_reg_buffer_2411_s_current_state_reg ( .D(
        new_AGEMA_signal_4298), .CK(clk), .Q(new_AGEMA_signal_4299) );
  DFF_X1 new_AGEMA_reg_buffer_2415_s_current_state_reg ( .D(
        new_AGEMA_signal_4302), .CK(clk), .Q(new_AGEMA_signal_4303) );
  DFF_X1 new_AGEMA_reg_buffer_2419_s_current_state_reg ( .D(
        new_AGEMA_signal_4306), .CK(clk), .Q(new_AGEMA_signal_4307) );
  DFF_X1 new_AGEMA_reg_buffer_2423_s_current_state_reg ( .D(
        new_AGEMA_signal_4310), .CK(clk), .Q(new_AGEMA_signal_4311) );
  DFF_X1 new_AGEMA_reg_buffer_2427_s_current_state_reg ( .D(
        new_AGEMA_signal_4314), .CK(clk), .Q(new_AGEMA_signal_4315) );
  DFF_X1 new_AGEMA_reg_buffer_2431_s_current_state_reg ( .D(
        new_AGEMA_signal_4318), .CK(clk), .Q(new_AGEMA_signal_4319) );
  DFF_X1 new_AGEMA_reg_buffer_2435_s_current_state_reg ( .D(
        new_AGEMA_signal_4322), .CK(clk), .Q(new_AGEMA_signal_4323) );
  DFF_X1 new_AGEMA_reg_buffer_2439_s_current_state_reg ( .D(
        new_AGEMA_signal_4326), .CK(clk), .Q(new_AGEMA_signal_4327) );
  DFF_X1 new_AGEMA_reg_buffer_2443_s_current_state_reg ( .D(
        new_AGEMA_signal_4330), .CK(clk), .Q(new_AGEMA_signal_4331) );
  DFF_X1 new_AGEMA_reg_buffer_2447_s_current_state_reg ( .D(
        new_AGEMA_signal_4334), .CK(clk), .Q(new_AGEMA_signal_4335) );
  DFF_X1 new_AGEMA_reg_buffer_2451_s_current_state_reg ( .D(
        new_AGEMA_signal_4338), .CK(clk), .Q(new_AGEMA_signal_4339) );
  DFF_X1 new_AGEMA_reg_buffer_2455_s_current_state_reg ( .D(
        new_AGEMA_signal_4342), .CK(clk), .Q(new_AGEMA_signal_4343) );
  DFF_X1 new_AGEMA_reg_buffer_2459_s_current_state_reg ( .D(
        new_AGEMA_signal_4346), .CK(clk), .Q(new_AGEMA_signal_4347) );
  DFF_X1 new_AGEMA_reg_buffer_2463_s_current_state_reg ( .D(
        new_AGEMA_signal_4350), .CK(clk), .Q(new_AGEMA_signal_4351) );
  DFF_X1 new_AGEMA_reg_buffer_2467_s_current_state_reg ( .D(
        new_AGEMA_signal_4354), .CK(clk), .Q(new_AGEMA_signal_4355) );
  DFF_X1 new_AGEMA_reg_buffer_2471_s_current_state_reg ( .D(
        new_AGEMA_signal_4358), .CK(clk), .Q(new_AGEMA_signal_4359) );
  DFF_X1 new_AGEMA_reg_buffer_2475_s_current_state_reg ( .D(
        new_AGEMA_signal_4362), .CK(clk), .Q(new_AGEMA_signal_4363) );
  DFF_X1 new_AGEMA_reg_buffer_2479_s_current_state_reg ( .D(
        new_AGEMA_signal_4366), .CK(clk), .Q(new_AGEMA_signal_4367) );
  DFF_X1 new_AGEMA_reg_buffer_2483_s_current_state_reg ( .D(
        new_AGEMA_signal_4370), .CK(clk), .Q(new_AGEMA_signal_4371) );
  DFF_X1 new_AGEMA_reg_buffer_2487_s_current_state_reg ( .D(
        new_AGEMA_signal_4374), .CK(clk), .Q(new_AGEMA_signal_4375) );
  DFF_X1 new_AGEMA_reg_buffer_2491_s_current_state_reg ( .D(
        new_AGEMA_signal_4378), .CK(clk), .Q(new_AGEMA_signal_4379) );
  DFF_X1 new_AGEMA_reg_buffer_2495_s_current_state_reg ( .D(
        new_AGEMA_signal_4382), .CK(clk), .Q(new_AGEMA_signal_4383) );
  DFF_X1 new_AGEMA_reg_buffer_2499_s_current_state_reg ( .D(
        new_AGEMA_signal_4386), .CK(clk), .Q(new_AGEMA_signal_4387) );
  DFF_X1 new_AGEMA_reg_buffer_2503_s_current_state_reg ( .D(
        new_AGEMA_signal_4390), .CK(clk), .Q(new_AGEMA_signal_4391) );
  DFF_X1 new_AGEMA_reg_buffer_2507_s_current_state_reg ( .D(
        new_AGEMA_signal_4394), .CK(clk), .Q(new_AGEMA_signal_4395) );
  DFF_X1 new_AGEMA_reg_buffer_2511_s_current_state_reg ( .D(
        new_AGEMA_signal_4398), .CK(clk), .Q(new_AGEMA_signal_4399) );
  DFF_X1 new_AGEMA_reg_buffer_2515_s_current_state_reg ( .D(
        new_AGEMA_signal_4402), .CK(clk), .Q(new_AGEMA_signal_4403) );
  DFF_X1 new_AGEMA_reg_buffer_2519_s_current_state_reg ( .D(
        new_AGEMA_signal_4406), .CK(clk), .Q(new_AGEMA_signal_4407) );
  DFF_X1 new_AGEMA_reg_buffer_2523_s_current_state_reg ( .D(
        new_AGEMA_signal_4410), .CK(clk), .Q(new_AGEMA_signal_4411) );
  DFF_X1 new_AGEMA_reg_buffer_2527_s_current_state_reg ( .D(
        new_AGEMA_signal_4414), .CK(clk), .Q(new_AGEMA_signal_4415) );
  DFF_X1 new_AGEMA_reg_buffer_2531_s_current_state_reg ( .D(
        new_AGEMA_signal_4418), .CK(clk), .Q(new_AGEMA_signal_4419) );
  DFF_X1 new_AGEMA_reg_buffer_2535_s_current_state_reg ( .D(
        new_AGEMA_signal_4422), .CK(clk), .Q(new_AGEMA_signal_4423) );
  DFF_X1 new_AGEMA_reg_buffer_2539_s_current_state_reg ( .D(
        new_AGEMA_signal_4426), .CK(clk), .Q(new_AGEMA_signal_4427) );
  DFF_X1 new_AGEMA_reg_buffer_2543_s_current_state_reg ( .D(
        new_AGEMA_signal_4430), .CK(clk), .Q(new_AGEMA_signal_4431) );
  DFF_X1 new_AGEMA_reg_buffer_2547_s_current_state_reg ( .D(
        new_AGEMA_signal_4434), .CK(clk), .Q(new_AGEMA_signal_4435) );
  DFF_X1 new_AGEMA_reg_buffer_2551_s_current_state_reg ( .D(
        new_AGEMA_signal_4438), .CK(clk), .Q(new_AGEMA_signal_4439) );
  DFF_X1 new_AGEMA_reg_buffer_2555_s_current_state_reg ( .D(
        new_AGEMA_signal_4442), .CK(clk), .Q(new_AGEMA_signal_4443) );
  DFF_X1 new_AGEMA_reg_buffer_2559_s_current_state_reg ( .D(
        new_AGEMA_signal_4446), .CK(clk), .Q(new_AGEMA_signal_4447) );
  DFF_X1 new_AGEMA_reg_buffer_2563_s_current_state_reg ( .D(
        new_AGEMA_signal_4450), .CK(clk), .Q(new_AGEMA_signal_4451) );
  DFF_X1 new_AGEMA_reg_buffer_2567_s_current_state_reg ( .D(
        new_AGEMA_signal_4454), .CK(clk), .Q(new_AGEMA_signal_4455) );
  DFF_X1 new_AGEMA_reg_buffer_2571_s_current_state_reg ( .D(
        new_AGEMA_signal_4458), .CK(clk), .Q(new_AGEMA_signal_4459) );
  DFF_X1 new_AGEMA_reg_buffer_2575_s_current_state_reg ( .D(
        new_AGEMA_signal_4462), .CK(clk), .Q(new_AGEMA_signal_4463) );
  DFF_X1 new_AGEMA_reg_buffer_2579_s_current_state_reg ( .D(
        new_AGEMA_signal_4466), .CK(clk), .Q(new_AGEMA_signal_4467) );
  DFF_X1 new_AGEMA_reg_buffer_2583_s_current_state_reg ( .D(
        new_AGEMA_signal_4470), .CK(clk), .Q(new_AGEMA_signal_4471) );
  DFF_X1 new_AGEMA_reg_buffer_2587_s_current_state_reg ( .D(
        new_AGEMA_signal_4474), .CK(clk), .Q(new_AGEMA_signal_4475) );
  DFF_X1 new_AGEMA_reg_buffer_2591_s_current_state_reg ( .D(
        new_AGEMA_signal_4478), .CK(clk), .Q(new_AGEMA_signal_4479) );
  DFF_X1 new_AGEMA_reg_buffer_2595_s_current_state_reg ( .D(
        new_AGEMA_signal_4482), .CK(clk), .Q(new_AGEMA_signal_4483) );
  DFF_X1 new_AGEMA_reg_buffer_2599_s_current_state_reg ( .D(
        new_AGEMA_signal_4486), .CK(clk), .Q(new_AGEMA_signal_4487) );
  DFF_X1 new_AGEMA_reg_buffer_2603_s_current_state_reg ( .D(
        new_AGEMA_signal_4490), .CK(clk), .Q(new_AGEMA_signal_4491) );
  DFF_X1 new_AGEMA_reg_buffer_2607_s_current_state_reg ( .D(
        new_AGEMA_signal_4494), .CK(clk), .Q(new_AGEMA_signal_4495) );
  DFF_X1 new_AGEMA_reg_buffer_2611_s_current_state_reg ( .D(
        new_AGEMA_signal_4498), .CK(clk), .Q(new_AGEMA_signal_4499) );
  DFF_X1 new_AGEMA_reg_buffer_2615_s_current_state_reg ( .D(
        new_AGEMA_signal_4502), .CK(clk), .Q(new_AGEMA_signal_4503) );
  DFF_X1 new_AGEMA_reg_buffer_2619_s_current_state_reg ( .D(
        new_AGEMA_signal_4506), .CK(clk), .Q(new_AGEMA_signal_4507) );
  DFF_X1 new_AGEMA_reg_buffer_2623_s_current_state_reg ( .D(
        new_AGEMA_signal_4510), .CK(clk), .Q(new_AGEMA_signal_4511) );
  DFF_X1 new_AGEMA_reg_buffer_2627_s_current_state_reg ( .D(
        new_AGEMA_signal_4514), .CK(clk), .Q(new_AGEMA_signal_4515) );
  DFF_X1 new_AGEMA_reg_buffer_2631_s_current_state_reg ( .D(
        new_AGEMA_signal_4518), .CK(clk), .Q(new_AGEMA_signal_4519) );
  DFF_X1 new_AGEMA_reg_buffer_2635_s_current_state_reg ( .D(
        new_AGEMA_signal_4522), .CK(clk), .Q(new_AGEMA_signal_4523) );
  DFF_X1 new_AGEMA_reg_buffer_2639_s_current_state_reg ( .D(
        new_AGEMA_signal_4526), .CK(clk), .Q(new_AGEMA_signal_4527) );
  DFF_X1 new_AGEMA_reg_buffer_2643_s_current_state_reg ( .D(
        new_AGEMA_signal_4530), .CK(clk), .Q(new_AGEMA_signal_4531) );
  DFF_X1 new_AGEMA_reg_buffer_2647_s_current_state_reg ( .D(
        new_AGEMA_signal_4534), .CK(clk), .Q(new_AGEMA_signal_4535) );
  DFF_X1 new_AGEMA_reg_buffer_2651_s_current_state_reg ( .D(
        new_AGEMA_signal_4538), .CK(clk), .Q(new_AGEMA_signal_4539) );
  DFF_X1 new_AGEMA_reg_buffer_2655_s_current_state_reg ( .D(
        new_AGEMA_signal_4542), .CK(clk), .Q(new_AGEMA_signal_4543) );
  DFF_X1 new_AGEMA_reg_buffer_2659_s_current_state_reg ( .D(
        new_AGEMA_signal_4546), .CK(clk), .Q(new_AGEMA_signal_4547) );
  DFF_X1 new_AGEMA_reg_buffer_2663_s_current_state_reg ( .D(
        new_AGEMA_signal_4550), .CK(clk), .Q(new_AGEMA_signal_4551) );
  DFF_X1 new_AGEMA_reg_buffer_2667_s_current_state_reg ( .D(
        new_AGEMA_signal_4554), .CK(clk), .Q(new_AGEMA_signal_4555) );
  DFF_X1 new_AGEMA_reg_buffer_2671_s_current_state_reg ( .D(
        new_AGEMA_signal_4558), .CK(clk), .Q(new_AGEMA_signal_4559) );
  DFF_X1 new_AGEMA_reg_buffer_2675_s_current_state_reg ( .D(
        new_AGEMA_signal_4562), .CK(clk), .Q(new_AGEMA_signal_4563) );
  DFF_X1 new_AGEMA_reg_buffer_2679_s_current_state_reg ( .D(
        new_AGEMA_signal_4566), .CK(clk), .Q(new_AGEMA_signal_4567) );
  DFF_X1 new_AGEMA_reg_buffer_2683_s_current_state_reg ( .D(
        new_AGEMA_signal_4570), .CK(clk), .Q(new_AGEMA_signal_4571) );
  DFF_X1 new_AGEMA_reg_buffer_2687_s_current_state_reg ( .D(
        new_AGEMA_signal_4574), .CK(clk), .Q(new_AGEMA_signal_4575) );
  DFF_X1 new_AGEMA_reg_buffer_2691_s_current_state_reg ( .D(
        new_AGEMA_signal_4578), .CK(clk), .Q(new_AGEMA_signal_4579) );
  DFF_X1 new_AGEMA_reg_buffer_2695_s_current_state_reg ( .D(
        new_AGEMA_signal_4582), .CK(clk), .Q(new_AGEMA_signal_4583) );
  DFF_X1 new_AGEMA_reg_buffer_2699_s_current_state_reg ( .D(
        new_AGEMA_signal_4586), .CK(clk), .Q(new_AGEMA_signal_4587) );
  DFF_X1 new_AGEMA_reg_buffer_2703_s_current_state_reg ( .D(
        new_AGEMA_signal_4590), .CK(clk), .Q(new_AGEMA_signal_4591) );
  DFF_X1 new_AGEMA_reg_buffer_2707_s_current_state_reg ( .D(
        new_AGEMA_signal_4594), .CK(clk), .Q(new_AGEMA_signal_4595) );
  DFF_X1 new_AGEMA_reg_buffer_2711_s_current_state_reg ( .D(
        new_AGEMA_signal_4598), .CK(clk), .Q(new_AGEMA_signal_4599) );
  DFF_X1 new_AGEMA_reg_buffer_2715_s_current_state_reg ( .D(
        new_AGEMA_signal_4602), .CK(clk), .Q(new_AGEMA_signal_4603) );
  DFF_X1 new_AGEMA_reg_buffer_2719_s_current_state_reg ( .D(
        new_AGEMA_signal_4606), .CK(clk), .Q(new_AGEMA_signal_4607) );
  DFF_X1 new_AGEMA_reg_buffer_2723_s_current_state_reg ( .D(
        new_AGEMA_signal_4610), .CK(clk), .Q(new_AGEMA_signal_4611) );
  DFF_X1 new_AGEMA_reg_buffer_2727_s_current_state_reg ( .D(
        new_AGEMA_signal_4614), .CK(clk), .Q(new_AGEMA_signal_4615) );
  DFF_X1 new_AGEMA_reg_buffer_2731_s_current_state_reg ( .D(
        new_AGEMA_signal_4618), .CK(clk), .Q(new_AGEMA_signal_4619) );
  DFF_X1 new_AGEMA_reg_buffer_2735_s_current_state_reg ( .D(
        new_AGEMA_signal_4622), .CK(clk), .Q(new_AGEMA_signal_4623) );
  DFF_X1 new_AGEMA_reg_buffer_2739_s_current_state_reg ( .D(
        new_AGEMA_signal_4626), .CK(clk), .Q(new_AGEMA_signal_4627) );
  DFF_X1 new_AGEMA_reg_buffer_2743_s_current_state_reg ( .D(
        new_AGEMA_signal_4630), .CK(clk), .Q(new_AGEMA_signal_4631) );
  DFF_X1 new_AGEMA_reg_buffer_2747_s_current_state_reg ( .D(
        new_AGEMA_signal_4634), .CK(clk), .Q(new_AGEMA_signal_4635) );
  DFF_X1 new_AGEMA_reg_buffer_2751_s_current_state_reg ( .D(
        new_AGEMA_signal_4638), .CK(clk), .Q(new_AGEMA_signal_4639) );
  DFF_X1 new_AGEMA_reg_buffer_2755_s_current_state_reg ( .D(
        new_AGEMA_signal_4642), .CK(clk), .Q(new_AGEMA_signal_4643) );
  DFF_X1 new_AGEMA_reg_buffer_2759_s_current_state_reg ( .D(
        new_AGEMA_signal_4646), .CK(clk), .Q(new_AGEMA_signal_4647) );
  DFF_X1 new_AGEMA_reg_buffer_2763_s_current_state_reg ( .D(
        new_AGEMA_signal_4650), .CK(clk), .Q(new_AGEMA_signal_4651) );
  DFF_X1 new_AGEMA_reg_buffer_2767_s_current_state_reg ( .D(
        new_AGEMA_signal_4654), .CK(clk), .Q(new_AGEMA_signal_4655) );
  DFF_X1 new_AGEMA_reg_buffer_2771_s_current_state_reg ( .D(
        new_AGEMA_signal_4658), .CK(clk), .Q(new_AGEMA_signal_4659) );
  DFF_X1 new_AGEMA_reg_buffer_2775_s_current_state_reg ( .D(
        new_AGEMA_signal_4662), .CK(clk), .Q(new_AGEMA_signal_4663) );
  DFF_X1 new_AGEMA_reg_buffer_2779_s_current_state_reg ( .D(
        new_AGEMA_signal_4666), .CK(clk), .Q(new_AGEMA_signal_4667) );
  DFF_X1 new_AGEMA_reg_buffer_2783_s_current_state_reg ( .D(
        new_AGEMA_signal_4670), .CK(clk), .Q(new_AGEMA_signal_4671) );
  DFF_X1 new_AGEMA_reg_buffer_2787_s_current_state_reg ( .D(
        new_AGEMA_signal_4674), .CK(clk), .Q(new_AGEMA_signal_4675) );
  DFF_X1 new_AGEMA_reg_buffer_2791_s_current_state_reg ( .D(
        new_AGEMA_signal_4678), .CK(clk), .Q(new_AGEMA_signal_4679) );
  DFF_X1 new_AGEMA_reg_buffer_2795_s_current_state_reg ( .D(
        new_AGEMA_signal_4682), .CK(clk), .Q(new_AGEMA_signal_4683) );
  DFF_X1 new_AGEMA_reg_buffer_2799_s_current_state_reg ( .D(
        new_AGEMA_signal_4686), .CK(clk), .Q(new_AGEMA_signal_4687) );
  DFF_X1 new_AGEMA_reg_buffer_2803_s_current_state_reg ( .D(
        new_AGEMA_signal_4690), .CK(clk), .Q(new_AGEMA_signal_4691) );
  DFF_X1 new_AGEMA_reg_buffer_2807_s_current_state_reg ( .D(
        new_AGEMA_signal_4694), .CK(clk), .Q(new_AGEMA_signal_4695) );
  DFF_X1 new_AGEMA_reg_buffer_2811_s_current_state_reg ( .D(
        new_AGEMA_signal_4698), .CK(clk), .Q(new_AGEMA_signal_4699) );
  DFF_X1 new_AGEMA_reg_buffer_2815_s_current_state_reg ( .D(
        new_AGEMA_signal_4702), .CK(clk), .Q(new_AGEMA_signal_4703) );
  DFF_X1 new_AGEMA_reg_buffer_2819_s_current_state_reg ( .D(
        new_AGEMA_signal_4706), .CK(clk), .Q(new_AGEMA_signal_4707) );
  DFF_X1 new_AGEMA_reg_buffer_2823_s_current_state_reg ( .D(
        new_AGEMA_signal_4710), .CK(clk), .Q(new_AGEMA_signal_4711) );
  DFF_X1 new_AGEMA_reg_buffer_2827_s_current_state_reg ( .D(
        new_AGEMA_signal_4714), .CK(clk), .Q(new_AGEMA_signal_4715) );
  DFF_X1 new_AGEMA_reg_buffer_2831_s_current_state_reg ( .D(
        new_AGEMA_signal_4718), .CK(clk), .Q(new_AGEMA_signal_4719) );
  DFF_X1 new_AGEMA_reg_buffer_2835_s_current_state_reg ( .D(
        new_AGEMA_signal_4722), .CK(clk), .Q(new_AGEMA_signal_4723) );
  DFF_X1 new_AGEMA_reg_buffer_2839_s_current_state_reg ( .D(
        new_AGEMA_signal_4726), .CK(clk), .Q(new_AGEMA_signal_4727) );
  DFF_X1 new_AGEMA_reg_buffer_2843_s_current_state_reg ( .D(
        new_AGEMA_signal_4730), .CK(clk), .Q(new_AGEMA_signal_4731) );
  DFF_X1 new_AGEMA_reg_buffer_2847_s_current_state_reg ( .D(
        new_AGEMA_signal_4734), .CK(clk), .Q(new_AGEMA_signal_4735) );
  DFF_X1 new_AGEMA_reg_buffer_2851_s_current_state_reg ( .D(
        new_AGEMA_signal_4738), .CK(clk), .Q(new_AGEMA_signal_4739) );
  DFF_X1 new_AGEMA_reg_buffer_2855_s_current_state_reg ( .D(
        new_AGEMA_signal_4742), .CK(clk), .Q(new_AGEMA_signal_4743) );
  DFF_X1 new_AGEMA_reg_buffer_2859_s_current_state_reg ( .D(
        new_AGEMA_signal_4746), .CK(clk), .Q(new_AGEMA_signal_4747) );
  DFF_X1 new_AGEMA_reg_buffer_2863_s_current_state_reg ( .D(
        new_AGEMA_signal_4750), .CK(clk), .Q(new_AGEMA_signal_4751) );
  DFF_X1 new_AGEMA_reg_buffer_2867_s_current_state_reg ( .D(
        new_AGEMA_signal_4754), .CK(clk), .Q(new_AGEMA_signal_4755) );
  DFF_X1 new_AGEMA_reg_buffer_2871_s_current_state_reg ( .D(
        new_AGEMA_signal_4758), .CK(clk), .Q(new_AGEMA_signal_4759) );
  DFF_X1 new_AGEMA_reg_buffer_2875_s_current_state_reg ( .D(
        new_AGEMA_signal_4762), .CK(clk), .Q(new_AGEMA_signal_4763) );
  DFF_X1 new_AGEMA_reg_buffer_2879_s_current_state_reg ( .D(
        new_AGEMA_signal_4766), .CK(clk), .Q(new_AGEMA_signal_4767) );
  DFF_X1 new_AGEMA_reg_buffer_2883_s_current_state_reg ( .D(
        new_AGEMA_signal_4770), .CK(clk), .Q(new_AGEMA_signal_4771) );
  DFF_X1 new_AGEMA_reg_buffer_2887_s_current_state_reg ( .D(
        new_AGEMA_signal_4774), .CK(clk), .Q(new_AGEMA_signal_4775) );
  DFF_X1 new_AGEMA_reg_buffer_2891_s_current_state_reg ( .D(
        new_AGEMA_signal_4778), .CK(clk), .Q(new_AGEMA_signal_4779) );
  DFF_X1 new_AGEMA_reg_buffer_2895_s_current_state_reg ( .D(
        new_AGEMA_signal_4782), .CK(clk), .Q(new_AGEMA_signal_4783) );
  DFF_X1 new_AGEMA_reg_buffer_2899_s_current_state_reg ( .D(
        new_AGEMA_signal_4786), .CK(clk), .Q(new_AGEMA_signal_4787) );
  DFF_X1 new_AGEMA_reg_buffer_2903_s_current_state_reg ( .D(
        new_AGEMA_signal_4790), .CK(clk), .Q(new_AGEMA_signal_4791) );
  DFF_X1 new_AGEMA_reg_buffer_2907_s_current_state_reg ( .D(
        new_AGEMA_signal_4794), .CK(clk), .Q(new_AGEMA_signal_4795) );
  DFF_X1 new_AGEMA_reg_buffer_2911_s_current_state_reg ( .D(
        new_AGEMA_signal_4798), .CK(clk), .Q(new_AGEMA_signal_4799) );
  DFF_X1 new_AGEMA_reg_buffer_2915_s_current_state_reg ( .D(
        new_AGEMA_signal_4802), .CK(clk), .Q(new_AGEMA_signal_4803) );
  DFF_X1 new_AGEMA_reg_buffer_2919_s_current_state_reg ( .D(
        new_AGEMA_signal_4806), .CK(clk), .Q(new_AGEMA_signal_4807) );
  DFF_X1 new_AGEMA_reg_buffer_2923_s_current_state_reg ( .D(
        new_AGEMA_signal_4810), .CK(clk), .Q(new_AGEMA_signal_4811) );
  DFF_X1 new_AGEMA_reg_buffer_2927_s_current_state_reg ( .D(
        new_AGEMA_signal_4814), .CK(clk), .Q(new_AGEMA_signal_4815) );
  DFF_X1 new_AGEMA_reg_buffer_2931_s_current_state_reg ( .D(
        new_AGEMA_signal_4818), .CK(clk), .Q(new_AGEMA_signal_4819) );
  DFF_X1 new_AGEMA_reg_buffer_2935_s_current_state_reg ( .D(
        new_AGEMA_signal_4822), .CK(clk), .Q(new_AGEMA_signal_4823) );
  DFF_X1 new_AGEMA_reg_buffer_2939_s_current_state_reg ( .D(
        new_AGEMA_signal_4826), .CK(clk), .Q(new_AGEMA_signal_4827) );
  DFF_X1 new_AGEMA_reg_buffer_2943_s_current_state_reg ( .D(
        new_AGEMA_signal_4830), .CK(clk), .Q(new_AGEMA_signal_4831) );
  DFF_X1 new_AGEMA_reg_buffer_2947_s_current_state_reg ( .D(
        new_AGEMA_signal_4834), .CK(clk), .Q(new_AGEMA_signal_4835) );
  DFF_X1 new_AGEMA_reg_buffer_2951_s_current_state_reg ( .D(
        new_AGEMA_signal_4838), .CK(clk), .Q(new_AGEMA_signal_4839) );
  DFF_X1 new_AGEMA_reg_buffer_2955_s_current_state_reg ( .D(
        new_AGEMA_signal_4842), .CK(clk), .Q(new_AGEMA_signal_4843) );
  DFF_X1 new_AGEMA_reg_buffer_2959_s_current_state_reg ( .D(
        new_AGEMA_signal_4846), .CK(clk), .Q(new_AGEMA_signal_4847) );
  DFF_X1 new_AGEMA_reg_buffer_2963_s_current_state_reg ( .D(
        new_AGEMA_signal_4850), .CK(clk), .Q(new_AGEMA_signal_4851) );
  DFF_X1 new_AGEMA_reg_buffer_2967_s_current_state_reg ( .D(
        new_AGEMA_signal_4854), .CK(clk), .Q(new_AGEMA_signal_4855) );
  DFF_X1 new_AGEMA_reg_buffer_2971_s_current_state_reg ( .D(
        new_AGEMA_signal_4858), .CK(clk), .Q(new_AGEMA_signal_4859) );
  DFF_X1 new_AGEMA_reg_buffer_2975_s_current_state_reg ( .D(
        new_AGEMA_signal_4862), .CK(clk), .Q(new_AGEMA_signal_4863) );
  DFF_X1 new_AGEMA_reg_buffer_2979_s_current_state_reg ( .D(
        new_AGEMA_signal_4866), .CK(clk), .Q(new_AGEMA_signal_4867) );
  DFF_X1 new_AGEMA_reg_buffer_2983_s_current_state_reg ( .D(
        new_AGEMA_signal_4870), .CK(clk), .Q(new_AGEMA_signal_4871) );
  DFF_X1 new_AGEMA_reg_buffer_2987_s_current_state_reg ( .D(
        new_AGEMA_signal_4874), .CK(clk), .Q(new_AGEMA_signal_4875) );
  DFF_X1 new_AGEMA_reg_buffer_2991_s_current_state_reg ( .D(
        new_AGEMA_signal_4878), .CK(clk), .Q(new_AGEMA_signal_4879) );
  DFF_X1 new_AGEMA_reg_buffer_2995_s_current_state_reg ( .D(
        new_AGEMA_signal_4882), .CK(clk), .Q(new_AGEMA_signal_4883) );
  DFF_X1 new_AGEMA_reg_buffer_2999_s_current_state_reg ( .D(
        new_AGEMA_signal_4886), .CK(clk), .Q(new_AGEMA_signal_4887) );
  DFF_X1 new_AGEMA_reg_buffer_3003_s_current_state_reg ( .D(
        new_AGEMA_signal_4890), .CK(clk), .Q(new_AGEMA_signal_4891) );
  DFF_X1 new_AGEMA_reg_buffer_3007_s_current_state_reg ( .D(
        new_AGEMA_signal_4894), .CK(clk), .Q(new_AGEMA_signal_4895) );
  DFF_X1 new_AGEMA_reg_buffer_3011_s_current_state_reg ( .D(
        new_AGEMA_signal_4898), .CK(clk), .Q(new_AGEMA_signal_4899) );
  DFF_X1 new_AGEMA_reg_buffer_3015_s_current_state_reg ( .D(
        new_AGEMA_signal_4902), .CK(clk), .Q(new_AGEMA_signal_4903) );
  DFF_X1 new_AGEMA_reg_buffer_3019_s_current_state_reg ( .D(
        new_AGEMA_signal_4906), .CK(clk), .Q(new_AGEMA_signal_4907) );
  DFF_X1 new_AGEMA_reg_buffer_3023_s_current_state_reg ( .D(
        new_AGEMA_signal_4910), .CK(clk), .Q(new_AGEMA_signal_4911) );
  DFF_X1 new_AGEMA_reg_buffer_3027_s_current_state_reg ( .D(
        new_AGEMA_signal_4914), .CK(clk), .Q(new_AGEMA_signal_4915) );
  DFF_X1 new_AGEMA_reg_buffer_3031_s_current_state_reg ( .D(
        new_AGEMA_signal_4918), .CK(clk), .Q(new_AGEMA_signal_4919) );
  DFF_X1 new_AGEMA_reg_buffer_3035_s_current_state_reg ( .D(
        new_AGEMA_signal_4922), .CK(clk), .Q(new_AGEMA_signal_4923) );
  DFF_X1 new_AGEMA_reg_buffer_3039_s_current_state_reg ( .D(
        new_AGEMA_signal_4926), .CK(clk), .Q(new_AGEMA_signal_4927) );
  DFF_X1 new_AGEMA_reg_buffer_3043_s_current_state_reg ( .D(
        new_AGEMA_signal_4930), .CK(clk), .Q(new_AGEMA_signal_4931) );
  DFF_X1 new_AGEMA_reg_buffer_3047_s_current_state_reg ( .D(
        new_AGEMA_signal_4934), .CK(clk), .Q(new_AGEMA_signal_4935) );
  DFF_X1 new_AGEMA_reg_buffer_3051_s_current_state_reg ( .D(
        new_AGEMA_signal_4938), .CK(clk), .Q(new_AGEMA_signal_4939) );
  DFF_X1 new_AGEMA_reg_buffer_3055_s_current_state_reg ( .D(
        new_AGEMA_signal_4942), .CK(clk), .Q(new_AGEMA_signal_4943) );
  DFF_X1 new_AGEMA_reg_buffer_3059_s_current_state_reg ( .D(
        new_AGEMA_signal_4946), .CK(clk), .Q(new_AGEMA_signal_4947) );
  DFF_X1 new_AGEMA_reg_buffer_3063_s_current_state_reg ( .D(
        new_AGEMA_signal_4950), .CK(clk), .Q(new_AGEMA_signal_4951) );
  DFF_X1 new_AGEMA_reg_buffer_3067_s_current_state_reg ( .D(
        new_AGEMA_signal_4954), .CK(clk), .Q(new_AGEMA_signal_4955) );
  DFF_X1 new_AGEMA_reg_buffer_3071_s_current_state_reg ( .D(
        new_AGEMA_signal_4958), .CK(clk), .Q(new_AGEMA_signal_4959) );
  DFF_X1 new_AGEMA_reg_buffer_3075_s_current_state_reg ( .D(
        new_AGEMA_signal_4962), .CK(clk), .Q(new_AGEMA_signal_4963) );
  DFF_X1 new_AGEMA_reg_buffer_3079_s_current_state_reg ( .D(
        new_AGEMA_signal_4966), .CK(clk), .Q(new_AGEMA_signal_4967) );
  DFF_X1 new_AGEMA_reg_buffer_3083_s_current_state_reg ( .D(
        new_AGEMA_signal_4970), .CK(clk), .Q(new_AGEMA_signal_4971) );
  DFF_X1 new_AGEMA_reg_buffer_3087_s_current_state_reg ( .D(
        new_AGEMA_signal_4974), .CK(clk), .Q(new_AGEMA_signal_4975) );
  DFF_X1 new_AGEMA_reg_buffer_3091_s_current_state_reg ( .D(
        new_AGEMA_signal_4978), .CK(clk), .Q(new_AGEMA_signal_4979) );
  DFF_X1 new_AGEMA_reg_buffer_3095_s_current_state_reg ( .D(
        new_AGEMA_signal_4982), .CK(clk), .Q(new_AGEMA_signal_4983) );
  DFF_X1 new_AGEMA_reg_buffer_3099_s_current_state_reg ( .D(
        new_AGEMA_signal_4986), .CK(clk), .Q(new_AGEMA_signal_4987) );
  DFF_X1 new_AGEMA_reg_buffer_3103_s_current_state_reg ( .D(
        new_AGEMA_signal_4990), .CK(clk), .Q(new_AGEMA_signal_4991) );
  DFF_X1 new_AGEMA_reg_buffer_3107_s_current_state_reg ( .D(
        new_AGEMA_signal_4994), .CK(clk), .Q(new_AGEMA_signal_4995) );
  DFF_X1 new_AGEMA_reg_buffer_3111_s_current_state_reg ( .D(
        new_AGEMA_signal_4998), .CK(clk), .Q(new_AGEMA_signal_4999) );
  DFF_X1 new_AGEMA_reg_buffer_3115_s_current_state_reg ( .D(
        new_AGEMA_signal_5002), .CK(clk), .Q(new_AGEMA_signal_5003) );
  DFF_X1 new_AGEMA_reg_buffer_3119_s_current_state_reg ( .D(
        new_AGEMA_signal_5006), .CK(clk), .Q(new_AGEMA_signal_5007) );
  DFF_X1 new_AGEMA_reg_buffer_3123_s_current_state_reg ( .D(
        new_AGEMA_signal_5010), .CK(clk), .Q(new_AGEMA_signal_5011) );
  DFF_X1 new_AGEMA_reg_buffer_3127_s_current_state_reg ( .D(
        new_AGEMA_signal_5014), .CK(clk), .Q(new_AGEMA_signal_5015) );
  DFF_X1 new_AGEMA_reg_buffer_3131_s_current_state_reg ( .D(
        new_AGEMA_signal_5018), .CK(clk), .Q(new_AGEMA_signal_5019) );
  DFF_X1 new_AGEMA_reg_buffer_3135_s_current_state_reg ( .D(
        new_AGEMA_signal_5022), .CK(clk), .Q(new_AGEMA_signal_5023) );
  DFF_X1 new_AGEMA_reg_buffer_3139_s_current_state_reg ( .D(
        new_AGEMA_signal_5026), .CK(clk), .Q(new_AGEMA_signal_5027) );
  DFF_X1 new_AGEMA_reg_buffer_3143_s_current_state_reg ( .D(
        new_AGEMA_signal_5030), .CK(clk), .Q(new_AGEMA_signal_5031) );
  DFF_X1 new_AGEMA_reg_buffer_3147_s_current_state_reg ( .D(
        new_AGEMA_signal_5034), .CK(clk), .Q(new_AGEMA_signal_5035) );
  DFF_X1 new_AGEMA_reg_buffer_3151_s_current_state_reg ( .D(
        new_AGEMA_signal_5038), .CK(clk), .Q(new_AGEMA_signal_5039) );
  DFF_X1 new_AGEMA_reg_buffer_3155_s_current_state_reg ( .D(
        new_AGEMA_signal_5042), .CK(clk), .Q(new_AGEMA_signal_5043) );
  DFF_X1 new_AGEMA_reg_buffer_3159_s_current_state_reg ( .D(
        new_AGEMA_signal_5046), .CK(clk), .Q(new_AGEMA_signal_5047) );
  DFF_X1 new_AGEMA_reg_buffer_3163_s_current_state_reg ( .D(
        new_AGEMA_signal_5050), .CK(clk), .Q(new_AGEMA_signal_5051) );
  DFF_X1 new_AGEMA_reg_buffer_3167_s_current_state_reg ( .D(
        new_AGEMA_signal_5054), .CK(clk), .Q(new_AGEMA_signal_5055) );
  DFF_X1 new_AGEMA_reg_buffer_3171_s_current_state_reg ( .D(
        new_AGEMA_signal_5058), .CK(clk), .Q(new_AGEMA_signal_5059) );
  DFF_X1 new_AGEMA_reg_buffer_3175_s_current_state_reg ( .D(
        new_AGEMA_signal_5062), .CK(clk), .Q(new_AGEMA_signal_5063) );
  DFF_X1 new_AGEMA_reg_buffer_3179_s_current_state_reg ( .D(
        new_AGEMA_signal_5066), .CK(clk), .Q(new_AGEMA_signal_5067) );
  DFF_X1 new_AGEMA_reg_buffer_3183_s_current_state_reg ( .D(
        new_AGEMA_signal_5070), .CK(clk), .Q(new_AGEMA_signal_5071) );
  DFF_X1 new_AGEMA_reg_buffer_3187_s_current_state_reg ( .D(
        new_AGEMA_signal_5074), .CK(clk), .Q(new_AGEMA_signal_5075) );
  DFF_X1 new_AGEMA_reg_buffer_3191_s_current_state_reg ( .D(
        new_AGEMA_signal_5078), .CK(clk), .Q(new_AGEMA_signal_5079) );
  DFF_X1 new_AGEMA_reg_buffer_3195_s_current_state_reg ( .D(
        new_AGEMA_signal_5082), .CK(clk), .Q(new_AGEMA_signal_5083) );
  DFF_X1 new_AGEMA_reg_buffer_3199_s_current_state_reg ( .D(
        new_AGEMA_signal_5086), .CK(clk), .Q(new_AGEMA_signal_5087) );
  DFF_X1 new_AGEMA_reg_buffer_3203_s_current_state_reg ( .D(
        new_AGEMA_signal_5090), .CK(clk), .Q(new_AGEMA_signal_5091) );
  DFF_X1 new_AGEMA_reg_buffer_3207_s_current_state_reg ( .D(
        new_AGEMA_signal_5094), .CK(clk), .Q(new_AGEMA_signal_5095) );
  DFF_X1 new_AGEMA_reg_buffer_3211_s_current_state_reg ( .D(
        new_AGEMA_signal_5098), .CK(clk), .Q(new_AGEMA_signal_5099) );
  DFF_X1 new_AGEMA_reg_buffer_3215_s_current_state_reg ( .D(
        new_AGEMA_signal_5102), .CK(clk), .Q(new_AGEMA_signal_5103) );
  DFF_X1 new_AGEMA_reg_buffer_3219_s_current_state_reg ( .D(
        new_AGEMA_signal_5106), .CK(clk), .Q(new_AGEMA_signal_5107) );
  DFF_X1 new_AGEMA_reg_buffer_3223_s_current_state_reg ( .D(
        new_AGEMA_signal_5110), .CK(clk), .Q(new_AGEMA_signal_5111) );
  DFF_X1 new_AGEMA_reg_buffer_3227_s_current_state_reg ( .D(
        new_AGEMA_signal_5114), .CK(clk), .Q(new_AGEMA_signal_5115) );
  DFF_X1 new_AGEMA_reg_buffer_3231_s_current_state_reg ( .D(
        new_AGEMA_signal_5118), .CK(clk), .Q(new_AGEMA_signal_5119) );
  DFF_X1 new_AGEMA_reg_buffer_3235_s_current_state_reg ( .D(
        new_AGEMA_signal_5122), .CK(clk), .Q(new_AGEMA_signal_5123) );
  DFF_X1 new_AGEMA_reg_buffer_3239_s_current_state_reg ( .D(
        new_AGEMA_signal_5126), .CK(clk), .Q(new_AGEMA_signal_5127) );
  DFF_X1 new_AGEMA_reg_buffer_3243_s_current_state_reg ( .D(
        new_AGEMA_signal_5130), .CK(clk), .Q(new_AGEMA_signal_5131) );
  DFF_X1 new_AGEMA_reg_buffer_3247_s_current_state_reg ( .D(
        new_AGEMA_signal_5134), .CK(clk), .Q(new_AGEMA_signal_5135) );
  DFF_X1 new_AGEMA_reg_buffer_3251_s_current_state_reg ( .D(
        new_AGEMA_signal_5138), .CK(clk), .Q(new_AGEMA_signal_5139) );
  DFF_X1 new_AGEMA_reg_buffer_3255_s_current_state_reg ( .D(
        new_AGEMA_signal_5142), .CK(clk), .Q(new_AGEMA_signal_5143) );
  DFF_X1 new_AGEMA_reg_buffer_3259_s_current_state_reg ( .D(
        new_AGEMA_signal_5146), .CK(clk), .Q(new_AGEMA_signal_5147) );
  DFF_X1 new_AGEMA_reg_buffer_3263_s_current_state_reg ( .D(
        new_AGEMA_signal_5150), .CK(clk), .Q(new_AGEMA_signal_5151) );
  DFF_X1 new_AGEMA_reg_buffer_3267_s_current_state_reg ( .D(
        new_AGEMA_signal_5154), .CK(clk), .Q(new_AGEMA_signal_5155) );
  DFF_X1 new_AGEMA_reg_buffer_3271_s_current_state_reg ( .D(
        new_AGEMA_signal_5158), .CK(clk), .Q(new_AGEMA_signal_5159) );
  DFF_X1 new_AGEMA_reg_buffer_3275_s_current_state_reg ( .D(
        new_AGEMA_signal_5162), .CK(clk), .Q(new_AGEMA_signal_5163) );
  DFF_X1 new_AGEMA_reg_buffer_3279_s_current_state_reg ( .D(
        new_AGEMA_signal_5166), .CK(clk), .Q(new_AGEMA_signal_5167) );
  DFF_X1 new_AGEMA_reg_buffer_3283_s_current_state_reg ( .D(
        new_AGEMA_signal_5170), .CK(clk), .Q(new_AGEMA_signal_5171) );
  DFF_X1 new_AGEMA_reg_buffer_3287_s_current_state_reg ( .D(
        new_AGEMA_signal_5174), .CK(clk), .Q(new_AGEMA_signal_5175) );
  DFF_X1 new_AGEMA_reg_buffer_3291_s_current_state_reg ( .D(
        new_AGEMA_signal_5178), .CK(clk), .Q(new_AGEMA_signal_5179) );
  DFF_X1 new_AGEMA_reg_buffer_3295_s_current_state_reg ( .D(
        new_AGEMA_signal_5182), .CK(clk), .Q(new_AGEMA_signal_5183) );
  DFF_X1 new_AGEMA_reg_buffer_3299_s_current_state_reg ( .D(
        new_AGEMA_signal_5186), .CK(clk), .Q(new_AGEMA_signal_5187) );
  DFF_X1 new_AGEMA_reg_buffer_3303_s_current_state_reg ( .D(
        new_AGEMA_signal_5190), .CK(clk), .Q(new_AGEMA_signal_5191) );
  DFF_X1 new_AGEMA_reg_buffer_3307_s_current_state_reg ( .D(
        new_AGEMA_signal_5194), .CK(clk), .Q(new_AGEMA_signal_5195) );
  DFF_X1 new_AGEMA_reg_buffer_3311_s_current_state_reg ( .D(
        new_AGEMA_signal_5198), .CK(clk), .Q(new_AGEMA_signal_5199) );
  DFF_X1 new_AGEMA_reg_buffer_3315_s_current_state_reg ( .D(
        new_AGEMA_signal_5202), .CK(clk), .Q(new_AGEMA_signal_5203) );
  DFF_X1 new_AGEMA_reg_buffer_3319_s_current_state_reg ( .D(
        new_AGEMA_signal_5206), .CK(clk), .Q(new_AGEMA_signal_5207) );
  DFF_X1 new_AGEMA_reg_buffer_3323_s_current_state_reg ( .D(
        new_AGEMA_signal_5210), .CK(clk), .Q(new_AGEMA_signal_5211) );
  DFF_X1 new_AGEMA_reg_buffer_3327_s_current_state_reg ( .D(
        new_AGEMA_signal_5214), .CK(clk), .Q(new_AGEMA_signal_5215) );
  DFF_X1 new_AGEMA_reg_buffer_3331_s_current_state_reg ( .D(
        new_AGEMA_signal_5218), .CK(clk), .Q(new_AGEMA_signal_5219) );
  DFF_X1 new_AGEMA_reg_buffer_3335_s_current_state_reg ( .D(
        new_AGEMA_signal_5222), .CK(clk), .Q(new_AGEMA_signal_5223) );
  DFF_X1 new_AGEMA_reg_buffer_3339_s_current_state_reg ( .D(
        new_AGEMA_signal_5226), .CK(clk), .Q(new_AGEMA_signal_5227) );
  DFF_X1 new_AGEMA_reg_buffer_3343_s_current_state_reg ( .D(
        new_AGEMA_signal_5230), .CK(clk), .Q(new_AGEMA_signal_5231) );
  DFF_X1 new_AGEMA_reg_buffer_3347_s_current_state_reg ( .D(
        new_AGEMA_signal_5234), .CK(clk), .Q(new_AGEMA_signal_5235) );
  DFF_X1 new_AGEMA_reg_buffer_3351_s_current_state_reg ( .D(
        new_AGEMA_signal_5238), .CK(clk), .Q(new_AGEMA_signal_5239) );
  DFF_X1 new_AGEMA_reg_buffer_3355_s_current_state_reg ( .D(
        new_AGEMA_signal_5242), .CK(clk), .Q(new_AGEMA_signal_5243) );
  DFF_X1 new_AGEMA_reg_buffer_3359_s_current_state_reg ( .D(
        new_AGEMA_signal_5246), .CK(clk), .Q(new_AGEMA_signal_5247) );
  DFF_X1 new_AGEMA_reg_buffer_3363_s_current_state_reg ( .D(
        new_AGEMA_signal_5250), .CK(clk), .Q(new_AGEMA_signal_5251) );
  DFF_X1 new_AGEMA_reg_buffer_3367_s_current_state_reg ( .D(
        new_AGEMA_signal_5254), .CK(clk), .Q(new_AGEMA_signal_5255) );
  DFF_X1 new_AGEMA_reg_buffer_3371_s_current_state_reg ( .D(
        new_AGEMA_signal_5258), .CK(clk), .Q(new_AGEMA_signal_5259) );
  DFF_X1 new_AGEMA_reg_buffer_3375_s_current_state_reg ( .D(
        new_AGEMA_signal_5262), .CK(clk), .Q(new_AGEMA_signal_5263) );
  DFF_X1 new_AGEMA_reg_buffer_3379_s_current_state_reg ( .D(
        new_AGEMA_signal_5266), .CK(clk), .Q(new_AGEMA_signal_5267) );
  DFF_X1 new_AGEMA_reg_buffer_3383_s_current_state_reg ( .D(
        new_AGEMA_signal_5270), .CK(clk), .Q(new_AGEMA_signal_5271) );
  DFF_X1 new_AGEMA_reg_buffer_3387_s_current_state_reg ( .D(
        new_AGEMA_signal_5274), .CK(clk), .Q(new_AGEMA_signal_5275) );
  DFF_X1 new_AGEMA_reg_buffer_3391_s_current_state_reg ( .D(
        new_AGEMA_signal_5278), .CK(clk), .Q(new_AGEMA_signal_5279) );
  DFF_X1 new_AGEMA_reg_buffer_3395_s_current_state_reg ( .D(
        new_AGEMA_signal_5282), .CK(clk), .Q(new_AGEMA_signal_5283) );
  DFF_X1 new_AGEMA_reg_buffer_3399_s_current_state_reg ( .D(
        new_AGEMA_signal_5286), .CK(clk), .Q(new_AGEMA_signal_5287) );
  DFF_X1 new_AGEMA_reg_buffer_3403_s_current_state_reg ( .D(
        new_AGEMA_signal_5290), .CK(clk), .Q(new_AGEMA_signal_5291) );
  DFF_X1 new_AGEMA_reg_buffer_3407_s_current_state_reg ( .D(
        new_AGEMA_signal_5294), .CK(clk), .Q(new_AGEMA_signal_5295) );
  DFF_X1 new_AGEMA_reg_buffer_3411_s_current_state_reg ( .D(
        new_AGEMA_signal_5298), .CK(clk), .Q(new_AGEMA_signal_5299) );
  DFF_X1 new_AGEMA_reg_buffer_3415_s_current_state_reg ( .D(
        new_AGEMA_signal_5302), .CK(clk), .Q(new_AGEMA_signal_5303) );
  DFF_X1 new_AGEMA_reg_buffer_3419_s_current_state_reg ( .D(
        new_AGEMA_signal_5306), .CK(clk), .Q(new_AGEMA_signal_5307) );
  DFF_X1 new_AGEMA_reg_buffer_3423_s_current_state_reg ( .D(
        new_AGEMA_signal_5310), .CK(clk), .Q(new_AGEMA_signal_5311) );
  DFF_X1 new_AGEMA_reg_buffer_3427_s_current_state_reg ( .D(
        new_AGEMA_signal_5314), .CK(clk), .Q(new_AGEMA_signal_5315) );
  DFF_X1 new_AGEMA_reg_buffer_3431_s_current_state_reg ( .D(
        new_AGEMA_signal_5318), .CK(clk), .Q(new_AGEMA_signal_5319) );
  DFF_X1 new_AGEMA_reg_buffer_3435_s_current_state_reg ( .D(
        new_AGEMA_signal_5322), .CK(clk), .Q(new_AGEMA_signal_5323) );
  DFF_X1 new_AGEMA_reg_buffer_3439_s_current_state_reg ( .D(
        new_AGEMA_signal_5326), .CK(clk), .Q(new_AGEMA_signal_5327) );
  DFF_X1 new_AGEMA_reg_buffer_3443_s_current_state_reg ( .D(
        new_AGEMA_signal_5330), .CK(clk), .Q(new_AGEMA_signal_5331) );
  DFF_X1 new_AGEMA_reg_buffer_3447_s_current_state_reg ( .D(
        new_AGEMA_signal_5334), .CK(clk), .Q(new_AGEMA_signal_5335) );
  DFF_X1 new_AGEMA_reg_buffer_3451_s_current_state_reg ( .D(
        new_AGEMA_signal_5338), .CK(clk), .Q(new_AGEMA_signal_5339) );
  DFF_X1 new_AGEMA_reg_buffer_3455_s_current_state_reg ( .D(
        new_AGEMA_signal_5342), .CK(clk), .Q(new_AGEMA_signal_5343) );
  DFF_X1 new_AGEMA_reg_buffer_3459_s_current_state_reg ( .D(
        new_AGEMA_signal_5346), .CK(clk), .Q(new_AGEMA_signal_5347) );
  DFF_X1 new_AGEMA_reg_buffer_3463_s_current_state_reg ( .D(
        new_AGEMA_signal_5350), .CK(clk), .Q(new_AGEMA_signal_5351) );
  DFF_X1 new_AGEMA_reg_buffer_3467_s_current_state_reg ( .D(
        new_AGEMA_signal_5354), .CK(clk), .Q(new_AGEMA_signal_5355) );
  DFF_X1 new_AGEMA_reg_buffer_3471_s_current_state_reg ( .D(
        new_AGEMA_signal_5358), .CK(clk), .Q(new_AGEMA_signal_5359) );
  DFF_X1 new_AGEMA_reg_buffer_3475_s_current_state_reg ( .D(
        new_AGEMA_signal_5362), .CK(clk), .Q(new_AGEMA_signal_5363) );
  DFF_X1 new_AGEMA_reg_buffer_3479_s_current_state_reg ( .D(
        new_AGEMA_signal_5366), .CK(clk), .Q(new_AGEMA_signal_5367) );
  DFF_X1 new_AGEMA_reg_buffer_3483_s_current_state_reg ( .D(
        new_AGEMA_signal_5370), .CK(clk), .Q(new_AGEMA_signal_5371) );
  DFF_X1 new_AGEMA_reg_buffer_3487_s_current_state_reg ( .D(
        new_AGEMA_signal_5374), .CK(clk), .Q(new_AGEMA_signal_5375) );
  DFF_X1 new_AGEMA_reg_buffer_3491_s_current_state_reg ( .D(
        new_AGEMA_signal_5378), .CK(clk), .Q(new_AGEMA_signal_5379) );
  DFF_X1 new_AGEMA_reg_buffer_3495_s_current_state_reg ( .D(
        new_AGEMA_signal_5382), .CK(clk), .Q(new_AGEMA_signal_5383) );
  DFF_X1 new_AGEMA_reg_buffer_3499_s_current_state_reg ( .D(
        new_AGEMA_signal_5386), .CK(clk), .Q(new_AGEMA_signal_5387) );
  DFF_X1 new_AGEMA_reg_buffer_3503_s_current_state_reg ( .D(
        new_AGEMA_signal_5390), .CK(clk), .Q(new_AGEMA_signal_5391) );
  DFF_X1 new_AGEMA_reg_buffer_3507_s_current_state_reg ( .D(
        new_AGEMA_signal_5394), .CK(clk), .Q(new_AGEMA_signal_5395) );
  DFF_X1 new_AGEMA_reg_buffer_3511_s_current_state_reg ( .D(
        new_AGEMA_signal_5398), .CK(clk), .Q(new_AGEMA_signal_5399) );
  DFF_X1 new_AGEMA_reg_buffer_3515_s_current_state_reg ( .D(
        new_AGEMA_signal_5402), .CK(clk), .Q(new_AGEMA_signal_5403) );
  DFF_X1 new_AGEMA_reg_buffer_3519_s_current_state_reg ( .D(
        new_AGEMA_signal_5406), .CK(clk), .Q(new_AGEMA_signal_5407) );
  DFF_X1 new_AGEMA_reg_buffer_3523_s_current_state_reg ( .D(
        new_AGEMA_signal_5410), .CK(clk), .Q(new_AGEMA_signal_5411) );
  DFF_X1 new_AGEMA_reg_buffer_3527_s_current_state_reg ( .D(
        new_AGEMA_signal_5414), .CK(clk), .Q(new_AGEMA_signal_5415) );
  DFF_X1 new_AGEMA_reg_buffer_3531_s_current_state_reg ( .D(
        new_AGEMA_signal_5418), .CK(clk), .Q(new_AGEMA_signal_5419) );
  DFF_X1 new_AGEMA_reg_buffer_3535_s_current_state_reg ( .D(
        new_AGEMA_signal_5422), .CK(clk), .Q(new_AGEMA_signal_5423) );
  DFF_X1 new_AGEMA_reg_buffer_3539_s_current_state_reg ( .D(
        new_AGEMA_signal_5426), .CK(clk), .Q(new_AGEMA_signal_5427) );
  DFF_X1 new_AGEMA_reg_buffer_3543_s_current_state_reg ( .D(
        new_AGEMA_signal_5430), .CK(clk), .Q(new_AGEMA_signal_5431) );
  DFF_X1 new_AGEMA_reg_buffer_3547_s_current_state_reg ( .D(
        new_AGEMA_signal_5434), .CK(clk), .Q(new_AGEMA_signal_5435) );
  DFF_X1 new_AGEMA_reg_buffer_3551_s_current_state_reg ( .D(
        new_AGEMA_signal_5438), .CK(clk), .Q(new_AGEMA_signal_5439) );
  DFF_X1 new_AGEMA_reg_buffer_3555_s_current_state_reg ( .D(
        new_AGEMA_signal_5442), .CK(clk), .Q(new_AGEMA_signal_5443) );
  DFF_X1 new_AGEMA_reg_buffer_3559_s_current_state_reg ( .D(
        new_AGEMA_signal_5446), .CK(clk), .Q(new_AGEMA_signal_5447) );
  DFF_X1 new_AGEMA_reg_buffer_3563_s_current_state_reg ( .D(
        new_AGEMA_signal_5450), .CK(clk), .Q(new_AGEMA_signal_5451) );
  DFF_X1 new_AGEMA_reg_buffer_3567_s_current_state_reg ( .D(
        new_AGEMA_signal_5454), .CK(clk), .Q(new_AGEMA_signal_5455) );
  DFF_X1 new_AGEMA_reg_buffer_3571_s_current_state_reg ( .D(
        new_AGEMA_signal_5458), .CK(clk), .Q(new_AGEMA_signal_5459) );
  DFF_X1 new_AGEMA_reg_buffer_3575_s_current_state_reg ( .D(
        new_AGEMA_signal_5462), .CK(clk), .Q(new_AGEMA_signal_5463) );
  DFF_X1 new_AGEMA_reg_buffer_3579_s_current_state_reg ( .D(
        new_AGEMA_signal_5466), .CK(clk), .Q(new_AGEMA_signal_5467) );
  DFF_X1 new_AGEMA_reg_buffer_3583_s_current_state_reg ( .D(
        new_AGEMA_signal_5470), .CK(clk), .Q(new_AGEMA_signal_5471) );
  DFF_X1 new_AGEMA_reg_buffer_3587_s_current_state_reg ( .D(
        new_AGEMA_signal_5474), .CK(clk), .Q(new_AGEMA_signal_5475) );
  DFF_X1 new_AGEMA_reg_buffer_3591_s_current_state_reg ( .D(
        new_AGEMA_signal_5478), .CK(clk), .Q(new_AGEMA_signal_5479) );
  DFF_X1 new_AGEMA_reg_buffer_3595_s_current_state_reg ( .D(
        new_AGEMA_signal_5482), .CK(clk), .Q(new_AGEMA_signal_5483) );
  DFF_X1 new_AGEMA_reg_buffer_3599_s_current_state_reg ( .D(
        new_AGEMA_signal_5486), .CK(clk), .Q(new_AGEMA_signal_5487) );
  DFF_X1 new_AGEMA_reg_buffer_3603_s_current_state_reg ( .D(
        new_AGEMA_signal_5490), .CK(clk), .Q(new_AGEMA_signal_5491) );
  DFF_X1 new_AGEMA_reg_buffer_3607_s_current_state_reg ( .D(
        new_AGEMA_signal_5494), .CK(clk), .Q(new_AGEMA_signal_5495) );
  DFF_X1 new_AGEMA_reg_buffer_3611_s_current_state_reg ( .D(
        new_AGEMA_signal_5498), .CK(clk), .Q(new_AGEMA_signal_5499) );
  DFF_X1 new_AGEMA_reg_buffer_3615_s_current_state_reg ( .D(
        new_AGEMA_signal_5502), .CK(clk), .Q(new_AGEMA_signal_5503) );
  DFF_X1 new_AGEMA_reg_buffer_3619_s_current_state_reg ( .D(
        new_AGEMA_signal_5506), .CK(clk), .Q(new_AGEMA_signal_5507) );
  DFF_X1 new_AGEMA_reg_buffer_3623_s_current_state_reg ( .D(
        new_AGEMA_signal_5510), .CK(clk), .Q(new_AGEMA_signal_5511) );
  DFF_X1 new_AGEMA_reg_buffer_3627_s_current_state_reg ( .D(
        new_AGEMA_signal_5514), .CK(clk), .Q(new_AGEMA_signal_5515) );
  DFF_X1 new_AGEMA_reg_buffer_3631_s_current_state_reg ( .D(
        new_AGEMA_signal_5518), .CK(clk), .Q(new_AGEMA_signal_5519) );
  DFF_X1 new_AGEMA_reg_buffer_3635_s_current_state_reg ( .D(
        new_AGEMA_signal_5522), .CK(clk), .Q(new_AGEMA_signal_5523) );
  DFF_X1 new_AGEMA_reg_buffer_3639_s_current_state_reg ( .D(
        new_AGEMA_signal_5526), .CK(clk), .Q(new_AGEMA_signal_5527) );
  DFF_X1 new_AGEMA_reg_buffer_3643_s_current_state_reg ( .D(
        new_AGEMA_signal_5530), .CK(clk), .Q(new_AGEMA_signal_5531) );
  DFF_X1 new_AGEMA_reg_buffer_3647_s_current_state_reg ( .D(
        new_AGEMA_signal_5534), .CK(clk), .Q(new_AGEMA_signal_5535) );
  DFF_X1 new_AGEMA_reg_buffer_3651_s_current_state_reg ( .D(
        new_AGEMA_signal_5538), .CK(clk), .Q(new_AGEMA_signal_5539) );
  DFF_X1 new_AGEMA_reg_buffer_3655_s_current_state_reg ( .D(
        new_AGEMA_signal_5542), .CK(clk), .Q(new_AGEMA_signal_5543) );
  DFF_X1 new_AGEMA_reg_buffer_3659_s_current_state_reg ( .D(
        new_AGEMA_signal_5546), .CK(clk), .Q(new_AGEMA_signal_5547) );
  DFF_X1 new_AGEMA_reg_buffer_3663_s_current_state_reg ( .D(
        new_AGEMA_signal_5550), .CK(clk), .Q(new_AGEMA_signal_5551) );
  DFF_X1 new_AGEMA_reg_buffer_3667_s_current_state_reg ( .D(
        new_AGEMA_signal_5554), .CK(clk), .Q(new_AGEMA_signal_5555) );
  DFF_X1 new_AGEMA_reg_buffer_3671_s_current_state_reg ( .D(
        new_AGEMA_signal_5558), .CK(clk), .Q(new_AGEMA_signal_5559) );
  DFF_X1 new_AGEMA_reg_buffer_3675_s_current_state_reg ( .D(
        new_AGEMA_signal_5562), .CK(clk), .Q(new_AGEMA_signal_5563) );
  DFF_X1 new_AGEMA_reg_buffer_3679_s_current_state_reg ( .D(
        new_AGEMA_signal_5566), .CK(clk), .Q(new_AGEMA_signal_5567) );
  DFF_X1 new_AGEMA_reg_buffer_3683_s_current_state_reg ( .D(
        new_AGEMA_signal_5570), .CK(clk), .Q(new_AGEMA_signal_5571) );
  DFF_X1 new_AGEMA_reg_buffer_3687_s_current_state_reg ( .D(
        new_AGEMA_signal_5574), .CK(clk), .Q(new_AGEMA_signal_5575) );
  DFF_X1 new_AGEMA_reg_buffer_3691_s_current_state_reg ( .D(
        new_AGEMA_signal_5578), .CK(clk), .Q(new_AGEMA_signal_5579) );
  DFF_X1 new_AGEMA_reg_buffer_3695_s_current_state_reg ( .D(
        new_AGEMA_signal_5582), .CK(clk), .Q(new_AGEMA_signal_5583) );
  DFF_X1 new_AGEMA_reg_buffer_3699_s_current_state_reg ( .D(
        new_AGEMA_signal_5586), .CK(clk), .Q(new_AGEMA_signal_5587) );
  DFF_X1 new_AGEMA_reg_buffer_3703_s_current_state_reg ( .D(
        new_AGEMA_signal_5590), .CK(clk), .Q(new_AGEMA_signal_5591) );
  DFF_X1 new_AGEMA_reg_buffer_3707_s_current_state_reg ( .D(
        new_AGEMA_signal_5594), .CK(clk), .Q(new_AGEMA_signal_5595) );
  DFF_X1 new_AGEMA_reg_buffer_3711_s_current_state_reg ( .D(
        new_AGEMA_signal_5598), .CK(clk), .Q(new_AGEMA_signal_5599) );
  DFF_X1 new_AGEMA_reg_buffer_3715_s_current_state_reg ( .D(
        new_AGEMA_signal_5602), .CK(clk), .Q(new_AGEMA_signal_5603) );
  DFF_X1 new_AGEMA_reg_buffer_3719_s_current_state_reg ( .D(
        new_AGEMA_signal_5606), .CK(clk), .Q(new_AGEMA_signal_5607) );
  DFF_X1 new_AGEMA_reg_buffer_3723_s_current_state_reg ( .D(
        new_AGEMA_signal_5610), .CK(clk), .Q(new_AGEMA_signal_5611) );
  DFF_X1 new_AGEMA_reg_buffer_3727_s_current_state_reg ( .D(
        new_AGEMA_signal_5614), .CK(clk), .Q(new_AGEMA_signal_5615) );
  DFF_X1 new_AGEMA_reg_buffer_3731_s_current_state_reg ( .D(
        new_AGEMA_signal_5618), .CK(clk), .Q(new_AGEMA_signal_5619) );
  DFF_X1 new_AGEMA_reg_buffer_3735_s_current_state_reg ( .D(
        new_AGEMA_signal_5622), .CK(clk), .Q(new_AGEMA_signal_5623) );
  DFF_X1 new_AGEMA_reg_buffer_3739_s_current_state_reg ( .D(
        new_AGEMA_signal_5626), .CK(clk), .Q(new_AGEMA_signal_5627) );
  DFF_X1 new_AGEMA_reg_buffer_3743_s_current_state_reg ( .D(
        new_AGEMA_signal_5630), .CK(clk), .Q(new_AGEMA_signal_5631) );
  DFF_X1 new_AGEMA_reg_buffer_3747_s_current_state_reg ( .D(
        new_AGEMA_signal_5634), .CK(clk), .Q(new_AGEMA_signal_5635) );
  DFF_X1 new_AGEMA_reg_buffer_3751_s_current_state_reg ( .D(
        new_AGEMA_signal_5638), .CK(clk), .Q(new_AGEMA_signal_5639) );
  DFF_X1 new_AGEMA_reg_buffer_3755_s_current_state_reg ( .D(
        new_AGEMA_signal_5642), .CK(clk), .Q(new_AGEMA_signal_5643) );
  DFF_X1 new_AGEMA_reg_buffer_3759_s_current_state_reg ( .D(
        new_AGEMA_signal_5646), .CK(clk), .Q(new_AGEMA_signal_5647) );
  DFF_X1 new_AGEMA_reg_buffer_3763_s_current_state_reg ( .D(
        new_AGEMA_signal_5650), .CK(clk), .Q(new_AGEMA_signal_5651) );
  DFF_X1 new_AGEMA_reg_buffer_3767_s_current_state_reg ( .D(
        new_AGEMA_signal_5654), .CK(clk), .Q(new_AGEMA_signal_5655) );
  DFF_X1 new_AGEMA_reg_buffer_3771_s_current_state_reg ( .D(
        new_AGEMA_signal_5658), .CK(clk), .Q(new_AGEMA_signal_5659) );
  DFF_X1 new_AGEMA_reg_buffer_3775_s_current_state_reg ( .D(
        new_AGEMA_signal_5662), .CK(clk), .Q(new_AGEMA_signal_5663) );
  DFF_X1 new_AGEMA_reg_buffer_3779_s_current_state_reg ( .D(
        new_AGEMA_signal_5666), .CK(clk), .Q(new_AGEMA_signal_5667) );
  DFF_X1 new_AGEMA_reg_buffer_3783_s_current_state_reg ( .D(
        new_AGEMA_signal_5670), .CK(clk), .Q(new_AGEMA_signal_5671) );
  DFF_X1 new_AGEMA_reg_buffer_3787_s_current_state_reg ( .D(
        new_AGEMA_signal_5674), .CK(clk), .Q(new_AGEMA_signal_5675) );
  DFF_X1 new_AGEMA_reg_buffer_3791_s_current_state_reg ( .D(
        new_AGEMA_signal_5678), .CK(clk), .Q(new_AGEMA_signal_5679) );
  DFF_X1 new_AGEMA_reg_buffer_3795_s_current_state_reg ( .D(
        new_AGEMA_signal_5682), .CK(clk), .Q(new_AGEMA_signal_5683) );
  DFF_X1 new_AGEMA_reg_buffer_3799_s_current_state_reg ( .D(
        new_AGEMA_signal_5686), .CK(clk), .Q(new_AGEMA_signal_5687) );
  DFF_X1 new_AGEMA_reg_buffer_3803_s_current_state_reg ( .D(
        new_AGEMA_signal_5690), .CK(clk), .Q(new_AGEMA_signal_5691) );
  DFF_X1 new_AGEMA_reg_buffer_3807_s_current_state_reg ( .D(
        new_AGEMA_signal_5694), .CK(clk), .Q(new_AGEMA_signal_5695) );
  DFF_X1 new_AGEMA_reg_buffer_3811_s_current_state_reg ( .D(
        new_AGEMA_signal_5698), .CK(clk), .Q(new_AGEMA_signal_5699) );
  DFF_X1 new_AGEMA_reg_buffer_3815_s_current_state_reg ( .D(
        new_AGEMA_signal_5702), .CK(clk), .Q(new_AGEMA_signal_5703) );
  DFF_X1 new_AGEMA_reg_buffer_3819_s_current_state_reg ( .D(
        new_AGEMA_signal_5706), .CK(clk), .Q(new_AGEMA_signal_5707) );
  DFF_X1 new_AGEMA_reg_buffer_3823_s_current_state_reg ( .D(
        new_AGEMA_signal_5710), .CK(clk), .Q(new_AGEMA_signal_5711) );
  DFF_X1 new_AGEMA_reg_buffer_3827_s_current_state_reg ( .D(
        new_AGEMA_signal_5714), .CK(clk), .Q(new_AGEMA_signal_5715) );
  DFF_X1 new_AGEMA_reg_buffer_3831_s_current_state_reg ( .D(
        new_AGEMA_signal_5718), .CK(clk), .Q(new_AGEMA_signal_5719) );
  DFF_X1 new_AGEMA_reg_buffer_3835_s_current_state_reg ( .D(
        new_AGEMA_signal_5722), .CK(clk), .Q(new_AGEMA_signal_5723) );
  DFF_X1 new_AGEMA_reg_buffer_3839_s_current_state_reg ( .D(
        new_AGEMA_signal_5726), .CK(clk), .Q(new_AGEMA_signal_5727) );
  DFF_X1 new_AGEMA_reg_buffer_3843_s_current_state_reg ( .D(
        new_AGEMA_signal_5730), .CK(clk), .Q(new_AGEMA_signal_5731) );
  DFF_X1 new_AGEMA_reg_buffer_3847_s_current_state_reg ( .D(
        new_AGEMA_signal_5734), .CK(clk), .Q(new_AGEMA_signal_5735) );
  DFF_X1 new_AGEMA_reg_buffer_3851_s_current_state_reg ( .D(
        new_AGEMA_signal_5738), .CK(clk), .Q(new_AGEMA_signal_5739) );
  DFF_X1 new_AGEMA_reg_buffer_3855_s_current_state_reg ( .D(
        new_AGEMA_signal_5742), .CK(clk), .Q(new_AGEMA_signal_5743) );
  DFF_X1 new_AGEMA_reg_buffer_3859_s_current_state_reg ( .D(
        new_AGEMA_signal_5746), .CK(clk), .Q(new_AGEMA_signal_5747) );
  DFF_X1 new_AGEMA_reg_buffer_3863_s_current_state_reg ( .D(
        new_AGEMA_signal_5750), .CK(clk), .Q(new_AGEMA_signal_5751) );
  DFF_X1 new_AGEMA_reg_buffer_3867_s_current_state_reg ( .D(
        new_AGEMA_signal_5754), .CK(clk), .Q(new_AGEMA_signal_5755) );
  DFF_X1 new_AGEMA_reg_buffer_3871_s_current_state_reg ( .D(
        new_AGEMA_signal_5758), .CK(clk), .Q(new_AGEMA_signal_5759) );
  DFF_X1 new_AGEMA_reg_buffer_3875_s_current_state_reg ( .D(
        new_AGEMA_signal_5762), .CK(clk), .Q(new_AGEMA_signal_5763) );
  DFF_X1 new_AGEMA_reg_buffer_3879_s_current_state_reg ( .D(
        new_AGEMA_signal_5766), .CK(clk), .Q(new_AGEMA_signal_5767) );
  DFF_X1 new_AGEMA_reg_buffer_3883_s_current_state_reg ( .D(
        new_AGEMA_signal_5770), .CK(clk), .Q(new_AGEMA_signal_5771) );
  DFF_X1 new_AGEMA_reg_buffer_3887_s_current_state_reg ( .D(
        new_AGEMA_signal_5774), .CK(clk), .Q(new_AGEMA_signal_5775) );
  DFF_X1 new_AGEMA_reg_buffer_3891_s_current_state_reg ( .D(
        new_AGEMA_signal_5778), .CK(clk), .Q(new_AGEMA_signal_5779) );
  DFF_X1 new_AGEMA_reg_buffer_3895_s_current_state_reg ( .D(
        new_AGEMA_signal_5782), .CK(clk), .Q(new_AGEMA_signal_5783) );
  DFF_X1 new_AGEMA_reg_buffer_3899_s_current_state_reg ( .D(
        new_AGEMA_signal_5786), .CK(clk), .Q(new_AGEMA_signal_5787) );
  DFF_X1 new_AGEMA_reg_buffer_3903_s_current_state_reg ( .D(
        new_AGEMA_signal_5790), .CK(clk), .Q(new_AGEMA_signal_5791) );
  DFF_X1 new_AGEMA_reg_buffer_3907_s_current_state_reg ( .D(
        new_AGEMA_signal_5794), .CK(clk), .Q(new_AGEMA_signal_5795) );
  DFF_X1 new_AGEMA_reg_buffer_3911_s_current_state_reg ( .D(
        new_AGEMA_signal_5798), .CK(clk), .Q(new_AGEMA_signal_5799) );
  DFF_X1 new_AGEMA_reg_buffer_3915_s_current_state_reg ( .D(
        new_AGEMA_signal_5802), .CK(clk), .Q(new_AGEMA_signal_5803) );
  DFF_X1 new_AGEMA_reg_buffer_3919_s_current_state_reg ( .D(
        new_AGEMA_signal_5806), .CK(clk), .Q(new_AGEMA_signal_5807) );
  DFF_X1 new_AGEMA_reg_buffer_3923_s_current_state_reg ( .D(
        new_AGEMA_signal_5810), .CK(clk), .Q(new_AGEMA_signal_5811) );
  DFF_X1 new_AGEMA_reg_buffer_3927_s_current_state_reg ( .D(
        new_AGEMA_signal_5814), .CK(clk), .Q(new_AGEMA_signal_5815) );
  DFF_X1 new_AGEMA_reg_buffer_3931_s_current_state_reg ( .D(
        new_AGEMA_signal_5818), .CK(clk), .Q(new_AGEMA_signal_5819) );
  DFF_X1 new_AGEMA_reg_buffer_3935_s_current_state_reg ( .D(
        new_AGEMA_signal_5822), .CK(clk), .Q(new_AGEMA_signal_5823) );
  DFF_X1 new_AGEMA_reg_buffer_3939_s_current_state_reg ( .D(
        new_AGEMA_signal_5826), .CK(clk), .Q(new_AGEMA_signal_5827) );
  DFF_X1 new_AGEMA_reg_buffer_3943_s_current_state_reg ( .D(
        new_AGEMA_signal_5830), .CK(clk), .Q(new_AGEMA_signal_5831) );
  DFF_X1 new_AGEMA_reg_buffer_3947_s_current_state_reg ( .D(
        new_AGEMA_signal_5834), .CK(clk), .Q(new_AGEMA_signal_5835) );
  DFF_X1 new_AGEMA_reg_buffer_3951_s_current_state_reg ( .D(
        new_AGEMA_signal_5838), .CK(clk), .Q(new_AGEMA_signal_5839) );
  DFF_X1 new_AGEMA_reg_buffer_3955_s_current_state_reg ( .D(
        new_AGEMA_signal_5842), .CK(clk), .Q(new_AGEMA_signal_5843) );
  DFF_X1 new_AGEMA_reg_buffer_3959_s_current_state_reg ( .D(
        new_AGEMA_signal_5846), .CK(clk), .Q(new_AGEMA_signal_5847) );
  DFF_X1 new_AGEMA_reg_buffer_3963_s_current_state_reg ( .D(
        new_AGEMA_signal_5850), .CK(clk), .Q(new_AGEMA_signal_5851) );
  DFF_X1 new_AGEMA_reg_buffer_3967_s_current_state_reg ( .D(
        new_AGEMA_signal_5854), .CK(clk), .Q(new_AGEMA_signal_5855) );
  DFF_X1 new_AGEMA_reg_buffer_3971_s_current_state_reg ( .D(
        new_AGEMA_signal_5858), .CK(clk), .Q(new_AGEMA_signal_5859) );
  DFF_X1 new_AGEMA_reg_buffer_3975_s_current_state_reg ( .D(
        new_AGEMA_signal_5862), .CK(clk), .Q(new_AGEMA_signal_5863) );
  DFF_X1 new_AGEMA_reg_buffer_3979_s_current_state_reg ( .D(
        new_AGEMA_signal_5866), .CK(clk), .Q(new_AGEMA_signal_5867) );
  DFF_X1 new_AGEMA_reg_buffer_3983_s_current_state_reg ( .D(
        new_AGEMA_signal_5870), .CK(clk), .Q(new_AGEMA_signal_5871) );
  DFF_X1 new_AGEMA_reg_buffer_3987_s_current_state_reg ( .D(
        new_AGEMA_signal_5874), .CK(clk), .Q(new_AGEMA_signal_5875) );
  DFF_X1 new_AGEMA_reg_buffer_3991_s_current_state_reg ( .D(
        new_AGEMA_signal_5878), .CK(clk), .Q(new_AGEMA_signal_5879) );
  DFF_X1 new_AGEMA_reg_buffer_3995_s_current_state_reg ( .D(
        new_AGEMA_signal_5882), .CK(clk), .Q(new_AGEMA_signal_5883) );
  DFF_X1 new_AGEMA_reg_buffer_3999_s_current_state_reg ( .D(
        new_AGEMA_signal_5886), .CK(clk), .Q(new_AGEMA_signal_5887) );
  DFF_X1 new_AGEMA_reg_buffer_4003_s_current_state_reg ( .D(
        new_AGEMA_signal_5890), .CK(clk), .Q(new_AGEMA_signal_5891) );
  DFF_X1 new_AGEMA_reg_buffer_4007_s_current_state_reg ( .D(
        new_AGEMA_signal_5894), .CK(clk), .Q(new_AGEMA_signal_5895) );
  DFF_X1 new_AGEMA_reg_buffer_4011_s_current_state_reg ( .D(
        new_AGEMA_signal_5898), .CK(clk), .Q(new_AGEMA_signal_5899) );
  DFF_X1 new_AGEMA_reg_buffer_4015_s_current_state_reg ( .D(
        new_AGEMA_signal_5902), .CK(clk), .Q(new_AGEMA_signal_5903) );
  DFF_X1 new_AGEMA_reg_buffer_4019_s_current_state_reg ( .D(
        new_AGEMA_signal_5906), .CK(clk), .Q(new_AGEMA_signal_5907) );
  DFF_X1 new_AGEMA_reg_buffer_4023_s_current_state_reg ( .D(
        new_AGEMA_signal_5910), .CK(clk), .Q(new_AGEMA_signal_5911) );
  DFF_X1 new_AGEMA_reg_buffer_4027_s_current_state_reg ( .D(
        new_AGEMA_signal_5914), .CK(clk), .Q(new_AGEMA_signal_5915) );
  DFF_X1 new_AGEMA_reg_buffer_4031_s_current_state_reg ( .D(
        new_AGEMA_signal_5918), .CK(clk), .Q(new_AGEMA_signal_5919) );
  DFF_X1 new_AGEMA_reg_buffer_4035_s_current_state_reg ( .D(
        new_AGEMA_signal_5922), .CK(clk), .Q(new_AGEMA_signal_5923) );
  DFF_X1 new_AGEMA_reg_buffer_4039_s_current_state_reg ( .D(
        new_AGEMA_signal_5926), .CK(clk), .Q(new_AGEMA_signal_5927) );
  DFF_X1 new_AGEMA_reg_buffer_4043_s_current_state_reg ( .D(
        new_AGEMA_signal_5930), .CK(clk), .Q(new_AGEMA_signal_5931) );
  DFF_X1 new_AGEMA_reg_buffer_4047_s_current_state_reg ( .D(
        new_AGEMA_signal_5934), .CK(clk), .Q(new_AGEMA_signal_5935) );
  DFF_X1 new_AGEMA_reg_buffer_4051_s_current_state_reg ( .D(
        new_AGEMA_signal_5938), .CK(clk), .Q(new_AGEMA_signal_5939) );
  DFF_X1 new_AGEMA_reg_buffer_4055_s_current_state_reg ( .D(
        new_AGEMA_signal_5942), .CK(clk), .Q(new_AGEMA_signal_5943) );
  DFF_X1 new_AGEMA_reg_buffer_4059_s_current_state_reg ( .D(
        new_AGEMA_signal_5946), .CK(clk), .Q(new_AGEMA_signal_5947) );
  DFF_X1 new_AGEMA_reg_buffer_4063_s_current_state_reg ( .D(
        new_AGEMA_signal_5950), .CK(clk), .Q(new_AGEMA_signal_5951) );
  DFF_X1 new_AGEMA_reg_buffer_4067_s_current_state_reg ( .D(
        new_AGEMA_signal_5954), .CK(clk), .Q(new_AGEMA_signal_5955) );
  DFF_X1 new_AGEMA_reg_buffer_4071_s_current_state_reg ( .D(
        new_AGEMA_signal_5958), .CK(clk), .Q(new_AGEMA_signal_5959) );
  DFF_X1 new_AGEMA_reg_buffer_4075_s_current_state_reg ( .D(
        new_AGEMA_signal_5962), .CK(clk), .Q(new_AGEMA_signal_5963) );
  DFF_X1 new_AGEMA_reg_buffer_4079_s_current_state_reg ( .D(
        new_AGEMA_signal_5966), .CK(clk), .Q(new_AGEMA_signal_5967) );
  DFF_X1 new_AGEMA_reg_buffer_4083_s_current_state_reg ( .D(
        new_AGEMA_signal_5970), .CK(clk), .Q(new_AGEMA_signal_5971) );
  DFF_X1 new_AGEMA_reg_buffer_4087_s_current_state_reg ( .D(
        new_AGEMA_signal_5974), .CK(clk), .Q(new_AGEMA_signal_5975) );
  DFF_X1 new_AGEMA_reg_buffer_4091_s_current_state_reg ( .D(
        new_AGEMA_signal_5978), .CK(clk), .Q(new_AGEMA_signal_5979) );
  DFF_X1 new_AGEMA_reg_buffer_4095_s_current_state_reg ( .D(
        new_AGEMA_signal_5982), .CK(clk), .Q(new_AGEMA_signal_5983) );
  DFF_X1 new_AGEMA_reg_buffer_4099_s_current_state_reg ( .D(
        new_AGEMA_signal_5986), .CK(clk), .Q(new_AGEMA_signal_5987) );
  DFF_X1 new_AGEMA_reg_buffer_4103_s_current_state_reg ( .D(
        new_AGEMA_signal_5990), .CK(clk), .Q(new_AGEMA_signal_5991) );
  DFF_X1 new_AGEMA_reg_buffer_4107_s_current_state_reg ( .D(
        new_AGEMA_signal_5994), .CK(clk), .Q(new_AGEMA_signal_5995) );
  DFF_X1 new_AGEMA_reg_buffer_4111_s_current_state_reg ( .D(
        new_AGEMA_signal_5998), .CK(clk), .Q(new_AGEMA_signal_5999) );
  DFF_X1 new_AGEMA_reg_buffer_4115_s_current_state_reg ( .D(
        new_AGEMA_signal_6002), .CK(clk), .Q(new_AGEMA_signal_6003) );
  DFF_X1 new_AGEMA_reg_buffer_4119_s_current_state_reg ( .D(
        new_AGEMA_signal_6006), .CK(clk), .Q(new_AGEMA_signal_6007) );
  DFF_X1 new_AGEMA_reg_buffer_4123_s_current_state_reg ( .D(
        new_AGEMA_signal_6010), .CK(clk), .Q(new_AGEMA_signal_6011) );
  DFF_X1 new_AGEMA_reg_buffer_4127_s_current_state_reg ( .D(
        new_AGEMA_signal_6014), .CK(clk), .Q(new_AGEMA_signal_6015) );
  DFF_X1 new_AGEMA_reg_buffer_4131_s_current_state_reg ( .D(
        new_AGEMA_signal_6018), .CK(clk), .Q(new_AGEMA_signal_6019) );
  DFF_X1 new_AGEMA_reg_buffer_4135_s_current_state_reg ( .D(
        new_AGEMA_signal_6022), .CK(clk), .Q(new_AGEMA_signal_6023) );
  DFF_X1 new_AGEMA_reg_buffer_4139_s_current_state_reg ( .D(
        new_AGEMA_signal_6026), .CK(clk), .Q(new_AGEMA_signal_6027) );
  DFF_X1 new_AGEMA_reg_buffer_4143_s_current_state_reg ( .D(
        new_AGEMA_signal_6030), .CK(clk), .Q(new_AGEMA_signal_6031) );
  DFF_X1 new_AGEMA_reg_buffer_4147_s_current_state_reg ( .D(
        new_AGEMA_signal_6034), .CK(clk), .Q(new_AGEMA_signal_6035) );
  DFF_X1 new_AGEMA_reg_buffer_4151_s_current_state_reg ( .D(
        new_AGEMA_signal_6038), .CK(clk), .Q(new_AGEMA_signal_6039) );
  DFF_X1 new_AGEMA_reg_buffer_4155_s_current_state_reg ( .D(
        new_AGEMA_signal_6042), .CK(clk), .Q(new_AGEMA_signal_6043) );
  DFF_X1 new_AGEMA_reg_buffer_4159_s_current_state_reg ( .D(
        new_AGEMA_signal_6046), .CK(clk), .Q(new_AGEMA_signal_6047) );
  DFF_X1 new_AGEMA_reg_buffer_4163_s_current_state_reg ( .D(
        new_AGEMA_signal_6050), .CK(clk), .Q(new_AGEMA_signal_6051) );
  DFF_X1 new_AGEMA_reg_buffer_4167_s_current_state_reg ( .D(
        new_AGEMA_signal_6054), .CK(clk), .Q(new_AGEMA_signal_6055) );
  DFF_X1 new_AGEMA_reg_buffer_4171_s_current_state_reg ( .D(
        new_AGEMA_signal_6058), .CK(clk), .Q(new_AGEMA_signal_6059) );
  DFF_X1 new_AGEMA_reg_buffer_4175_s_current_state_reg ( .D(
        new_AGEMA_signal_6062), .CK(clk), .Q(new_AGEMA_signal_6063) );
  DFF_X1 new_AGEMA_reg_buffer_4179_s_current_state_reg ( .D(
        new_AGEMA_signal_6066), .CK(clk), .Q(new_AGEMA_signal_6067) );
  DFF_X1 new_AGEMA_reg_buffer_4183_s_current_state_reg ( .D(
        new_AGEMA_signal_6070), .CK(clk), .Q(new_AGEMA_signal_6071) );
  DFF_X1 new_AGEMA_reg_buffer_4187_s_current_state_reg ( .D(
        new_AGEMA_signal_6074), .CK(clk), .Q(new_AGEMA_signal_6075) );
  DFF_X1 new_AGEMA_reg_buffer_4191_s_current_state_reg ( .D(
        new_AGEMA_signal_6078), .CK(clk), .Q(new_AGEMA_signal_6079) );
  DFF_X1 new_AGEMA_reg_buffer_4195_s_current_state_reg ( .D(
        new_AGEMA_signal_6082), .CK(clk), .Q(new_AGEMA_signal_6083) );
  DFF_X1 new_AGEMA_reg_buffer_4199_s_current_state_reg ( .D(
        new_AGEMA_signal_6086), .CK(clk), .Q(new_AGEMA_signal_6087) );
  DFF_X1 new_AGEMA_reg_buffer_4203_s_current_state_reg ( .D(
        new_AGEMA_signal_6090), .CK(clk), .Q(new_AGEMA_signal_6091) );
  DFF_X1 new_AGEMA_reg_buffer_4207_s_current_state_reg ( .D(
        new_AGEMA_signal_6094), .CK(clk), .Q(new_AGEMA_signal_6095) );
  DFF_X1 new_AGEMA_reg_buffer_4211_s_current_state_reg ( .D(
        new_AGEMA_signal_6098), .CK(clk), .Q(new_AGEMA_signal_6099) );
  DFF_X1 new_AGEMA_reg_buffer_4215_s_current_state_reg ( .D(
        new_AGEMA_signal_6102), .CK(clk), .Q(new_AGEMA_signal_6103) );
  DFF_X1 new_AGEMA_reg_buffer_4219_s_current_state_reg ( .D(
        new_AGEMA_signal_6106), .CK(clk), .Q(new_AGEMA_signal_6107) );
  DFF_X1 new_AGEMA_reg_buffer_4223_s_current_state_reg ( .D(
        new_AGEMA_signal_6110), .CK(clk), .Q(new_AGEMA_signal_6111) );
  DFF_X1 new_AGEMA_reg_buffer_4227_s_current_state_reg ( .D(
        new_AGEMA_signal_6114), .CK(clk), .Q(new_AGEMA_signal_6115) );
  DFF_X1 new_AGEMA_reg_buffer_4231_s_current_state_reg ( .D(
        new_AGEMA_signal_6118), .CK(clk), .Q(new_AGEMA_signal_6119) );
  DFF_X1 new_AGEMA_reg_buffer_4235_s_current_state_reg ( .D(
        new_AGEMA_signal_6122), .CK(clk), .Q(new_AGEMA_signal_6123) );
  DFF_X1 new_AGEMA_reg_buffer_4239_s_current_state_reg ( .D(
        new_AGEMA_signal_6126), .CK(clk), .Q(new_AGEMA_signal_6127) );
  DFF_X1 new_AGEMA_reg_buffer_4243_s_current_state_reg ( .D(
        new_AGEMA_signal_6130), .CK(clk), .Q(new_AGEMA_signal_6131) );
  DFF_X1 new_AGEMA_reg_buffer_4247_s_current_state_reg ( .D(
        new_AGEMA_signal_6134), .CK(clk), .Q(new_AGEMA_signal_6135) );
  DFF_X1 new_AGEMA_reg_buffer_4251_s_current_state_reg ( .D(
        new_AGEMA_signal_6138), .CK(clk), .Q(new_AGEMA_signal_6139) );
  DFF_X1 new_AGEMA_reg_buffer_4255_s_current_state_reg ( .D(
        new_AGEMA_signal_6142), .CK(clk), .Q(new_AGEMA_signal_6143) );
  DFF_X1 new_AGEMA_reg_buffer_4259_s_current_state_reg ( .D(
        new_AGEMA_signal_6146), .CK(clk), .Q(new_AGEMA_signal_6147) );
  DFF_X1 new_AGEMA_reg_buffer_4263_s_current_state_reg ( .D(
        new_AGEMA_signal_6150), .CK(clk), .Q(new_AGEMA_signal_6151) );
  DFF_X1 new_AGEMA_reg_buffer_4267_s_current_state_reg ( .D(
        new_AGEMA_signal_6154), .CK(clk), .Q(new_AGEMA_signal_6155) );
  DFF_X1 new_AGEMA_reg_buffer_4271_s_current_state_reg ( .D(
        new_AGEMA_signal_6158), .CK(clk), .Q(new_AGEMA_signal_6159) );
  DFF_X1 new_AGEMA_reg_buffer_4275_s_current_state_reg ( .D(
        new_AGEMA_signal_6162), .CK(clk), .Q(new_AGEMA_signal_6163) );
  DFF_X1 new_AGEMA_reg_buffer_4279_s_current_state_reg ( .D(
        new_AGEMA_signal_6166), .CK(clk), .Q(new_AGEMA_signal_6167) );
  DFF_X1 new_AGEMA_reg_buffer_4283_s_current_state_reg ( .D(
        new_AGEMA_signal_6170), .CK(clk), .Q(new_AGEMA_signal_6171) );
  DFF_X1 new_AGEMA_reg_buffer_4287_s_current_state_reg ( .D(
        new_AGEMA_signal_6174), .CK(clk), .Q(new_AGEMA_signal_6175) );
  DFF_X1 new_AGEMA_reg_buffer_4291_s_current_state_reg ( .D(
        new_AGEMA_signal_6178), .CK(clk), .Q(new_AGEMA_signal_6179) );
  DFF_X1 new_AGEMA_reg_buffer_4295_s_current_state_reg ( .D(
        new_AGEMA_signal_6182), .CK(clk), .Q(new_AGEMA_signal_6183) );
  DFF_X1 new_AGEMA_reg_buffer_4299_s_current_state_reg ( .D(
        new_AGEMA_signal_6186), .CK(clk), .Q(new_AGEMA_signal_6187) );
  DFF_X1 new_AGEMA_reg_buffer_4303_s_current_state_reg ( .D(
        new_AGEMA_signal_6190), .CK(clk), .Q(new_AGEMA_signal_6191) );
  DFF_X1 new_AGEMA_reg_buffer_4307_s_current_state_reg ( .D(
        new_AGEMA_signal_6194), .CK(clk), .Q(new_AGEMA_signal_6195) );
  DFF_X1 new_AGEMA_reg_buffer_4311_s_current_state_reg ( .D(
        new_AGEMA_signal_6198), .CK(clk), .Q(new_AGEMA_signal_6199) );
  DFF_X1 new_AGEMA_reg_buffer_4315_s_current_state_reg ( .D(
        new_AGEMA_signal_6202), .CK(clk), .Q(new_AGEMA_signal_6203) );
  DFF_X1 new_AGEMA_reg_buffer_4319_s_current_state_reg ( .D(
        new_AGEMA_signal_6206), .CK(clk), .Q(new_AGEMA_signal_6207) );
  DFF_X1 new_AGEMA_reg_buffer_4323_s_current_state_reg ( .D(
        new_AGEMA_signal_6210), .CK(clk), .Q(new_AGEMA_signal_6211) );
  DFF_X1 new_AGEMA_reg_buffer_4327_s_current_state_reg ( .D(
        new_AGEMA_signal_6214), .CK(clk), .Q(new_AGEMA_signal_6215) );
  DFF_X1 new_AGEMA_reg_buffer_4331_s_current_state_reg ( .D(
        new_AGEMA_signal_6218), .CK(clk), .Q(new_AGEMA_signal_6219) );
  DFF_X1 new_AGEMA_reg_buffer_4335_s_current_state_reg ( .D(
        new_AGEMA_signal_6222), .CK(clk), .Q(new_AGEMA_signal_6223) );
  DFF_X1 new_AGEMA_reg_buffer_4339_s_current_state_reg ( .D(
        new_AGEMA_signal_6226), .CK(clk), .Q(new_AGEMA_signal_6227) );
  AND2_X1 Inst_bSbox_AND_M29_U1_U16 ( .A1(new_AGEMA_signal_3389), .A2(
        new_AGEMA_signal_3615), .ZN(Inst_bSbox_AND_M29_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M29_U1_U15 ( .A1(Inst_bSbox_M28), .A2(
        new_AGEMA_signal_3614), .ZN(Inst_bSbox_AND_M29_U1_mul[0]) );
  XOR2_X1 Inst_bSbox_AND_M29_U1_U14 ( .A(Fresh[24]), .B(
        Inst_bSbox_AND_M29_U1_n23), .Z(Inst_bSbox_AND_M29_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M29_U1_U13 ( .A1(new_AGEMA_signal_3389), .A2(
        Inst_bSbox_AND_M29_U1_n22), .ZN(Inst_bSbox_AND_M29_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M29_U1_U12 ( .A(Fresh[24]), .B(
        Inst_bSbox_AND_M29_U1_n21), .Z(Inst_bSbox_AND_M29_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M29_U1_U11 ( .A1(Inst_bSbox_M28), .A2(
        Inst_bSbox_AND_M29_U1_n22), .ZN(Inst_bSbox_AND_M29_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M29_U1_U10 ( .A(Inst_bSbox_AND_M29_U1_n20), .B(
        Inst_bSbox_AND_M29_U1_n19), .ZN(Inst_bSbox_M29) );
  NAND2_X1 Inst_bSbox_AND_M29_U1_U9 ( .A1(Inst_bSbox_AND_M29_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M29_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M29_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M29_U1_U8 ( .A(Inst_bSbox_AND_M29_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M29_U1_z[0]), .Z(Inst_bSbox_AND_M29_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M29_U1_U7 ( .A(Inst_bSbox_AND_M29_U1_n18), .B(
        Inst_bSbox_AND_M29_U1_n17), .ZN(new_AGEMA_signal_3392) );
  NAND2_X1 Inst_bSbox_AND_M29_U1_U6 ( .A1(Inst_bSbox_AND_M29_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M29_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M29_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M29_U1_U5 ( .A(Inst_bSbox_AND_M29_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M29_U1_z[1]), .Z(Inst_bSbox_AND_M29_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M29_U1_U4 ( .A(new_AGEMA_signal_3615), .B(
        Inst_bSbox_AND_M29_U1_n22), .ZN(Inst_bSbox_AND_M29_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M29_U1_U3 ( .A(new_AGEMA_signal_3614), .B(
        Inst_bSbox_AND_M29_U1_n22), .ZN(Inst_bSbox_AND_M29_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M29_U1_U2 ( .A(Fresh[25]), .ZN(
        Inst_bSbox_AND_M29_U1_n22) );
  DFF_X1 Inst_bSbox_AND_M29_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M29_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M29_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M28),
        .CK(clk), .Q(Inst_bSbox_AND_M29_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M29_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M29_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M29_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M29_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M29_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M29_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M29_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3389), .CK(clk), .Q(Inst_bSbox_AND_M29_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M29_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M29_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M29_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M29_U1_p_0_out_1__0_) );
  AND2_X1 Inst_bSbox_AND_M30_U1_U16 ( .A1(new_AGEMA_signal_3388), .A2(
        new_AGEMA_signal_3617), .ZN(Inst_bSbox_AND_M30_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M30_U1_U15 ( .A1(Inst_bSbox_M26), .A2(
        new_AGEMA_signal_3616), .ZN(Inst_bSbox_AND_M30_U1_mul[0]) );
  XOR2_X1 Inst_bSbox_AND_M30_U1_U14 ( .A(Fresh[26]), .B(
        Inst_bSbox_AND_M30_U1_n23), .Z(Inst_bSbox_AND_M30_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M30_U1_U13 ( .A1(new_AGEMA_signal_3388), .A2(
        Inst_bSbox_AND_M30_U1_n22), .ZN(Inst_bSbox_AND_M30_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M30_U1_U12 ( .A(Fresh[26]), .B(
        Inst_bSbox_AND_M30_U1_n21), .Z(Inst_bSbox_AND_M30_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M30_U1_U11 ( .A1(Inst_bSbox_M26), .A2(
        Inst_bSbox_AND_M30_U1_n22), .ZN(Inst_bSbox_AND_M30_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M30_U1_U10 ( .A(Inst_bSbox_AND_M30_U1_n20), .B(
        Inst_bSbox_AND_M30_U1_n19), .ZN(Inst_bSbox_M30) );
  NAND2_X1 Inst_bSbox_AND_M30_U1_U9 ( .A1(Inst_bSbox_AND_M30_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M30_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M30_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M30_U1_U8 ( .A(Inst_bSbox_AND_M30_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M30_U1_z[0]), .Z(Inst_bSbox_AND_M30_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M30_U1_U7 ( .A(Inst_bSbox_AND_M30_U1_n18), .B(
        Inst_bSbox_AND_M30_U1_n17), .ZN(new_AGEMA_signal_3393) );
  NAND2_X1 Inst_bSbox_AND_M30_U1_U6 ( .A1(Inst_bSbox_AND_M30_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M30_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M30_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M30_U1_U5 ( .A(Inst_bSbox_AND_M30_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M30_U1_z[1]), .Z(Inst_bSbox_AND_M30_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M30_U1_U4 ( .A(new_AGEMA_signal_3617), .B(
        Inst_bSbox_AND_M30_U1_n22), .ZN(Inst_bSbox_AND_M30_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M30_U1_U3 ( .A(new_AGEMA_signal_3616), .B(
        Inst_bSbox_AND_M30_U1_n22), .ZN(Inst_bSbox_AND_M30_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M30_U1_U2 ( .A(Fresh[27]), .ZN(
        Inst_bSbox_AND_M30_U1_n22) );
  DFF_X1 Inst_bSbox_AND_M30_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M30_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M30_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M26),
        .CK(clk), .Q(Inst_bSbox_AND_M30_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M30_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M30_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M30_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M30_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M30_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M30_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M30_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3388), .CK(clk), .Q(Inst_bSbox_AND_M30_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M30_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M30_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M30_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M30_U1_p_0_out_1__0_) );
  AND2_X1 Inst_bSbox_AND_M32_U1_U16 ( .A1(new_AGEMA_signal_3615), .A2(
        new_AGEMA_signal_3390), .ZN(Inst_bSbox_AND_M32_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M32_U1_U15 ( .A1(new_AGEMA_signal_3614), .A2(
        Inst_bSbox_M31), .ZN(Inst_bSbox_AND_M32_U1_mul[0]) );
  XOR2_X1 Inst_bSbox_AND_M32_U1_U14 ( .A(Fresh[28]), .B(
        Inst_bSbox_AND_M32_U1_n23), .Z(Inst_bSbox_AND_M32_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M32_U1_U13 ( .A1(new_AGEMA_signal_3615), .A2(
        Inst_bSbox_AND_M32_U1_n22), .ZN(Inst_bSbox_AND_M32_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M32_U1_U12 ( .A(Fresh[28]), .B(
        Inst_bSbox_AND_M32_U1_n21), .Z(Inst_bSbox_AND_M32_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M32_U1_U11 ( .A1(new_AGEMA_signal_3614), .A2(
        Inst_bSbox_AND_M32_U1_n22), .ZN(Inst_bSbox_AND_M32_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M32_U1_U10 ( .A(Inst_bSbox_AND_M32_U1_n20), .B(
        Inst_bSbox_AND_M32_U1_n19), .ZN(Inst_bSbox_M32) );
  NAND2_X1 Inst_bSbox_AND_M32_U1_U9 ( .A1(Inst_bSbox_AND_M32_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M32_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M32_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M32_U1_U8 ( .A(Inst_bSbox_AND_M32_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M32_U1_z[0]), .Z(Inst_bSbox_AND_M32_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M32_U1_U7 ( .A(Inst_bSbox_AND_M32_U1_n18), .B(
        Inst_bSbox_AND_M32_U1_n17), .ZN(new_AGEMA_signal_3394) );
  NAND2_X1 Inst_bSbox_AND_M32_U1_U6 ( .A1(Inst_bSbox_AND_M32_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M32_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M32_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M32_U1_U5 ( .A(Inst_bSbox_AND_M32_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M32_U1_z[1]), .Z(Inst_bSbox_AND_M32_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M32_U1_U4 ( .A(new_AGEMA_signal_3390), .B(
        Inst_bSbox_AND_M32_U1_n22), .ZN(Inst_bSbox_AND_M32_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M32_U1_U3 ( .A(Inst_bSbox_M31), .B(
        Inst_bSbox_AND_M32_U1_n22), .ZN(Inst_bSbox_AND_M32_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M32_U1_U2 ( .A(Fresh[29]), .ZN(
        Inst_bSbox_AND_M32_U1_n22) );
  DFF_X1 Inst_bSbox_AND_M32_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M32_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M32_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3614), .CK(clk), .Q(Inst_bSbox_AND_M32_U1_a_reg[0])
         );
  DFF_X1 Inst_bSbox_AND_M32_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M32_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M32_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M32_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M32_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M32_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M32_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3615), .CK(clk), .Q(Inst_bSbox_AND_M32_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M32_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M32_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M32_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M32_U1_p_0_out_1__0_) );
  AND2_X1 Inst_bSbox_AND_M35_U1_U16 ( .A1(new_AGEMA_signal_3617), .A2(
        new_AGEMA_signal_3386), .ZN(Inst_bSbox_AND_M35_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M35_U1_U15 ( .A1(new_AGEMA_signal_3616), .A2(
        Inst_bSbox_M34), .ZN(Inst_bSbox_AND_M35_U1_mul[0]) );
  XOR2_X1 Inst_bSbox_AND_M35_U1_U14 ( .A(Fresh[30]), .B(
        Inst_bSbox_AND_M35_U1_n23), .Z(Inst_bSbox_AND_M35_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M35_U1_U13 ( .A1(new_AGEMA_signal_3617), .A2(
        Inst_bSbox_AND_M35_U1_n22), .ZN(Inst_bSbox_AND_M35_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M35_U1_U12 ( .A(Fresh[30]), .B(
        Inst_bSbox_AND_M35_U1_n21), .Z(Inst_bSbox_AND_M35_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M35_U1_U11 ( .A1(new_AGEMA_signal_3616), .A2(
        Inst_bSbox_AND_M35_U1_n22), .ZN(Inst_bSbox_AND_M35_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M35_U1_U10 ( .A(Inst_bSbox_AND_M35_U1_n20), .B(
        Inst_bSbox_AND_M35_U1_n19), .ZN(Inst_bSbox_M35) );
  NAND2_X1 Inst_bSbox_AND_M35_U1_U9 ( .A1(Inst_bSbox_AND_M35_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M35_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M35_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M35_U1_U8 ( .A(Inst_bSbox_AND_M35_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M35_U1_z[0]), .Z(Inst_bSbox_AND_M35_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M35_U1_U7 ( .A(Inst_bSbox_AND_M35_U1_n18), .B(
        Inst_bSbox_AND_M35_U1_n17), .ZN(new_AGEMA_signal_3395) );
  NAND2_X1 Inst_bSbox_AND_M35_U1_U6 ( .A1(Inst_bSbox_AND_M35_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M35_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M35_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M35_U1_U5 ( .A(Inst_bSbox_AND_M35_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M35_U1_z[1]), .Z(Inst_bSbox_AND_M35_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M35_U1_U4 ( .A(new_AGEMA_signal_3386), .B(
        Inst_bSbox_AND_M35_U1_n22), .ZN(Inst_bSbox_AND_M35_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M35_U1_U3 ( .A(Inst_bSbox_M34), .B(
        Inst_bSbox_AND_M35_U1_n22), .ZN(Inst_bSbox_AND_M35_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M35_U1_U2 ( .A(Fresh[31]), .ZN(
        Inst_bSbox_AND_M35_U1_n22) );
  DFF_X1 Inst_bSbox_AND_M35_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M35_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M35_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3616), .CK(clk), .Q(Inst_bSbox_AND_M35_U1_a_reg[0])
         );
  DFF_X1 Inst_bSbox_AND_M35_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M35_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M35_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M35_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M35_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M35_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M35_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3617), .CK(clk), .Q(Inst_bSbox_AND_M35_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M35_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M35_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M35_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M35_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_M37_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3618), .B(
        Inst_bSbox_M29), .Z(Inst_bSbox_M37) );
  XOR2_X1 Inst_bSbox_XOR_M37_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3619), .B(
        new_AGEMA_signal_3392), .Z(new_AGEMA_signal_3397) );
  XOR2_X1 Inst_bSbox_XOR_M38_U1_Ins_0_U1 ( .A(Inst_bSbox_M32), .B(
        new_AGEMA_signal_3620), .Z(Inst_bSbox_M38) );
  XOR2_X1 Inst_bSbox_XOR_M38_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3394), .B(
        new_AGEMA_signal_3621), .Z(new_AGEMA_signal_3398) );
  XOR2_X1 Inst_bSbox_XOR_M39_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3622), .B(
        Inst_bSbox_M30), .Z(Inst_bSbox_M39) );
  XOR2_X1 Inst_bSbox_XOR_M39_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3623), .B(
        new_AGEMA_signal_3393), .Z(new_AGEMA_signal_3399) );
  XOR2_X1 Inst_bSbox_XOR_M40_U1_Ins_0_U1 ( .A(Inst_bSbox_M35), .B(
        new_AGEMA_signal_3624), .Z(Inst_bSbox_M40) );
  XOR2_X1 Inst_bSbox_XOR_M40_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3395), .B(
        new_AGEMA_signal_3625), .Z(new_AGEMA_signal_3400) );
  XOR2_X1 Inst_bSbox_XOR_M41_U1_Ins_0_U1 ( .A(Inst_bSbox_M38), .B(
        Inst_bSbox_M40), .Z(Inst_bSbox_M41) );
  XOR2_X1 Inst_bSbox_XOR_M41_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3398), .B(
        new_AGEMA_signal_3400), .Z(new_AGEMA_signal_3401) );
  XOR2_X1 Inst_bSbox_XOR_M42_U1_Ins_0_U1 ( .A(Inst_bSbox_M37), .B(
        Inst_bSbox_M39), .Z(Inst_bSbox_M42) );
  XOR2_X1 Inst_bSbox_XOR_M42_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3397), .B(
        new_AGEMA_signal_3399), .Z(new_AGEMA_signal_3402) );
  XOR2_X1 Inst_bSbox_XOR_M43_U1_Ins_0_U1 ( .A(Inst_bSbox_M37), .B(
        Inst_bSbox_M38), .Z(Inst_bSbox_M43) );
  XOR2_X1 Inst_bSbox_XOR_M43_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3397), .B(
        new_AGEMA_signal_3398), .Z(new_AGEMA_signal_3403) );
  XOR2_X1 Inst_bSbox_XOR_M44_U1_Ins_0_U1 ( .A(Inst_bSbox_M39), .B(
        Inst_bSbox_M40), .Z(Inst_bSbox_M44) );
  XOR2_X1 Inst_bSbox_XOR_M44_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3399), .B(
        new_AGEMA_signal_3400), .Z(new_AGEMA_signal_3404) );
  XOR2_X1 Inst_bSbox_XOR_M45_U1_Ins_0_U1 ( .A(Inst_bSbox_M42), .B(
        Inst_bSbox_M41), .Z(Inst_bSbox_M45) );
  XOR2_X1 Inst_bSbox_XOR_M45_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3402), .B(
        new_AGEMA_signal_3401), .Z(new_AGEMA_signal_3413) );
  DFF_X1 new_AGEMA_reg_buffer_1730_s_current_state_reg ( .D(
        new_AGEMA_signal_3610), .CK(clk), .Q(new_AGEMA_signal_3618) );
  DFF_X1 new_AGEMA_reg_buffer_1731_s_current_state_reg ( .D(
        new_AGEMA_signal_3611), .CK(clk), .Q(new_AGEMA_signal_3619) );
  DFF_X1 new_AGEMA_reg_buffer_1732_s_current_state_reg ( .D(Inst_bSbox_M33),
        .CK(clk), .Q(new_AGEMA_signal_3620) );
  DFF_X1 new_AGEMA_reg_buffer_1733_s_current_state_reg ( .D(
        new_AGEMA_signal_3391), .CK(clk), .Q(new_AGEMA_signal_3621) );
  DFF_X1 new_AGEMA_reg_buffer_1734_s_current_state_reg ( .D(
        new_AGEMA_signal_3612), .CK(clk), .Q(new_AGEMA_signal_3622) );
  DFF_X1 new_AGEMA_reg_buffer_1735_s_current_state_reg ( .D(
        new_AGEMA_signal_3613), .CK(clk), .Q(new_AGEMA_signal_3623) );
  DFF_X1 new_AGEMA_reg_buffer_1736_s_current_state_reg ( .D(Inst_bSbox_M36),
        .CK(clk), .Q(new_AGEMA_signal_3624) );
  DFF_X1 new_AGEMA_reg_buffer_1737_s_current_state_reg ( .D(
        new_AGEMA_signal_3396), .CK(clk), .Q(new_AGEMA_signal_3625) );
  DFF_X1 new_AGEMA_reg_buffer_1740_s_current_state_reg ( .D(
        new_AGEMA_signal_3627), .CK(clk), .Q(new_AGEMA_signal_3628) );
  DFF_X1 new_AGEMA_reg_buffer_1744_s_current_state_reg ( .D(
        new_AGEMA_signal_3631), .CK(clk), .Q(new_AGEMA_signal_3632) );
  DFF_X1 new_AGEMA_reg_buffer_1748_s_current_state_reg ( .D(
        new_AGEMA_signal_3635), .CK(clk), .Q(new_AGEMA_signal_3636) );
  DFF_X1 new_AGEMA_reg_buffer_1752_s_current_state_reg ( .D(
        new_AGEMA_signal_3639), .CK(clk), .Q(new_AGEMA_signal_3640) );
  DFF_X1 new_AGEMA_reg_buffer_1756_s_current_state_reg ( .D(
        new_AGEMA_signal_3643), .CK(clk), .Q(new_AGEMA_signal_3644) );
  DFF_X1 new_AGEMA_reg_buffer_1760_s_current_state_reg ( .D(
        new_AGEMA_signal_3647), .CK(clk), .Q(new_AGEMA_signal_3648) );
  DFF_X1 new_AGEMA_reg_buffer_1764_s_current_state_reg ( .D(
        new_AGEMA_signal_3651), .CK(clk), .Q(new_AGEMA_signal_3652) );
  DFF_X1 new_AGEMA_reg_buffer_1768_s_current_state_reg ( .D(
        new_AGEMA_signal_3655), .CK(clk), .Q(new_AGEMA_signal_3656) );
  DFF_X1 new_AGEMA_reg_buffer_1772_s_current_state_reg ( .D(
        new_AGEMA_signal_3659), .CK(clk), .Q(new_AGEMA_signal_3660) );
  DFF_X1 new_AGEMA_reg_buffer_1776_s_current_state_reg ( .D(
        new_AGEMA_signal_3663), .CK(clk), .Q(new_AGEMA_signal_3664) );
  DFF_X1 new_AGEMA_reg_buffer_1780_s_current_state_reg ( .D(
        new_AGEMA_signal_3667), .CK(clk), .Q(new_AGEMA_signal_3668) );
  DFF_X1 new_AGEMA_reg_buffer_1784_s_current_state_reg ( .D(
        new_AGEMA_signal_3671), .CK(clk), .Q(new_AGEMA_signal_3672) );
  DFF_X1 new_AGEMA_reg_buffer_1788_s_current_state_reg ( .D(
        new_AGEMA_signal_3675), .CK(clk), .Q(new_AGEMA_signal_3676) );
  DFF_X1 new_AGEMA_reg_buffer_1792_s_current_state_reg ( .D(
        new_AGEMA_signal_3679), .CK(clk), .Q(new_AGEMA_signal_3680) );
  DFF_X1 new_AGEMA_reg_buffer_1796_s_current_state_reg ( .D(
        new_AGEMA_signal_3683), .CK(clk), .Q(new_AGEMA_signal_3684) );
  DFF_X1 new_AGEMA_reg_buffer_1800_s_current_state_reg ( .D(
        new_AGEMA_signal_3687), .CK(clk), .Q(new_AGEMA_signal_3688) );
  DFF_X1 new_AGEMA_reg_buffer_1804_s_current_state_reg ( .D(
        new_AGEMA_signal_3691), .CK(clk), .Q(new_AGEMA_signal_3692) );
  DFF_X1 new_AGEMA_reg_buffer_1808_s_current_state_reg ( .D(
        new_AGEMA_signal_3695), .CK(clk), .Q(new_AGEMA_signal_3696) );
  DFF_X1 new_AGEMA_reg_buffer_1812_s_current_state_reg ( .D(
        new_AGEMA_signal_3699), .CK(clk), .Q(new_AGEMA_signal_3700) );
  DFF_X1 new_AGEMA_reg_buffer_1816_s_current_state_reg ( .D(
        new_AGEMA_signal_3703), .CK(clk), .Q(new_AGEMA_signal_3704) );
  DFF_X1 new_AGEMA_reg_buffer_1820_s_current_state_reg ( .D(
        new_AGEMA_signal_3707), .CK(clk), .Q(new_AGEMA_signal_3708) );
  DFF_X1 new_AGEMA_reg_buffer_1824_s_current_state_reg ( .D(
        new_AGEMA_signal_3711), .CK(clk), .Q(new_AGEMA_signal_3712) );
  DFF_X1 new_AGEMA_reg_buffer_1828_s_current_state_reg ( .D(
        new_AGEMA_signal_3715), .CK(clk), .Q(new_AGEMA_signal_3716) );
  DFF_X1 new_AGEMA_reg_buffer_1832_s_current_state_reg ( .D(
        new_AGEMA_signal_3719), .CK(clk), .Q(new_AGEMA_signal_3720) );
  DFF_X1 new_AGEMA_reg_buffer_1836_s_current_state_reg ( .D(
        new_AGEMA_signal_3723), .CK(clk), .Q(new_AGEMA_signal_3724) );
  DFF_X1 new_AGEMA_reg_buffer_1840_s_current_state_reg ( .D(
        new_AGEMA_signal_3727), .CK(clk), .Q(new_AGEMA_signal_3728) );
  DFF_X1 new_AGEMA_reg_buffer_1844_s_current_state_reg ( .D(
        new_AGEMA_signal_3731), .CK(clk), .Q(new_AGEMA_signal_3732) );
  DFF_X1 new_AGEMA_reg_buffer_1848_s_current_state_reg ( .D(
        new_AGEMA_signal_3735), .CK(clk), .Q(new_AGEMA_signal_3736) );
  DFF_X1 new_AGEMA_reg_buffer_1852_s_current_state_reg ( .D(
        new_AGEMA_signal_3739), .CK(clk), .Q(new_AGEMA_signal_3740) );
  DFF_X1 new_AGEMA_reg_buffer_1856_s_current_state_reg ( .D(
        new_AGEMA_signal_3743), .CK(clk), .Q(new_AGEMA_signal_3744) );
  DFF_X1 new_AGEMA_reg_buffer_1860_s_current_state_reg ( .D(
        new_AGEMA_signal_3747), .CK(clk), .Q(new_AGEMA_signal_3748) );
  DFF_X1 new_AGEMA_reg_buffer_1864_s_current_state_reg ( .D(
        new_AGEMA_signal_3751), .CK(clk), .Q(new_AGEMA_signal_3752) );
  DFF_X1 new_AGEMA_reg_buffer_1868_s_current_state_reg ( .D(
        new_AGEMA_signal_3755), .CK(clk), .Q(new_AGEMA_signal_3756) );
  DFF_X1 new_AGEMA_reg_buffer_1872_s_current_state_reg ( .D(
        new_AGEMA_signal_3759), .CK(clk), .Q(new_AGEMA_signal_3760) );
  DFF_X1 new_AGEMA_reg_buffer_1876_s_current_state_reg ( .D(
        new_AGEMA_signal_3763), .CK(clk), .Q(new_AGEMA_signal_3764) );
  DFF_X1 new_AGEMA_reg_buffer_1880_s_current_state_reg ( .D(
        new_AGEMA_signal_3767), .CK(clk), .Q(new_AGEMA_signal_3768) );
  DFF_X1 new_AGEMA_reg_buffer_1884_s_current_state_reg ( .D(
        new_AGEMA_signal_3771), .CK(clk), .Q(new_AGEMA_signal_3772) );
  DFF_X1 new_AGEMA_reg_buffer_1888_s_current_state_reg ( .D(
        new_AGEMA_signal_3775), .CK(clk), .Q(new_AGEMA_signal_3776) );
  DFF_X1 new_AGEMA_reg_buffer_1892_s_current_state_reg ( .D(
        new_AGEMA_signal_3779), .CK(clk), .Q(new_AGEMA_signal_3780) );
  DFF_X1 new_AGEMA_reg_buffer_1896_s_current_state_reg ( .D(
        new_AGEMA_signal_3783), .CK(clk), .Q(new_AGEMA_signal_3784) );
  DFF_X1 new_AGEMA_reg_buffer_1900_s_current_state_reg ( .D(
        new_AGEMA_signal_3787), .CK(clk), .Q(new_AGEMA_signal_3788) );
  DFF_X1 new_AGEMA_reg_buffer_1904_s_current_state_reg ( .D(
        new_AGEMA_signal_3791), .CK(clk), .Q(new_AGEMA_signal_3792) );
  DFF_X1 new_AGEMA_reg_buffer_1908_s_current_state_reg ( .D(
        new_AGEMA_signal_3795), .CK(clk), .Q(new_AGEMA_signal_3796) );
  DFF_X1 new_AGEMA_reg_buffer_1912_s_current_state_reg ( .D(
        new_AGEMA_signal_3799), .CK(clk), .Q(new_AGEMA_signal_3800) );
  DFF_X1 new_AGEMA_reg_buffer_1916_s_current_state_reg ( .D(
        new_AGEMA_signal_3803), .CK(clk), .Q(new_AGEMA_signal_3804) );
  DFF_X1 new_AGEMA_reg_buffer_1920_s_current_state_reg ( .D(
        new_AGEMA_signal_3807), .CK(clk), .Q(new_AGEMA_signal_3808) );
  DFF_X1 new_AGEMA_reg_buffer_1924_s_current_state_reg ( .D(
        new_AGEMA_signal_3811), .CK(clk), .Q(new_AGEMA_signal_3812) );
  DFF_X1 new_AGEMA_reg_buffer_1928_s_current_state_reg ( .D(
        new_AGEMA_signal_3815), .CK(clk), .Q(new_AGEMA_signal_3816) );
  DFF_X1 new_AGEMA_reg_buffer_1932_s_current_state_reg ( .D(
        new_AGEMA_signal_3819), .CK(clk), .Q(new_AGEMA_signal_3820) );
  DFF_X1 new_AGEMA_reg_buffer_1936_s_current_state_reg ( .D(
        new_AGEMA_signal_3823), .CK(clk), .Q(new_AGEMA_signal_3824) );
  DFF_X1 new_AGEMA_reg_buffer_1940_s_current_state_reg ( .D(
        new_AGEMA_signal_3827), .CK(clk), .Q(new_AGEMA_signal_3828) );
  DFF_X1 new_AGEMA_reg_buffer_1944_s_current_state_reg ( .D(
        new_AGEMA_signal_3831), .CK(clk), .Q(new_AGEMA_signal_3832) );
  DFF_X1 new_AGEMA_reg_buffer_1948_s_current_state_reg ( .D(
        new_AGEMA_signal_3835), .CK(clk), .Q(new_AGEMA_signal_3836) );
  DFF_X1 new_AGEMA_reg_buffer_1952_s_current_state_reg ( .D(
        new_AGEMA_signal_3839), .CK(clk), .Q(new_AGEMA_signal_3840) );
  DFF_X1 new_AGEMA_reg_buffer_1956_s_current_state_reg ( .D(
        new_AGEMA_signal_3843), .CK(clk), .Q(new_AGEMA_signal_3844) );
  DFF_X1 new_AGEMA_reg_buffer_1960_s_current_state_reg ( .D(
        new_AGEMA_signal_3847), .CK(clk), .Q(new_AGEMA_signal_3848) );
  DFF_X1 new_AGEMA_reg_buffer_1964_s_current_state_reg ( .D(
        new_AGEMA_signal_3851), .CK(clk), .Q(new_AGEMA_signal_3852) );
  DFF_X1 new_AGEMA_reg_buffer_1968_s_current_state_reg ( .D(
        new_AGEMA_signal_3855), .CK(clk), .Q(new_AGEMA_signal_3856) );
  DFF_X1 new_AGEMA_reg_buffer_1972_s_current_state_reg ( .D(
        new_AGEMA_signal_3859), .CK(clk), .Q(new_AGEMA_signal_3860) );
  DFF_X1 new_AGEMA_reg_buffer_1976_s_current_state_reg ( .D(
        new_AGEMA_signal_3863), .CK(clk), .Q(new_AGEMA_signal_3864) );
  DFF_X1 new_AGEMA_reg_buffer_1980_s_current_state_reg ( .D(
        new_AGEMA_signal_3867), .CK(clk), .Q(new_AGEMA_signal_3868) );
  DFF_X1 new_AGEMA_reg_buffer_1984_s_current_state_reg ( .D(
        new_AGEMA_signal_3871), .CK(clk), .Q(new_AGEMA_signal_3872) );
  DFF_X1 new_AGEMA_reg_buffer_1988_s_current_state_reg ( .D(
        new_AGEMA_signal_3875), .CK(clk), .Q(new_AGEMA_signal_3876) );
  DFF_X1 new_AGEMA_reg_buffer_1992_s_current_state_reg ( .D(
        new_AGEMA_signal_3879), .CK(clk), .Q(new_AGEMA_signal_3880) );
  DFF_X1 new_AGEMA_reg_buffer_1996_s_current_state_reg ( .D(
        new_AGEMA_signal_3883), .CK(clk), .Q(new_AGEMA_signal_3884) );
  DFF_X1 new_AGEMA_reg_buffer_2000_s_current_state_reg ( .D(
        new_AGEMA_signal_3887), .CK(clk), .Q(new_AGEMA_signal_3888) );
  DFF_X1 new_AGEMA_reg_buffer_2004_s_current_state_reg ( .D(
        new_AGEMA_signal_3891), .CK(clk), .Q(new_AGEMA_signal_3892) );
  DFF_X1 new_AGEMA_reg_buffer_2008_s_current_state_reg ( .D(
        new_AGEMA_signal_3895), .CK(clk), .Q(new_AGEMA_signal_3896) );
  DFF_X1 new_AGEMA_reg_buffer_2012_s_current_state_reg ( .D(
        new_AGEMA_signal_3899), .CK(clk), .Q(new_AGEMA_signal_3900) );
  DFF_X1 new_AGEMA_reg_buffer_2016_s_current_state_reg ( .D(
        new_AGEMA_signal_3903), .CK(clk), .Q(new_AGEMA_signal_3904) );
  DFF_X1 new_AGEMA_reg_buffer_2020_s_current_state_reg ( .D(
        new_AGEMA_signal_3907), .CK(clk), .Q(new_AGEMA_signal_3908) );
  DFF_X1 new_AGEMA_reg_buffer_2024_s_current_state_reg ( .D(
        new_AGEMA_signal_3911), .CK(clk), .Q(new_AGEMA_signal_3912) );
  DFF_X1 new_AGEMA_reg_buffer_2028_s_current_state_reg ( .D(
        new_AGEMA_signal_3915), .CK(clk), .Q(new_AGEMA_signal_3916) );
  DFF_X1 new_AGEMA_reg_buffer_2032_s_current_state_reg ( .D(
        new_AGEMA_signal_3919), .CK(clk), .Q(new_AGEMA_signal_3920) );
  DFF_X1 new_AGEMA_reg_buffer_2036_s_current_state_reg ( .D(
        new_AGEMA_signal_3923), .CK(clk), .Q(new_AGEMA_signal_3924) );
  DFF_X1 new_AGEMA_reg_buffer_2040_s_current_state_reg ( .D(
        new_AGEMA_signal_3927), .CK(clk), .Q(new_AGEMA_signal_3928) );
  DFF_X1 new_AGEMA_reg_buffer_2044_s_current_state_reg ( .D(
        new_AGEMA_signal_3931), .CK(clk), .Q(new_AGEMA_signal_3932) );
  DFF_X1 new_AGEMA_reg_buffer_2048_s_current_state_reg ( .D(
        new_AGEMA_signal_3935), .CK(clk), .Q(new_AGEMA_signal_3936) );
  DFF_X1 new_AGEMA_reg_buffer_2052_s_current_state_reg ( .D(
        new_AGEMA_signal_3939), .CK(clk), .Q(new_AGEMA_signal_3940) );
  DFF_X1 new_AGEMA_reg_buffer_2056_s_current_state_reg ( .D(
        new_AGEMA_signal_3943), .CK(clk), .Q(new_AGEMA_signal_3944) );
  DFF_X1 new_AGEMA_reg_buffer_2060_s_current_state_reg ( .D(
        new_AGEMA_signal_3947), .CK(clk), .Q(new_AGEMA_signal_3948) );
  DFF_X1 new_AGEMA_reg_buffer_2064_s_current_state_reg ( .D(
        new_AGEMA_signal_3951), .CK(clk), .Q(new_AGEMA_signal_3952) );
  DFF_X1 new_AGEMA_reg_buffer_2068_s_current_state_reg ( .D(
        new_AGEMA_signal_3955), .CK(clk), .Q(new_AGEMA_signal_3956) );
  DFF_X1 new_AGEMA_reg_buffer_2072_s_current_state_reg ( .D(
        new_AGEMA_signal_3959), .CK(clk), .Q(new_AGEMA_signal_3960) );
  DFF_X1 new_AGEMA_reg_buffer_2076_s_current_state_reg ( .D(
        new_AGEMA_signal_3963), .CK(clk), .Q(new_AGEMA_signal_3964) );
  DFF_X1 new_AGEMA_reg_buffer_2080_s_current_state_reg ( .D(
        new_AGEMA_signal_3967), .CK(clk), .Q(new_AGEMA_signal_3968) );
  DFF_X1 new_AGEMA_reg_buffer_2084_s_current_state_reg ( .D(
        new_AGEMA_signal_3971), .CK(clk), .Q(new_AGEMA_signal_3972) );
  DFF_X1 new_AGEMA_reg_buffer_2088_s_current_state_reg ( .D(
        new_AGEMA_signal_3975), .CK(clk), .Q(new_AGEMA_signal_3976) );
  DFF_X1 new_AGEMA_reg_buffer_2092_s_current_state_reg ( .D(
        new_AGEMA_signal_3979), .CK(clk), .Q(new_AGEMA_signal_3980) );
  DFF_X1 new_AGEMA_reg_buffer_2096_s_current_state_reg ( .D(
        new_AGEMA_signal_3983), .CK(clk), .Q(new_AGEMA_signal_3984) );
  DFF_X1 new_AGEMA_reg_buffer_2100_s_current_state_reg ( .D(
        new_AGEMA_signal_3987), .CK(clk), .Q(new_AGEMA_signal_3988) );
  DFF_X1 new_AGEMA_reg_buffer_2104_s_current_state_reg ( .D(
        new_AGEMA_signal_3991), .CK(clk), .Q(new_AGEMA_signal_3992) );
  DFF_X1 new_AGEMA_reg_buffer_2108_s_current_state_reg ( .D(
        new_AGEMA_signal_3995), .CK(clk), .Q(new_AGEMA_signal_3996) );
  DFF_X1 new_AGEMA_reg_buffer_2112_s_current_state_reg ( .D(
        new_AGEMA_signal_3999), .CK(clk), .Q(new_AGEMA_signal_4000) );
  DFF_X1 new_AGEMA_reg_buffer_2116_s_current_state_reg ( .D(
        new_AGEMA_signal_4003), .CK(clk), .Q(new_AGEMA_signal_4004) );
  DFF_X1 new_AGEMA_reg_buffer_2120_s_current_state_reg ( .D(
        new_AGEMA_signal_4007), .CK(clk), .Q(new_AGEMA_signal_4008) );
  DFF_X1 new_AGEMA_reg_buffer_2124_s_current_state_reg ( .D(
        new_AGEMA_signal_4011), .CK(clk), .Q(new_AGEMA_signal_4012) );
  DFF_X1 new_AGEMA_reg_buffer_2128_s_current_state_reg ( .D(
        new_AGEMA_signal_4015), .CK(clk), .Q(new_AGEMA_signal_4016) );
  DFF_X1 new_AGEMA_reg_buffer_2132_s_current_state_reg ( .D(
        new_AGEMA_signal_4019), .CK(clk), .Q(new_AGEMA_signal_4020) );
  DFF_X1 new_AGEMA_reg_buffer_2136_s_current_state_reg ( .D(
        new_AGEMA_signal_4023), .CK(clk), .Q(new_AGEMA_signal_4024) );
  DFF_X1 new_AGEMA_reg_buffer_2140_s_current_state_reg ( .D(
        new_AGEMA_signal_4027), .CK(clk), .Q(new_AGEMA_signal_4028) );
  DFF_X1 new_AGEMA_reg_buffer_2144_s_current_state_reg ( .D(
        new_AGEMA_signal_4031), .CK(clk), .Q(new_AGEMA_signal_4032) );
  DFF_X1 new_AGEMA_reg_buffer_2148_s_current_state_reg ( .D(
        new_AGEMA_signal_4035), .CK(clk), .Q(new_AGEMA_signal_4036) );
  DFF_X1 new_AGEMA_reg_buffer_2152_s_current_state_reg ( .D(
        new_AGEMA_signal_4039), .CK(clk), .Q(new_AGEMA_signal_4040) );
  DFF_X1 new_AGEMA_reg_buffer_2156_s_current_state_reg ( .D(
        new_AGEMA_signal_4043), .CK(clk), .Q(new_AGEMA_signal_4044) );
  DFF_X1 new_AGEMA_reg_buffer_2160_s_current_state_reg ( .D(
        new_AGEMA_signal_4047), .CK(clk), .Q(new_AGEMA_signal_4048) );
  DFF_X1 new_AGEMA_reg_buffer_2164_s_current_state_reg ( .D(
        new_AGEMA_signal_4051), .CK(clk), .Q(new_AGEMA_signal_4052) );
  DFF_X1 new_AGEMA_reg_buffer_2168_s_current_state_reg ( .D(
        new_AGEMA_signal_4055), .CK(clk), .Q(new_AGEMA_signal_4056) );
  DFF_X1 new_AGEMA_reg_buffer_2172_s_current_state_reg ( .D(
        new_AGEMA_signal_4059), .CK(clk), .Q(new_AGEMA_signal_4060) );
  DFF_X1 new_AGEMA_reg_buffer_2176_s_current_state_reg ( .D(
        new_AGEMA_signal_4063), .CK(clk), .Q(new_AGEMA_signal_4064) );
  DFF_X1 new_AGEMA_reg_buffer_2180_s_current_state_reg ( .D(
        new_AGEMA_signal_4067), .CK(clk), .Q(new_AGEMA_signal_4068) );
  DFF_X1 new_AGEMA_reg_buffer_2184_s_current_state_reg ( .D(
        new_AGEMA_signal_4071), .CK(clk), .Q(new_AGEMA_signal_4072) );
  DFF_X1 new_AGEMA_reg_buffer_2188_s_current_state_reg ( .D(
        new_AGEMA_signal_4075), .CK(clk), .Q(new_AGEMA_signal_4076) );
  DFF_X1 new_AGEMA_reg_buffer_2192_s_current_state_reg ( .D(
        new_AGEMA_signal_4079), .CK(clk), .Q(new_AGEMA_signal_4080) );
  DFF_X1 new_AGEMA_reg_buffer_2196_s_current_state_reg ( .D(
        new_AGEMA_signal_4083), .CK(clk), .Q(new_AGEMA_signal_4084) );
  DFF_X1 new_AGEMA_reg_buffer_2200_s_current_state_reg ( .D(
        new_AGEMA_signal_4087), .CK(clk), .Q(new_AGEMA_signal_4088) );
  DFF_X1 new_AGEMA_reg_buffer_2204_s_current_state_reg ( .D(
        new_AGEMA_signal_4091), .CK(clk), .Q(new_AGEMA_signal_4092) );
  DFF_X1 new_AGEMA_reg_buffer_2208_s_current_state_reg ( .D(
        new_AGEMA_signal_4095), .CK(clk), .Q(new_AGEMA_signal_4096) );
  DFF_X1 new_AGEMA_reg_buffer_2212_s_current_state_reg ( .D(
        new_AGEMA_signal_4099), .CK(clk), .Q(new_AGEMA_signal_4100) );
  DFF_X1 new_AGEMA_reg_buffer_2216_s_current_state_reg ( .D(
        new_AGEMA_signal_4103), .CK(clk), .Q(new_AGEMA_signal_4104) );
  DFF_X1 new_AGEMA_reg_buffer_2220_s_current_state_reg ( .D(
        new_AGEMA_signal_4107), .CK(clk), .Q(new_AGEMA_signal_4108) );
  DFF_X1 new_AGEMA_reg_buffer_2224_s_current_state_reg ( .D(
        new_AGEMA_signal_4111), .CK(clk), .Q(new_AGEMA_signal_4112) );
  DFF_X1 new_AGEMA_reg_buffer_2228_s_current_state_reg ( .D(
        new_AGEMA_signal_4115), .CK(clk), .Q(new_AGEMA_signal_4116) );
  DFF_X1 new_AGEMA_reg_buffer_2232_s_current_state_reg ( .D(
        new_AGEMA_signal_4119), .CK(clk), .Q(new_AGEMA_signal_4120) );
  DFF_X1 new_AGEMA_reg_buffer_2236_s_current_state_reg ( .D(
        new_AGEMA_signal_4123), .CK(clk), .Q(new_AGEMA_signal_4124) );
  DFF_X1 new_AGEMA_reg_buffer_2240_s_current_state_reg ( .D(
        new_AGEMA_signal_4127), .CK(clk), .Q(new_AGEMA_signal_4128) );
  DFF_X1 new_AGEMA_reg_buffer_2244_s_current_state_reg ( .D(
        new_AGEMA_signal_4131), .CK(clk), .Q(new_AGEMA_signal_4132) );
  DFF_X1 new_AGEMA_reg_buffer_2247_s_current_state_reg ( .D(
        new_AGEMA_signal_4134), .CK(clk), .Q(new_AGEMA_signal_4135) );
  DFF_X1 new_AGEMA_reg_buffer_2250_s_current_state_reg ( .D(
        new_AGEMA_signal_4137), .CK(clk), .Q(new_AGEMA_signal_4138) );
  DFF_X1 new_AGEMA_reg_buffer_2253_s_current_state_reg ( .D(
        new_AGEMA_signal_4140), .CK(clk), .Q(new_AGEMA_signal_4141) );
  DFF_X1 new_AGEMA_reg_buffer_2256_s_current_state_reg ( .D(
        new_AGEMA_signal_4143), .CK(clk), .Q(new_AGEMA_signal_4144) );
  DFF_X1 new_AGEMA_reg_buffer_2259_s_current_state_reg ( .D(
        new_AGEMA_signal_4146), .CK(clk), .Q(new_AGEMA_signal_4147) );
  DFF_X1 new_AGEMA_reg_buffer_2262_s_current_state_reg ( .D(
        new_AGEMA_signal_4149), .CK(clk), .Q(new_AGEMA_signal_4150) );
  DFF_X1 new_AGEMA_reg_buffer_2265_s_current_state_reg ( .D(
        new_AGEMA_signal_4152), .CK(clk), .Q(new_AGEMA_signal_4153) );
  DFF_X1 new_AGEMA_reg_buffer_2268_s_current_state_reg ( .D(
        new_AGEMA_signal_4155), .CK(clk), .Q(new_AGEMA_signal_4156) );
  DFF_X1 new_AGEMA_reg_buffer_2271_s_current_state_reg ( .D(
        new_AGEMA_signal_4158), .CK(clk), .Q(new_AGEMA_signal_4159) );
  DFF_X1 new_AGEMA_reg_buffer_2274_s_current_state_reg ( .D(
        new_AGEMA_signal_4161), .CK(clk), .Q(new_AGEMA_signal_4162) );
  DFF_X1 new_AGEMA_reg_buffer_2277_s_current_state_reg ( .D(
        new_AGEMA_signal_4164), .CK(clk), .Q(new_AGEMA_signal_4165) );
  DFF_X1 new_AGEMA_reg_buffer_2280_s_current_state_reg ( .D(
        new_AGEMA_signal_4167), .CK(clk), .Q(new_AGEMA_signal_4168) );
  DFF_X1 new_AGEMA_reg_buffer_2283_s_current_state_reg ( .D(
        new_AGEMA_signal_4170), .CK(clk), .Q(new_AGEMA_signal_4171) );
  DFF_X1 new_AGEMA_reg_buffer_2286_s_current_state_reg ( .D(
        new_AGEMA_signal_4173), .CK(clk), .Q(new_AGEMA_signal_4174) );
  DFF_X1 new_AGEMA_reg_buffer_2289_s_current_state_reg ( .D(
        new_AGEMA_signal_4176), .CK(clk), .Q(new_AGEMA_signal_4177) );
  DFF_X1 new_AGEMA_reg_buffer_2292_s_current_state_reg ( .D(
        new_AGEMA_signal_4179), .CK(clk), .Q(new_AGEMA_signal_4180) );
  DFF_X1 new_AGEMA_reg_buffer_2295_s_current_state_reg ( .D(
        new_AGEMA_signal_4182), .CK(clk), .Q(new_AGEMA_signal_4183) );
  DFF_X1 new_AGEMA_reg_buffer_2298_s_current_state_reg ( .D(
        new_AGEMA_signal_4185), .CK(clk), .Q(new_AGEMA_signal_4186) );
  DFF_X1 new_AGEMA_reg_buffer_2301_s_current_state_reg ( .D(
        new_AGEMA_signal_4188), .CK(clk), .Q(new_AGEMA_signal_4189) );
  DFF_X1 new_AGEMA_reg_buffer_2304_s_current_state_reg ( .D(
        new_AGEMA_signal_4191), .CK(clk), .Q(new_AGEMA_signal_4192) );
  DFF_X1 new_AGEMA_reg_buffer_2307_s_current_state_reg ( .D(
        new_AGEMA_signal_4194), .CK(clk), .Q(new_AGEMA_signal_4195) );
  DFF_X1 new_AGEMA_reg_buffer_2310_s_current_state_reg ( .D(
        new_AGEMA_signal_4197), .CK(clk), .Q(new_AGEMA_signal_4198) );
  DFF_X1 new_AGEMA_reg_buffer_2313_s_current_state_reg ( .D(
        new_AGEMA_signal_4200), .CK(clk), .Q(new_AGEMA_signal_4201) );
  DFF_X1 new_AGEMA_reg_buffer_2316_s_current_state_reg ( .D(
        new_AGEMA_signal_4203), .CK(clk), .Q(new_AGEMA_signal_4204) );
  DFF_X1 new_AGEMA_reg_buffer_2319_s_current_state_reg ( .D(
        new_AGEMA_signal_4206), .CK(clk), .Q(new_AGEMA_signal_4207) );
  DFF_X1 new_AGEMA_reg_buffer_2322_s_current_state_reg ( .D(
        new_AGEMA_signal_4209), .CK(clk), .Q(new_AGEMA_signal_4210) );
  DFF_X1 new_AGEMA_reg_buffer_2325_s_current_state_reg ( .D(
        new_AGEMA_signal_4212), .CK(clk), .Q(new_AGEMA_signal_4213) );
  DFF_X1 new_AGEMA_reg_buffer_2328_s_current_state_reg ( .D(
        new_AGEMA_signal_4215), .CK(clk), .Q(new_AGEMA_signal_4216) );
  DFF_X1 new_AGEMA_reg_buffer_2331_s_current_state_reg ( .D(
        new_AGEMA_signal_4218), .CK(clk), .Q(new_AGEMA_signal_4219) );
  DFF_X1 new_AGEMA_reg_buffer_2334_s_current_state_reg ( .D(
        new_AGEMA_signal_4221), .CK(clk), .Q(new_AGEMA_signal_4222) );
  DFF_X1 new_AGEMA_reg_buffer_2337_s_current_state_reg ( .D(
        new_AGEMA_signal_4224), .CK(clk), .Q(new_AGEMA_signal_4225) );
  DFF_X1 new_AGEMA_reg_buffer_2340_s_current_state_reg ( .D(
        new_AGEMA_signal_4227), .CK(clk), .Q(new_AGEMA_signal_4228) );
  DFF_X1 new_AGEMA_reg_buffer_2343_s_current_state_reg ( .D(
        new_AGEMA_signal_4230), .CK(clk), .Q(new_AGEMA_signal_4231) );
  DFF_X1 new_AGEMA_reg_buffer_2346_s_current_state_reg ( .D(
        new_AGEMA_signal_4233), .CK(clk), .Q(new_AGEMA_signal_4234) );
  DFF_X1 new_AGEMA_reg_buffer_2349_s_current_state_reg ( .D(
        new_AGEMA_signal_4236), .CK(clk), .Q(new_AGEMA_signal_4237) );
  DFF_X1 new_AGEMA_reg_buffer_2352_s_current_state_reg ( .D(
        new_AGEMA_signal_4239), .CK(clk), .Q(new_AGEMA_signal_4240) );
  DFF_X1 new_AGEMA_reg_buffer_2356_s_current_state_reg ( .D(
        new_AGEMA_signal_4243), .CK(clk), .Q(new_AGEMA_signal_4244) );
  DFF_X1 new_AGEMA_reg_buffer_2360_s_current_state_reg ( .D(
        new_AGEMA_signal_4247), .CK(clk), .Q(new_AGEMA_signal_4248) );
  DFF_X1 new_AGEMA_reg_buffer_2364_s_current_state_reg ( .D(
        new_AGEMA_signal_4251), .CK(clk), .Q(new_AGEMA_signal_4252) );
  DFF_X1 new_AGEMA_reg_buffer_2368_s_current_state_reg ( .D(
        new_AGEMA_signal_4255), .CK(clk), .Q(new_AGEMA_signal_4256) );
  DFF_X1 new_AGEMA_reg_buffer_2372_s_current_state_reg ( .D(
        new_AGEMA_signal_4259), .CK(clk), .Q(new_AGEMA_signal_4260) );
  DFF_X1 new_AGEMA_reg_buffer_2376_s_current_state_reg ( .D(
        new_AGEMA_signal_4263), .CK(clk), .Q(new_AGEMA_signal_4264) );
  DFF_X1 new_AGEMA_reg_buffer_2380_s_current_state_reg ( .D(
        new_AGEMA_signal_4267), .CK(clk), .Q(new_AGEMA_signal_4268) );
  DFF_X1 new_AGEMA_reg_buffer_2384_s_current_state_reg ( .D(
        new_AGEMA_signal_4271), .CK(clk), .Q(new_AGEMA_signal_4272) );
  DFF_X1 new_AGEMA_reg_buffer_2388_s_current_state_reg ( .D(
        new_AGEMA_signal_4275), .CK(clk), .Q(new_AGEMA_signal_4276) );
  DFF_X1 new_AGEMA_reg_buffer_2392_s_current_state_reg ( .D(
        new_AGEMA_signal_4279), .CK(clk), .Q(new_AGEMA_signal_4280) );
  DFF_X1 new_AGEMA_reg_buffer_2396_s_current_state_reg ( .D(
        new_AGEMA_signal_4283), .CK(clk), .Q(new_AGEMA_signal_4284) );
  DFF_X1 new_AGEMA_reg_buffer_2400_s_current_state_reg ( .D(
        new_AGEMA_signal_4287), .CK(clk), .Q(new_AGEMA_signal_4288) );
  DFF_X1 new_AGEMA_reg_buffer_2404_s_current_state_reg ( .D(
        new_AGEMA_signal_4291), .CK(clk), .Q(new_AGEMA_signal_4292) );
  DFF_X1 new_AGEMA_reg_buffer_2408_s_current_state_reg ( .D(
        new_AGEMA_signal_4295), .CK(clk), .Q(new_AGEMA_signal_4296) );
  DFF_X1 new_AGEMA_reg_buffer_2412_s_current_state_reg ( .D(
        new_AGEMA_signal_4299), .CK(clk), .Q(new_AGEMA_signal_4300) );
  DFF_X1 new_AGEMA_reg_buffer_2416_s_current_state_reg ( .D(
        new_AGEMA_signal_4303), .CK(clk), .Q(new_AGEMA_signal_4304) );
  DFF_X1 new_AGEMA_reg_buffer_2420_s_current_state_reg ( .D(
        new_AGEMA_signal_4307), .CK(clk), .Q(new_AGEMA_signal_4308) );
  DFF_X1 new_AGEMA_reg_buffer_2424_s_current_state_reg ( .D(
        new_AGEMA_signal_4311), .CK(clk), .Q(new_AGEMA_signal_4312) );
  DFF_X1 new_AGEMA_reg_buffer_2428_s_current_state_reg ( .D(
        new_AGEMA_signal_4315), .CK(clk), .Q(new_AGEMA_signal_4316) );
  DFF_X1 new_AGEMA_reg_buffer_2432_s_current_state_reg ( .D(
        new_AGEMA_signal_4319), .CK(clk), .Q(new_AGEMA_signal_4320) );
  DFF_X1 new_AGEMA_reg_buffer_2436_s_current_state_reg ( .D(
        new_AGEMA_signal_4323), .CK(clk), .Q(new_AGEMA_signal_4324) );
  DFF_X1 new_AGEMA_reg_buffer_2440_s_current_state_reg ( .D(
        new_AGEMA_signal_4327), .CK(clk), .Q(new_AGEMA_signal_4328) );
  DFF_X1 new_AGEMA_reg_buffer_2444_s_current_state_reg ( .D(
        new_AGEMA_signal_4331), .CK(clk), .Q(new_AGEMA_signal_4332) );
  DFF_X1 new_AGEMA_reg_buffer_2448_s_current_state_reg ( .D(
        new_AGEMA_signal_4335), .CK(clk), .Q(new_AGEMA_signal_4336) );
  DFF_X1 new_AGEMA_reg_buffer_2452_s_current_state_reg ( .D(
        new_AGEMA_signal_4339), .CK(clk), .Q(new_AGEMA_signal_4340) );
  DFF_X1 new_AGEMA_reg_buffer_2456_s_current_state_reg ( .D(
        new_AGEMA_signal_4343), .CK(clk), .Q(new_AGEMA_signal_4344) );
  DFF_X1 new_AGEMA_reg_buffer_2460_s_current_state_reg ( .D(
        new_AGEMA_signal_4347), .CK(clk), .Q(new_AGEMA_signal_4348) );
  DFF_X1 new_AGEMA_reg_buffer_2464_s_current_state_reg ( .D(
        new_AGEMA_signal_4351), .CK(clk), .Q(new_AGEMA_signal_4352) );
  DFF_X1 new_AGEMA_reg_buffer_2468_s_current_state_reg ( .D(
        new_AGEMA_signal_4355), .CK(clk), .Q(new_AGEMA_signal_4356) );
  DFF_X1 new_AGEMA_reg_buffer_2472_s_current_state_reg ( .D(
        new_AGEMA_signal_4359), .CK(clk), .Q(new_AGEMA_signal_4360) );
  DFF_X1 new_AGEMA_reg_buffer_2476_s_current_state_reg ( .D(
        new_AGEMA_signal_4363), .CK(clk), .Q(new_AGEMA_signal_4364) );
  DFF_X1 new_AGEMA_reg_buffer_2480_s_current_state_reg ( .D(
        new_AGEMA_signal_4367), .CK(clk), .Q(new_AGEMA_signal_4368) );
  DFF_X1 new_AGEMA_reg_buffer_2484_s_current_state_reg ( .D(
        new_AGEMA_signal_4371), .CK(clk), .Q(new_AGEMA_signal_4372) );
  DFF_X1 new_AGEMA_reg_buffer_2488_s_current_state_reg ( .D(
        new_AGEMA_signal_4375), .CK(clk), .Q(new_AGEMA_signal_4376) );
  DFF_X1 new_AGEMA_reg_buffer_2492_s_current_state_reg ( .D(
        new_AGEMA_signal_4379), .CK(clk), .Q(new_AGEMA_signal_4380) );
  DFF_X1 new_AGEMA_reg_buffer_2496_s_current_state_reg ( .D(
        new_AGEMA_signal_4383), .CK(clk), .Q(new_AGEMA_signal_4384) );
  DFF_X1 new_AGEMA_reg_buffer_2500_s_current_state_reg ( .D(
        new_AGEMA_signal_4387), .CK(clk), .Q(new_AGEMA_signal_4388) );
  DFF_X1 new_AGEMA_reg_buffer_2504_s_current_state_reg ( .D(
        new_AGEMA_signal_4391), .CK(clk), .Q(new_AGEMA_signal_4392) );
  DFF_X1 new_AGEMA_reg_buffer_2508_s_current_state_reg ( .D(
        new_AGEMA_signal_4395), .CK(clk), .Q(new_AGEMA_signal_4396) );
  DFF_X1 new_AGEMA_reg_buffer_2512_s_current_state_reg ( .D(
        new_AGEMA_signal_4399), .CK(clk), .Q(new_AGEMA_signal_4400) );
  DFF_X1 new_AGEMA_reg_buffer_2516_s_current_state_reg ( .D(
        new_AGEMA_signal_4403), .CK(clk), .Q(new_AGEMA_signal_4404) );
  DFF_X1 new_AGEMA_reg_buffer_2520_s_current_state_reg ( .D(
        new_AGEMA_signal_4407), .CK(clk), .Q(new_AGEMA_signal_4408) );
  DFF_X1 new_AGEMA_reg_buffer_2524_s_current_state_reg ( .D(
        new_AGEMA_signal_4411), .CK(clk), .Q(new_AGEMA_signal_4412) );
  DFF_X1 new_AGEMA_reg_buffer_2528_s_current_state_reg ( .D(
        new_AGEMA_signal_4415), .CK(clk), .Q(new_AGEMA_signal_4416) );
  DFF_X1 new_AGEMA_reg_buffer_2532_s_current_state_reg ( .D(
        new_AGEMA_signal_4419), .CK(clk), .Q(new_AGEMA_signal_4420) );
  DFF_X1 new_AGEMA_reg_buffer_2536_s_current_state_reg ( .D(
        new_AGEMA_signal_4423), .CK(clk), .Q(new_AGEMA_signal_4424) );
  DFF_X1 new_AGEMA_reg_buffer_2540_s_current_state_reg ( .D(
        new_AGEMA_signal_4427), .CK(clk), .Q(new_AGEMA_signal_4428) );
  DFF_X1 new_AGEMA_reg_buffer_2544_s_current_state_reg ( .D(
        new_AGEMA_signal_4431), .CK(clk), .Q(new_AGEMA_signal_4432) );
  DFF_X1 new_AGEMA_reg_buffer_2548_s_current_state_reg ( .D(
        new_AGEMA_signal_4435), .CK(clk), .Q(new_AGEMA_signal_4436) );
  DFF_X1 new_AGEMA_reg_buffer_2552_s_current_state_reg ( .D(
        new_AGEMA_signal_4439), .CK(clk), .Q(new_AGEMA_signal_4440) );
  DFF_X1 new_AGEMA_reg_buffer_2556_s_current_state_reg ( .D(
        new_AGEMA_signal_4443), .CK(clk), .Q(new_AGEMA_signal_4444) );
  DFF_X1 new_AGEMA_reg_buffer_2560_s_current_state_reg ( .D(
        new_AGEMA_signal_4447), .CK(clk), .Q(new_AGEMA_signal_4448) );
  DFF_X1 new_AGEMA_reg_buffer_2564_s_current_state_reg ( .D(
        new_AGEMA_signal_4451), .CK(clk), .Q(new_AGEMA_signal_4452) );
  DFF_X1 new_AGEMA_reg_buffer_2568_s_current_state_reg ( .D(
        new_AGEMA_signal_4455), .CK(clk), .Q(new_AGEMA_signal_4456) );
  DFF_X1 new_AGEMA_reg_buffer_2572_s_current_state_reg ( .D(
        new_AGEMA_signal_4459), .CK(clk), .Q(new_AGEMA_signal_4460) );
  DFF_X1 new_AGEMA_reg_buffer_2576_s_current_state_reg ( .D(
        new_AGEMA_signal_4463), .CK(clk), .Q(new_AGEMA_signal_4464) );
  DFF_X1 new_AGEMA_reg_buffer_2580_s_current_state_reg ( .D(
        new_AGEMA_signal_4467), .CK(clk), .Q(new_AGEMA_signal_4468) );
  DFF_X1 new_AGEMA_reg_buffer_2584_s_current_state_reg ( .D(
        new_AGEMA_signal_4471), .CK(clk), .Q(new_AGEMA_signal_4472) );
  DFF_X1 new_AGEMA_reg_buffer_2588_s_current_state_reg ( .D(
        new_AGEMA_signal_4475), .CK(clk), .Q(new_AGEMA_signal_4476) );
  DFF_X1 new_AGEMA_reg_buffer_2592_s_current_state_reg ( .D(
        new_AGEMA_signal_4479), .CK(clk), .Q(new_AGEMA_signal_4480) );
  DFF_X1 new_AGEMA_reg_buffer_2596_s_current_state_reg ( .D(
        new_AGEMA_signal_4483), .CK(clk), .Q(new_AGEMA_signal_4484) );
  DFF_X1 new_AGEMA_reg_buffer_2600_s_current_state_reg ( .D(
        new_AGEMA_signal_4487), .CK(clk), .Q(new_AGEMA_signal_4488) );
  DFF_X1 new_AGEMA_reg_buffer_2604_s_current_state_reg ( .D(
        new_AGEMA_signal_4491), .CK(clk), .Q(new_AGEMA_signal_4492) );
  DFF_X1 new_AGEMA_reg_buffer_2608_s_current_state_reg ( .D(
        new_AGEMA_signal_4495), .CK(clk), .Q(new_AGEMA_signal_4496) );
  DFF_X1 new_AGEMA_reg_buffer_2612_s_current_state_reg ( .D(
        new_AGEMA_signal_4499), .CK(clk), .Q(new_AGEMA_signal_4500) );
  DFF_X1 new_AGEMA_reg_buffer_2616_s_current_state_reg ( .D(
        new_AGEMA_signal_4503), .CK(clk), .Q(new_AGEMA_signal_4504) );
  DFF_X1 new_AGEMA_reg_buffer_2620_s_current_state_reg ( .D(
        new_AGEMA_signal_4507), .CK(clk), .Q(new_AGEMA_signal_4508) );
  DFF_X1 new_AGEMA_reg_buffer_2624_s_current_state_reg ( .D(
        new_AGEMA_signal_4511), .CK(clk), .Q(new_AGEMA_signal_4512) );
  DFF_X1 new_AGEMA_reg_buffer_2628_s_current_state_reg ( .D(
        new_AGEMA_signal_4515), .CK(clk), .Q(new_AGEMA_signal_4516) );
  DFF_X1 new_AGEMA_reg_buffer_2632_s_current_state_reg ( .D(
        new_AGEMA_signal_4519), .CK(clk), .Q(new_AGEMA_signal_4520) );
  DFF_X1 new_AGEMA_reg_buffer_2636_s_current_state_reg ( .D(
        new_AGEMA_signal_4523), .CK(clk), .Q(new_AGEMA_signal_4524) );
  DFF_X1 new_AGEMA_reg_buffer_2640_s_current_state_reg ( .D(
        new_AGEMA_signal_4527), .CK(clk), .Q(new_AGEMA_signal_4528) );
  DFF_X1 new_AGEMA_reg_buffer_2644_s_current_state_reg ( .D(
        new_AGEMA_signal_4531), .CK(clk), .Q(new_AGEMA_signal_4532) );
  DFF_X1 new_AGEMA_reg_buffer_2648_s_current_state_reg ( .D(
        new_AGEMA_signal_4535), .CK(clk), .Q(new_AGEMA_signal_4536) );
  DFF_X1 new_AGEMA_reg_buffer_2652_s_current_state_reg ( .D(
        new_AGEMA_signal_4539), .CK(clk), .Q(new_AGEMA_signal_4540) );
  DFF_X1 new_AGEMA_reg_buffer_2656_s_current_state_reg ( .D(
        new_AGEMA_signal_4543), .CK(clk), .Q(new_AGEMA_signal_4544) );
  DFF_X1 new_AGEMA_reg_buffer_2660_s_current_state_reg ( .D(
        new_AGEMA_signal_4547), .CK(clk), .Q(new_AGEMA_signal_4548) );
  DFF_X1 new_AGEMA_reg_buffer_2664_s_current_state_reg ( .D(
        new_AGEMA_signal_4551), .CK(clk), .Q(new_AGEMA_signal_4552) );
  DFF_X1 new_AGEMA_reg_buffer_2668_s_current_state_reg ( .D(
        new_AGEMA_signal_4555), .CK(clk), .Q(new_AGEMA_signal_4556) );
  DFF_X1 new_AGEMA_reg_buffer_2672_s_current_state_reg ( .D(
        new_AGEMA_signal_4559), .CK(clk), .Q(new_AGEMA_signal_4560) );
  DFF_X1 new_AGEMA_reg_buffer_2676_s_current_state_reg ( .D(
        new_AGEMA_signal_4563), .CK(clk), .Q(new_AGEMA_signal_4564) );
  DFF_X1 new_AGEMA_reg_buffer_2680_s_current_state_reg ( .D(
        new_AGEMA_signal_4567), .CK(clk), .Q(new_AGEMA_signal_4568) );
  DFF_X1 new_AGEMA_reg_buffer_2684_s_current_state_reg ( .D(
        new_AGEMA_signal_4571), .CK(clk), .Q(new_AGEMA_signal_4572) );
  DFF_X1 new_AGEMA_reg_buffer_2688_s_current_state_reg ( .D(
        new_AGEMA_signal_4575), .CK(clk), .Q(new_AGEMA_signal_4576) );
  DFF_X1 new_AGEMA_reg_buffer_2692_s_current_state_reg ( .D(
        new_AGEMA_signal_4579), .CK(clk), .Q(new_AGEMA_signal_4580) );
  DFF_X1 new_AGEMA_reg_buffer_2696_s_current_state_reg ( .D(
        new_AGEMA_signal_4583), .CK(clk), .Q(new_AGEMA_signal_4584) );
  DFF_X1 new_AGEMA_reg_buffer_2700_s_current_state_reg ( .D(
        new_AGEMA_signal_4587), .CK(clk), .Q(new_AGEMA_signal_4588) );
  DFF_X1 new_AGEMA_reg_buffer_2704_s_current_state_reg ( .D(
        new_AGEMA_signal_4591), .CK(clk), .Q(new_AGEMA_signal_4592) );
  DFF_X1 new_AGEMA_reg_buffer_2708_s_current_state_reg ( .D(
        new_AGEMA_signal_4595), .CK(clk), .Q(new_AGEMA_signal_4596) );
  DFF_X1 new_AGEMA_reg_buffer_2712_s_current_state_reg ( .D(
        new_AGEMA_signal_4599), .CK(clk), .Q(new_AGEMA_signal_4600) );
  DFF_X1 new_AGEMA_reg_buffer_2716_s_current_state_reg ( .D(
        new_AGEMA_signal_4603), .CK(clk), .Q(new_AGEMA_signal_4604) );
  DFF_X1 new_AGEMA_reg_buffer_2720_s_current_state_reg ( .D(
        new_AGEMA_signal_4607), .CK(clk), .Q(new_AGEMA_signal_4608) );
  DFF_X1 new_AGEMA_reg_buffer_2724_s_current_state_reg ( .D(
        new_AGEMA_signal_4611), .CK(clk), .Q(new_AGEMA_signal_4612) );
  DFF_X1 new_AGEMA_reg_buffer_2728_s_current_state_reg ( .D(
        new_AGEMA_signal_4615), .CK(clk), .Q(new_AGEMA_signal_4616) );
  DFF_X1 new_AGEMA_reg_buffer_2732_s_current_state_reg ( .D(
        new_AGEMA_signal_4619), .CK(clk), .Q(new_AGEMA_signal_4620) );
  DFF_X1 new_AGEMA_reg_buffer_2736_s_current_state_reg ( .D(
        new_AGEMA_signal_4623), .CK(clk), .Q(new_AGEMA_signal_4624) );
  DFF_X1 new_AGEMA_reg_buffer_2740_s_current_state_reg ( .D(
        new_AGEMA_signal_4627), .CK(clk), .Q(new_AGEMA_signal_4628) );
  DFF_X1 new_AGEMA_reg_buffer_2744_s_current_state_reg ( .D(
        new_AGEMA_signal_4631), .CK(clk), .Q(new_AGEMA_signal_4632) );
  DFF_X1 new_AGEMA_reg_buffer_2748_s_current_state_reg ( .D(
        new_AGEMA_signal_4635), .CK(clk), .Q(new_AGEMA_signal_4636) );
  DFF_X1 new_AGEMA_reg_buffer_2752_s_current_state_reg ( .D(
        new_AGEMA_signal_4639), .CK(clk), .Q(new_AGEMA_signal_4640) );
  DFF_X1 new_AGEMA_reg_buffer_2756_s_current_state_reg ( .D(
        new_AGEMA_signal_4643), .CK(clk), .Q(new_AGEMA_signal_4644) );
  DFF_X1 new_AGEMA_reg_buffer_2760_s_current_state_reg ( .D(
        new_AGEMA_signal_4647), .CK(clk), .Q(new_AGEMA_signal_4648) );
  DFF_X1 new_AGEMA_reg_buffer_2764_s_current_state_reg ( .D(
        new_AGEMA_signal_4651), .CK(clk), .Q(new_AGEMA_signal_4652) );
  DFF_X1 new_AGEMA_reg_buffer_2768_s_current_state_reg ( .D(
        new_AGEMA_signal_4655), .CK(clk), .Q(new_AGEMA_signal_4656) );
  DFF_X1 new_AGEMA_reg_buffer_2772_s_current_state_reg ( .D(
        new_AGEMA_signal_4659), .CK(clk), .Q(new_AGEMA_signal_4660) );
  DFF_X1 new_AGEMA_reg_buffer_2776_s_current_state_reg ( .D(
        new_AGEMA_signal_4663), .CK(clk), .Q(new_AGEMA_signal_4664) );
  DFF_X1 new_AGEMA_reg_buffer_2780_s_current_state_reg ( .D(
        new_AGEMA_signal_4667), .CK(clk), .Q(new_AGEMA_signal_4668) );
  DFF_X1 new_AGEMA_reg_buffer_2784_s_current_state_reg ( .D(
        new_AGEMA_signal_4671), .CK(clk), .Q(new_AGEMA_signal_4672) );
  DFF_X1 new_AGEMA_reg_buffer_2788_s_current_state_reg ( .D(
        new_AGEMA_signal_4675), .CK(clk), .Q(new_AGEMA_signal_4676) );
  DFF_X1 new_AGEMA_reg_buffer_2792_s_current_state_reg ( .D(
        new_AGEMA_signal_4679), .CK(clk), .Q(new_AGEMA_signal_4680) );
  DFF_X1 new_AGEMA_reg_buffer_2796_s_current_state_reg ( .D(
        new_AGEMA_signal_4683), .CK(clk), .Q(new_AGEMA_signal_4684) );
  DFF_X1 new_AGEMA_reg_buffer_2800_s_current_state_reg ( .D(
        new_AGEMA_signal_4687), .CK(clk), .Q(new_AGEMA_signal_4688) );
  DFF_X1 new_AGEMA_reg_buffer_2804_s_current_state_reg ( .D(
        new_AGEMA_signal_4691), .CK(clk), .Q(new_AGEMA_signal_4692) );
  DFF_X1 new_AGEMA_reg_buffer_2808_s_current_state_reg ( .D(
        new_AGEMA_signal_4695), .CK(clk), .Q(new_AGEMA_signal_4696) );
  DFF_X1 new_AGEMA_reg_buffer_2812_s_current_state_reg ( .D(
        new_AGEMA_signal_4699), .CK(clk), .Q(new_AGEMA_signal_4700) );
  DFF_X1 new_AGEMA_reg_buffer_2816_s_current_state_reg ( .D(
        new_AGEMA_signal_4703), .CK(clk), .Q(new_AGEMA_signal_4704) );
  DFF_X1 new_AGEMA_reg_buffer_2820_s_current_state_reg ( .D(
        new_AGEMA_signal_4707), .CK(clk), .Q(new_AGEMA_signal_4708) );
  DFF_X1 new_AGEMA_reg_buffer_2824_s_current_state_reg ( .D(
        new_AGEMA_signal_4711), .CK(clk), .Q(new_AGEMA_signal_4712) );
  DFF_X1 new_AGEMA_reg_buffer_2828_s_current_state_reg ( .D(
        new_AGEMA_signal_4715), .CK(clk), .Q(new_AGEMA_signal_4716) );
  DFF_X1 new_AGEMA_reg_buffer_2832_s_current_state_reg ( .D(
        new_AGEMA_signal_4719), .CK(clk), .Q(new_AGEMA_signal_4720) );
  DFF_X1 new_AGEMA_reg_buffer_2836_s_current_state_reg ( .D(
        new_AGEMA_signal_4723), .CK(clk), .Q(new_AGEMA_signal_4724) );
  DFF_X1 new_AGEMA_reg_buffer_2840_s_current_state_reg ( .D(
        new_AGEMA_signal_4727), .CK(clk), .Q(new_AGEMA_signal_4728) );
  DFF_X1 new_AGEMA_reg_buffer_2844_s_current_state_reg ( .D(
        new_AGEMA_signal_4731), .CK(clk), .Q(new_AGEMA_signal_4732) );
  DFF_X1 new_AGEMA_reg_buffer_2848_s_current_state_reg ( .D(
        new_AGEMA_signal_4735), .CK(clk), .Q(new_AGEMA_signal_4736) );
  DFF_X1 new_AGEMA_reg_buffer_2852_s_current_state_reg ( .D(
        new_AGEMA_signal_4739), .CK(clk), .Q(new_AGEMA_signal_4740) );
  DFF_X1 new_AGEMA_reg_buffer_2856_s_current_state_reg ( .D(
        new_AGEMA_signal_4743), .CK(clk), .Q(new_AGEMA_signal_4744) );
  DFF_X1 new_AGEMA_reg_buffer_2860_s_current_state_reg ( .D(
        new_AGEMA_signal_4747), .CK(clk), .Q(new_AGEMA_signal_4748) );
  DFF_X1 new_AGEMA_reg_buffer_2864_s_current_state_reg ( .D(
        new_AGEMA_signal_4751), .CK(clk), .Q(new_AGEMA_signal_4752) );
  DFF_X1 new_AGEMA_reg_buffer_2868_s_current_state_reg ( .D(
        new_AGEMA_signal_4755), .CK(clk), .Q(new_AGEMA_signal_4756) );
  DFF_X1 new_AGEMA_reg_buffer_2872_s_current_state_reg ( .D(
        new_AGEMA_signal_4759), .CK(clk), .Q(new_AGEMA_signal_4760) );
  DFF_X1 new_AGEMA_reg_buffer_2876_s_current_state_reg ( .D(
        new_AGEMA_signal_4763), .CK(clk), .Q(new_AGEMA_signal_4764) );
  DFF_X1 new_AGEMA_reg_buffer_2880_s_current_state_reg ( .D(
        new_AGEMA_signal_4767), .CK(clk), .Q(new_AGEMA_signal_4768) );
  DFF_X1 new_AGEMA_reg_buffer_2884_s_current_state_reg ( .D(
        new_AGEMA_signal_4771), .CK(clk), .Q(new_AGEMA_signal_4772) );
  DFF_X1 new_AGEMA_reg_buffer_2888_s_current_state_reg ( .D(
        new_AGEMA_signal_4775), .CK(clk), .Q(new_AGEMA_signal_4776) );
  DFF_X1 new_AGEMA_reg_buffer_2892_s_current_state_reg ( .D(
        new_AGEMA_signal_4779), .CK(clk), .Q(new_AGEMA_signal_4780) );
  DFF_X1 new_AGEMA_reg_buffer_2896_s_current_state_reg ( .D(
        new_AGEMA_signal_4783), .CK(clk), .Q(new_AGEMA_signal_4784) );
  DFF_X1 new_AGEMA_reg_buffer_2900_s_current_state_reg ( .D(
        new_AGEMA_signal_4787), .CK(clk), .Q(new_AGEMA_signal_4788) );
  DFF_X1 new_AGEMA_reg_buffer_2904_s_current_state_reg ( .D(
        new_AGEMA_signal_4791), .CK(clk), .Q(new_AGEMA_signal_4792) );
  DFF_X1 new_AGEMA_reg_buffer_2908_s_current_state_reg ( .D(
        new_AGEMA_signal_4795), .CK(clk), .Q(new_AGEMA_signal_4796) );
  DFF_X1 new_AGEMA_reg_buffer_2912_s_current_state_reg ( .D(
        new_AGEMA_signal_4799), .CK(clk), .Q(new_AGEMA_signal_4800) );
  DFF_X1 new_AGEMA_reg_buffer_2916_s_current_state_reg ( .D(
        new_AGEMA_signal_4803), .CK(clk), .Q(new_AGEMA_signal_4804) );
  DFF_X1 new_AGEMA_reg_buffer_2920_s_current_state_reg ( .D(
        new_AGEMA_signal_4807), .CK(clk), .Q(new_AGEMA_signal_4808) );
  DFF_X1 new_AGEMA_reg_buffer_2924_s_current_state_reg ( .D(
        new_AGEMA_signal_4811), .CK(clk), .Q(new_AGEMA_signal_4812) );
  DFF_X1 new_AGEMA_reg_buffer_2928_s_current_state_reg ( .D(
        new_AGEMA_signal_4815), .CK(clk), .Q(new_AGEMA_signal_4816) );
  DFF_X1 new_AGEMA_reg_buffer_2932_s_current_state_reg ( .D(
        new_AGEMA_signal_4819), .CK(clk), .Q(new_AGEMA_signal_4820) );
  DFF_X1 new_AGEMA_reg_buffer_2936_s_current_state_reg ( .D(
        new_AGEMA_signal_4823), .CK(clk), .Q(new_AGEMA_signal_4824) );
  DFF_X1 new_AGEMA_reg_buffer_2940_s_current_state_reg ( .D(
        new_AGEMA_signal_4827), .CK(clk), .Q(new_AGEMA_signal_4828) );
  DFF_X1 new_AGEMA_reg_buffer_2944_s_current_state_reg ( .D(
        new_AGEMA_signal_4831), .CK(clk), .Q(new_AGEMA_signal_4832) );
  DFF_X1 new_AGEMA_reg_buffer_2948_s_current_state_reg ( .D(
        new_AGEMA_signal_4835), .CK(clk), .Q(new_AGEMA_signal_4836) );
  DFF_X1 new_AGEMA_reg_buffer_2952_s_current_state_reg ( .D(
        new_AGEMA_signal_4839), .CK(clk), .Q(new_AGEMA_signal_4840) );
  DFF_X1 new_AGEMA_reg_buffer_2956_s_current_state_reg ( .D(
        new_AGEMA_signal_4843), .CK(clk), .Q(new_AGEMA_signal_4844) );
  DFF_X1 new_AGEMA_reg_buffer_2960_s_current_state_reg ( .D(
        new_AGEMA_signal_4847), .CK(clk), .Q(new_AGEMA_signal_4848) );
  DFF_X1 new_AGEMA_reg_buffer_2964_s_current_state_reg ( .D(
        new_AGEMA_signal_4851), .CK(clk), .Q(new_AGEMA_signal_4852) );
  DFF_X1 new_AGEMA_reg_buffer_2968_s_current_state_reg ( .D(
        new_AGEMA_signal_4855), .CK(clk), .Q(new_AGEMA_signal_4856) );
  DFF_X1 new_AGEMA_reg_buffer_2972_s_current_state_reg ( .D(
        new_AGEMA_signal_4859), .CK(clk), .Q(new_AGEMA_signal_4860) );
  DFF_X1 new_AGEMA_reg_buffer_2976_s_current_state_reg ( .D(
        new_AGEMA_signal_4863), .CK(clk), .Q(new_AGEMA_signal_4864) );
  DFF_X1 new_AGEMA_reg_buffer_2980_s_current_state_reg ( .D(
        new_AGEMA_signal_4867), .CK(clk), .Q(new_AGEMA_signal_4868) );
  DFF_X1 new_AGEMA_reg_buffer_2984_s_current_state_reg ( .D(
        new_AGEMA_signal_4871), .CK(clk), .Q(new_AGEMA_signal_4872) );
  DFF_X1 new_AGEMA_reg_buffer_2988_s_current_state_reg ( .D(
        new_AGEMA_signal_4875), .CK(clk), .Q(new_AGEMA_signal_4876) );
  DFF_X1 new_AGEMA_reg_buffer_2992_s_current_state_reg ( .D(
        new_AGEMA_signal_4879), .CK(clk), .Q(new_AGEMA_signal_4880) );
  DFF_X1 new_AGEMA_reg_buffer_2996_s_current_state_reg ( .D(
        new_AGEMA_signal_4883), .CK(clk), .Q(new_AGEMA_signal_4884) );
  DFF_X1 new_AGEMA_reg_buffer_3000_s_current_state_reg ( .D(
        new_AGEMA_signal_4887), .CK(clk), .Q(new_AGEMA_signal_4888) );
  DFF_X1 new_AGEMA_reg_buffer_3004_s_current_state_reg ( .D(
        new_AGEMA_signal_4891), .CK(clk), .Q(new_AGEMA_signal_4892) );
  DFF_X1 new_AGEMA_reg_buffer_3008_s_current_state_reg ( .D(
        new_AGEMA_signal_4895), .CK(clk), .Q(new_AGEMA_signal_4896) );
  DFF_X1 new_AGEMA_reg_buffer_3012_s_current_state_reg ( .D(
        new_AGEMA_signal_4899), .CK(clk), .Q(new_AGEMA_signal_4900) );
  DFF_X1 new_AGEMA_reg_buffer_3016_s_current_state_reg ( .D(
        new_AGEMA_signal_4903), .CK(clk), .Q(new_AGEMA_signal_4904) );
  DFF_X1 new_AGEMA_reg_buffer_3020_s_current_state_reg ( .D(
        new_AGEMA_signal_4907), .CK(clk), .Q(new_AGEMA_signal_4908) );
  DFF_X1 new_AGEMA_reg_buffer_3024_s_current_state_reg ( .D(
        new_AGEMA_signal_4911), .CK(clk), .Q(new_AGEMA_signal_4912) );
  DFF_X1 new_AGEMA_reg_buffer_3028_s_current_state_reg ( .D(
        new_AGEMA_signal_4915), .CK(clk), .Q(new_AGEMA_signal_4916) );
  DFF_X1 new_AGEMA_reg_buffer_3032_s_current_state_reg ( .D(
        new_AGEMA_signal_4919), .CK(clk), .Q(new_AGEMA_signal_4920) );
  DFF_X1 new_AGEMA_reg_buffer_3036_s_current_state_reg ( .D(
        new_AGEMA_signal_4923), .CK(clk), .Q(new_AGEMA_signal_4924) );
  DFF_X1 new_AGEMA_reg_buffer_3040_s_current_state_reg ( .D(
        new_AGEMA_signal_4927), .CK(clk), .Q(new_AGEMA_signal_4928) );
  DFF_X1 new_AGEMA_reg_buffer_3044_s_current_state_reg ( .D(
        new_AGEMA_signal_4931), .CK(clk), .Q(new_AGEMA_signal_4932) );
  DFF_X1 new_AGEMA_reg_buffer_3048_s_current_state_reg ( .D(
        new_AGEMA_signal_4935), .CK(clk), .Q(new_AGEMA_signal_4936) );
  DFF_X1 new_AGEMA_reg_buffer_3052_s_current_state_reg ( .D(
        new_AGEMA_signal_4939), .CK(clk), .Q(new_AGEMA_signal_4940) );
  DFF_X1 new_AGEMA_reg_buffer_3056_s_current_state_reg ( .D(
        new_AGEMA_signal_4943), .CK(clk), .Q(new_AGEMA_signal_4944) );
  DFF_X1 new_AGEMA_reg_buffer_3060_s_current_state_reg ( .D(
        new_AGEMA_signal_4947), .CK(clk), .Q(new_AGEMA_signal_4948) );
  DFF_X1 new_AGEMA_reg_buffer_3064_s_current_state_reg ( .D(
        new_AGEMA_signal_4951), .CK(clk), .Q(new_AGEMA_signal_4952) );
  DFF_X1 new_AGEMA_reg_buffer_3068_s_current_state_reg ( .D(
        new_AGEMA_signal_4955), .CK(clk), .Q(new_AGEMA_signal_4956) );
  DFF_X1 new_AGEMA_reg_buffer_3072_s_current_state_reg ( .D(
        new_AGEMA_signal_4959), .CK(clk), .Q(new_AGEMA_signal_4960) );
  DFF_X1 new_AGEMA_reg_buffer_3076_s_current_state_reg ( .D(
        new_AGEMA_signal_4963), .CK(clk), .Q(new_AGEMA_signal_4964) );
  DFF_X1 new_AGEMA_reg_buffer_3080_s_current_state_reg ( .D(
        new_AGEMA_signal_4967), .CK(clk), .Q(new_AGEMA_signal_4968) );
  DFF_X1 new_AGEMA_reg_buffer_3084_s_current_state_reg ( .D(
        new_AGEMA_signal_4971), .CK(clk), .Q(new_AGEMA_signal_4972) );
  DFF_X1 new_AGEMA_reg_buffer_3088_s_current_state_reg ( .D(
        new_AGEMA_signal_4975), .CK(clk), .Q(new_AGEMA_signal_4976) );
  DFF_X1 new_AGEMA_reg_buffer_3092_s_current_state_reg ( .D(
        new_AGEMA_signal_4979), .CK(clk), .Q(new_AGEMA_signal_4980) );
  DFF_X1 new_AGEMA_reg_buffer_3096_s_current_state_reg ( .D(
        new_AGEMA_signal_4983), .CK(clk), .Q(new_AGEMA_signal_4984) );
  DFF_X1 new_AGEMA_reg_buffer_3100_s_current_state_reg ( .D(
        new_AGEMA_signal_4987), .CK(clk), .Q(new_AGEMA_signal_4988) );
  DFF_X1 new_AGEMA_reg_buffer_3104_s_current_state_reg ( .D(
        new_AGEMA_signal_4991), .CK(clk), .Q(new_AGEMA_signal_4992) );
  DFF_X1 new_AGEMA_reg_buffer_3108_s_current_state_reg ( .D(
        new_AGEMA_signal_4995), .CK(clk), .Q(new_AGEMA_signal_4996) );
  DFF_X1 new_AGEMA_reg_buffer_3112_s_current_state_reg ( .D(
        new_AGEMA_signal_4999), .CK(clk), .Q(new_AGEMA_signal_5000) );
  DFF_X1 new_AGEMA_reg_buffer_3116_s_current_state_reg ( .D(
        new_AGEMA_signal_5003), .CK(clk), .Q(new_AGEMA_signal_5004) );
  DFF_X1 new_AGEMA_reg_buffer_3120_s_current_state_reg ( .D(
        new_AGEMA_signal_5007), .CK(clk), .Q(new_AGEMA_signal_5008) );
  DFF_X1 new_AGEMA_reg_buffer_3124_s_current_state_reg ( .D(
        new_AGEMA_signal_5011), .CK(clk), .Q(new_AGEMA_signal_5012) );
  DFF_X1 new_AGEMA_reg_buffer_3128_s_current_state_reg ( .D(
        new_AGEMA_signal_5015), .CK(clk), .Q(new_AGEMA_signal_5016) );
  DFF_X1 new_AGEMA_reg_buffer_3132_s_current_state_reg ( .D(
        new_AGEMA_signal_5019), .CK(clk), .Q(new_AGEMA_signal_5020) );
  DFF_X1 new_AGEMA_reg_buffer_3136_s_current_state_reg ( .D(
        new_AGEMA_signal_5023), .CK(clk), .Q(new_AGEMA_signal_5024) );
  DFF_X1 new_AGEMA_reg_buffer_3140_s_current_state_reg ( .D(
        new_AGEMA_signal_5027), .CK(clk), .Q(new_AGEMA_signal_5028) );
  DFF_X1 new_AGEMA_reg_buffer_3144_s_current_state_reg ( .D(
        new_AGEMA_signal_5031), .CK(clk), .Q(new_AGEMA_signal_5032) );
  DFF_X1 new_AGEMA_reg_buffer_3148_s_current_state_reg ( .D(
        new_AGEMA_signal_5035), .CK(clk), .Q(new_AGEMA_signal_5036) );
  DFF_X1 new_AGEMA_reg_buffer_3152_s_current_state_reg ( .D(
        new_AGEMA_signal_5039), .CK(clk), .Q(new_AGEMA_signal_5040) );
  DFF_X1 new_AGEMA_reg_buffer_3156_s_current_state_reg ( .D(
        new_AGEMA_signal_5043), .CK(clk), .Q(new_AGEMA_signal_5044) );
  DFF_X1 new_AGEMA_reg_buffer_3160_s_current_state_reg ( .D(
        new_AGEMA_signal_5047), .CK(clk), .Q(new_AGEMA_signal_5048) );
  DFF_X1 new_AGEMA_reg_buffer_3164_s_current_state_reg ( .D(
        new_AGEMA_signal_5051), .CK(clk), .Q(new_AGEMA_signal_5052) );
  DFF_X1 new_AGEMA_reg_buffer_3168_s_current_state_reg ( .D(
        new_AGEMA_signal_5055), .CK(clk), .Q(new_AGEMA_signal_5056) );
  DFF_X1 new_AGEMA_reg_buffer_3172_s_current_state_reg ( .D(
        new_AGEMA_signal_5059), .CK(clk), .Q(new_AGEMA_signal_5060) );
  DFF_X1 new_AGEMA_reg_buffer_3176_s_current_state_reg ( .D(
        new_AGEMA_signal_5063), .CK(clk), .Q(new_AGEMA_signal_5064) );
  DFF_X1 new_AGEMA_reg_buffer_3180_s_current_state_reg ( .D(
        new_AGEMA_signal_5067), .CK(clk), .Q(new_AGEMA_signal_5068) );
  DFF_X1 new_AGEMA_reg_buffer_3184_s_current_state_reg ( .D(
        new_AGEMA_signal_5071), .CK(clk), .Q(new_AGEMA_signal_5072) );
  DFF_X1 new_AGEMA_reg_buffer_3188_s_current_state_reg ( .D(
        new_AGEMA_signal_5075), .CK(clk), .Q(new_AGEMA_signal_5076) );
  DFF_X1 new_AGEMA_reg_buffer_3192_s_current_state_reg ( .D(
        new_AGEMA_signal_5079), .CK(clk), .Q(new_AGEMA_signal_5080) );
  DFF_X1 new_AGEMA_reg_buffer_3196_s_current_state_reg ( .D(
        new_AGEMA_signal_5083), .CK(clk), .Q(new_AGEMA_signal_5084) );
  DFF_X1 new_AGEMA_reg_buffer_3200_s_current_state_reg ( .D(
        new_AGEMA_signal_5087), .CK(clk), .Q(new_AGEMA_signal_5088) );
  DFF_X1 new_AGEMA_reg_buffer_3204_s_current_state_reg ( .D(
        new_AGEMA_signal_5091), .CK(clk), .Q(new_AGEMA_signal_5092) );
  DFF_X1 new_AGEMA_reg_buffer_3208_s_current_state_reg ( .D(
        new_AGEMA_signal_5095), .CK(clk), .Q(new_AGEMA_signal_5096) );
  DFF_X1 new_AGEMA_reg_buffer_3212_s_current_state_reg ( .D(
        new_AGEMA_signal_5099), .CK(clk), .Q(new_AGEMA_signal_5100) );
  DFF_X1 new_AGEMA_reg_buffer_3216_s_current_state_reg ( .D(
        new_AGEMA_signal_5103), .CK(clk), .Q(new_AGEMA_signal_5104) );
  DFF_X1 new_AGEMA_reg_buffer_3220_s_current_state_reg ( .D(
        new_AGEMA_signal_5107), .CK(clk), .Q(new_AGEMA_signal_5108) );
  DFF_X1 new_AGEMA_reg_buffer_3224_s_current_state_reg ( .D(
        new_AGEMA_signal_5111), .CK(clk), .Q(new_AGEMA_signal_5112) );
  DFF_X1 new_AGEMA_reg_buffer_3228_s_current_state_reg ( .D(
        new_AGEMA_signal_5115), .CK(clk), .Q(new_AGEMA_signal_5116) );
  DFF_X1 new_AGEMA_reg_buffer_3232_s_current_state_reg ( .D(
        new_AGEMA_signal_5119), .CK(clk), .Q(new_AGEMA_signal_5120) );
  DFF_X1 new_AGEMA_reg_buffer_3236_s_current_state_reg ( .D(
        new_AGEMA_signal_5123), .CK(clk), .Q(new_AGEMA_signal_5124) );
  DFF_X1 new_AGEMA_reg_buffer_3240_s_current_state_reg ( .D(
        new_AGEMA_signal_5127), .CK(clk), .Q(new_AGEMA_signal_5128) );
  DFF_X1 new_AGEMA_reg_buffer_3244_s_current_state_reg ( .D(
        new_AGEMA_signal_5131), .CK(clk), .Q(new_AGEMA_signal_5132) );
  DFF_X1 new_AGEMA_reg_buffer_3248_s_current_state_reg ( .D(
        new_AGEMA_signal_5135), .CK(clk), .Q(new_AGEMA_signal_5136) );
  DFF_X1 new_AGEMA_reg_buffer_3252_s_current_state_reg ( .D(
        new_AGEMA_signal_5139), .CK(clk), .Q(new_AGEMA_signal_5140) );
  DFF_X1 new_AGEMA_reg_buffer_3256_s_current_state_reg ( .D(
        new_AGEMA_signal_5143), .CK(clk), .Q(new_AGEMA_signal_5144) );
  DFF_X1 new_AGEMA_reg_buffer_3260_s_current_state_reg ( .D(
        new_AGEMA_signal_5147), .CK(clk), .Q(new_AGEMA_signal_5148) );
  DFF_X1 new_AGEMA_reg_buffer_3264_s_current_state_reg ( .D(
        new_AGEMA_signal_5151), .CK(clk), .Q(new_AGEMA_signal_5152) );
  DFF_X1 new_AGEMA_reg_buffer_3268_s_current_state_reg ( .D(
        new_AGEMA_signal_5155), .CK(clk), .Q(new_AGEMA_signal_5156) );
  DFF_X1 new_AGEMA_reg_buffer_3272_s_current_state_reg ( .D(
        new_AGEMA_signal_5159), .CK(clk), .Q(new_AGEMA_signal_5160) );
  DFF_X1 new_AGEMA_reg_buffer_3276_s_current_state_reg ( .D(
        new_AGEMA_signal_5163), .CK(clk), .Q(new_AGEMA_signal_5164) );
  DFF_X1 new_AGEMA_reg_buffer_3280_s_current_state_reg ( .D(
        new_AGEMA_signal_5167), .CK(clk), .Q(new_AGEMA_signal_5168) );
  DFF_X1 new_AGEMA_reg_buffer_3284_s_current_state_reg ( .D(
        new_AGEMA_signal_5171), .CK(clk), .Q(new_AGEMA_signal_5172) );
  DFF_X1 new_AGEMA_reg_buffer_3288_s_current_state_reg ( .D(
        new_AGEMA_signal_5175), .CK(clk), .Q(new_AGEMA_signal_5176) );
  DFF_X1 new_AGEMA_reg_buffer_3292_s_current_state_reg ( .D(
        new_AGEMA_signal_5179), .CK(clk), .Q(new_AGEMA_signal_5180) );
  DFF_X1 new_AGEMA_reg_buffer_3296_s_current_state_reg ( .D(
        new_AGEMA_signal_5183), .CK(clk), .Q(new_AGEMA_signal_5184) );
  DFF_X1 new_AGEMA_reg_buffer_3300_s_current_state_reg ( .D(
        new_AGEMA_signal_5187), .CK(clk), .Q(new_AGEMA_signal_5188) );
  DFF_X1 new_AGEMA_reg_buffer_3304_s_current_state_reg ( .D(
        new_AGEMA_signal_5191), .CK(clk), .Q(new_AGEMA_signal_5192) );
  DFF_X1 new_AGEMA_reg_buffer_3308_s_current_state_reg ( .D(
        new_AGEMA_signal_5195), .CK(clk), .Q(new_AGEMA_signal_5196) );
  DFF_X1 new_AGEMA_reg_buffer_3312_s_current_state_reg ( .D(
        new_AGEMA_signal_5199), .CK(clk), .Q(new_AGEMA_signal_5200) );
  DFF_X1 new_AGEMA_reg_buffer_3316_s_current_state_reg ( .D(
        new_AGEMA_signal_5203), .CK(clk), .Q(new_AGEMA_signal_5204) );
  DFF_X1 new_AGEMA_reg_buffer_3320_s_current_state_reg ( .D(
        new_AGEMA_signal_5207), .CK(clk), .Q(new_AGEMA_signal_5208) );
  DFF_X1 new_AGEMA_reg_buffer_3324_s_current_state_reg ( .D(
        new_AGEMA_signal_5211), .CK(clk), .Q(new_AGEMA_signal_5212) );
  DFF_X1 new_AGEMA_reg_buffer_3328_s_current_state_reg ( .D(
        new_AGEMA_signal_5215), .CK(clk), .Q(new_AGEMA_signal_5216) );
  DFF_X1 new_AGEMA_reg_buffer_3332_s_current_state_reg ( .D(
        new_AGEMA_signal_5219), .CK(clk), .Q(new_AGEMA_signal_5220) );
  DFF_X1 new_AGEMA_reg_buffer_3336_s_current_state_reg ( .D(
        new_AGEMA_signal_5223), .CK(clk), .Q(new_AGEMA_signal_5224) );
  DFF_X1 new_AGEMA_reg_buffer_3340_s_current_state_reg ( .D(
        new_AGEMA_signal_5227), .CK(clk), .Q(new_AGEMA_signal_5228) );
  DFF_X1 new_AGEMA_reg_buffer_3344_s_current_state_reg ( .D(
        new_AGEMA_signal_5231), .CK(clk), .Q(new_AGEMA_signal_5232) );
  DFF_X1 new_AGEMA_reg_buffer_3348_s_current_state_reg ( .D(
        new_AGEMA_signal_5235), .CK(clk), .Q(new_AGEMA_signal_5236) );
  DFF_X1 new_AGEMA_reg_buffer_3352_s_current_state_reg ( .D(
        new_AGEMA_signal_5239), .CK(clk), .Q(new_AGEMA_signal_5240) );
  DFF_X1 new_AGEMA_reg_buffer_3356_s_current_state_reg ( .D(
        new_AGEMA_signal_5243), .CK(clk), .Q(new_AGEMA_signal_5244) );
  DFF_X1 new_AGEMA_reg_buffer_3360_s_current_state_reg ( .D(
        new_AGEMA_signal_5247), .CK(clk), .Q(new_AGEMA_signal_5248) );
  DFF_X1 new_AGEMA_reg_buffer_3364_s_current_state_reg ( .D(
        new_AGEMA_signal_5251), .CK(clk), .Q(new_AGEMA_signal_5252) );
  DFF_X1 new_AGEMA_reg_buffer_3368_s_current_state_reg ( .D(
        new_AGEMA_signal_5255), .CK(clk), .Q(new_AGEMA_signal_5256) );
  DFF_X1 new_AGEMA_reg_buffer_3372_s_current_state_reg ( .D(
        new_AGEMA_signal_5259), .CK(clk), .Q(new_AGEMA_signal_5260) );
  DFF_X1 new_AGEMA_reg_buffer_3376_s_current_state_reg ( .D(
        new_AGEMA_signal_5263), .CK(clk), .Q(new_AGEMA_signal_5264) );
  DFF_X1 new_AGEMA_reg_buffer_3380_s_current_state_reg ( .D(
        new_AGEMA_signal_5267), .CK(clk), .Q(new_AGEMA_signal_5268) );
  DFF_X1 new_AGEMA_reg_buffer_3384_s_current_state_reg ( .D(
        new_AGEMA_signal_5271), .CK(clk), .Q(new_AGEMA_signal_5272) );
  DFF_X1 new_AGEMA_reg_buffer_3388_s_current_state_reg ( .D(
        new_AGEMA_signal_5275), .CK(clk), .Q(new_AGEMA_signal_5276) );
  DFF_X1 new_AGEMA_reg_buffer_3392_s_current_state_reg ( .D(
        new_AGEMA_signal_5279), .CK(clk), .Q(new_AGEMA_signal_5280) );
  DFF_X1 new_AGEMA_reg_buffer_3396_s_current_state_reg ( .D(
        new_AGEMA_signal_5283), .CK(clk), .Q(new_AGEMA_signal_5284) );
  DFF_X1 new_AGEMA_reg_buffer_3400_s_current_state_reg ( .D(
        new_AGEMA_signal_5287), .CK(clk), .Q(new_AGEMA_signal_5288) );
  DFF_X1 new_AGEMA_reg_buffer_3404_s_current_state_reg ( .D(
        new_AGEMA_signal_5291), .CK(clk), .Q(new_AGEMA_signal_5292) );
  DFF_X1 new_AGEMA_reg_buffer_3408_s_current_state_reg ( .D(
        new_AGEMA_signal_5295), .CK(clk), .Q(new_AGEMA_signal_5296) );
  DFF_X1 new_AGEMA_reg_buffer_3412_s_current_state_reg ( .D(
        new_AGEMA_signal_5299), .CK(clk), .Q(new_AGEMA_signal_5300) );
  DFF_X1 new_AGEMA_reg_buffer_3416_s_current_state_reg ( .D(
        new_AGEMA_signal_5303), .CK(clk), .Q(new_AGEMA_signal_5304) );
  DFF_X1 new_AGEMA_reg_buffer_3420_s_current_state_reg ( .D(
        new_AGEMA_signal_5307), .CK(clk), .Q(new_AGEMA_signal_5308) );
  DFF_X1 new_AGEMA_reg_buffer_3424_s_current_state_reg ( .D(
        new_AGEMA_signal_5311), .CK(clk), .Q(new_AGEMA_signal_5312) );
  DFF_X1 new_AGEMA_reg_buffer_3428_s_current_state_reg ( .D(
        new_AGEMA_signal_5315), .CK(clk), .Q(new_AGEMA_signal_5316) );
  DFF_X1 new_AGEMA_reg_buffer_3432_s_current_state_reg ( .D(
        new_AGEMA_signal_5319), .CK(clk), .Q(new_AGEMA_signal_5320) );
  DFF_X1 new_AGEMA_reg_buffer_3436_s_current_state_reg ( .D(
        new_AGEMA_signal_5323), .CK(clk), .Q(new_AGEMA_signal_5324) );
  DFF_X1 new_AGEMA_reg_buffer_3440_s_current_state_reg ( .D(
        new_AGEMA_signal_5327), .CK(clk), .Q(new_AGEMA_signal_5328) );
  DFF_X1 new_AGEMA_reg_buffer_3444_s_current_state_reg ( .D(
        new_AGEMA_signal_5331), .CK(clk), .Q(new_AGEMA_signal_5332) );
  DFF_X1 new_AGEMA_reg_buffer_3448_s_current_state_reg ( .D(
        new_AGEMA_signal_5335), .CK(clk), .Q(new_AGEMA_signal_5336) );
  DFF_X1 new_AGEMA_reg_buffer_3452_s_current_state_reg ( .D(
        new_AGEMA_signal_5339), .CK(clk), .Q(new_AGEMA_signal_5340) );
  DFF_X1 new_AGEMA_reg_buffer_3456_s_current_state_reg ( .D(
        new_AGEMA_signal_5343), .CK(clk), .Q(new_AGEMA_signal_5344) );
  DFF_X1 new_AGEMA_reg_buffer_3460_s_current_state_reg ( .D(
        new_AGEMA_signal_5347), .CK(clk), .Q(new_AGEMA_signal_5348) );
  DFF_X1 new_AGEMA_reg_buffer_3464_s_current_state_reg ( .D(
        new_AGEMA_signal_5351), .CK(clk), .Q(new_AGEMA_signal_5352) );
  DFF_X1 new_AGEMA_reg_buffer_3468_s_current_state_reg ( .D(
        new_AGEMA_signal_5355), .CK(clk), .Q(new_AGEMA_signal_5356) );
  DFF_X1 new_AGEMA_reg_buffer_3472_s_current_state_reg ( .D(
        new_AGEMA_signal_5359), .CK(clk), .Q(new_AGEMA_signal_5360) );
  DFF_X1 new_AGEMA_reg_buffer_3476_s_current_state_reg ( .D(
        new_AGEMA_signal_5363), .CK(clk), .Q(new_AGEMA_signal_5364) );
  DFF_X1 new_AGEMA_reg_buffer_3480_s_current_state_reg ( .D(
        new_AGEMA_signal_5367), .CK(clk), .Q(new_AGEMA_signal_5368) );
  DFF_X1 new_AGEMA_reg_buffer_3484_s_current_state_reg ( .D(
        new_AGEMA_signal_5371), .CK(clk), .Q(new_AGEMA_signal_5372) );
  DFF_X1 new_AGEMA_reg_buffer_3488_s_current_state_reg ( .D(
        new_AGEMA_signal_5375), .CK(clk), .Q(new_AGEMA_signal_5376) );
  DFF_X1 new_AGEMA_reg_buffer_3492_s_current_state_reg ( .D(
        new_AGEMA_signal_5379), .CK(clk), .Q(new_AGEMA_signal_5380) );
  DFF_X1 new_AGEMA_reg_buffer_3496_s_current_state_reg ( .D(
        new_AGEMA_signal_5383), .CK(clk), .Q(new_AGEMA_signal_5384) );
  DFF_X1 new_AGEMA_reg_buffer_3500_s_current_state_reg ( .D(
        new_AGEMA_signal_5387), .CK(clk), .Q(new_AGEMA_signal_5388) );
  DFF_X1 new_AGEMA_reg_buffer_3504_s_current_state_reg ( .D(
        new_AGEMA_signal_5391), .CK(clk), .Q(new_AGEMA_signal_5392) );
  DFF_X1 new_AGEMA_reg_buffer_3508_s_current_state_reg ( .D(
        new_AGEMA_signal_5395), .CK(clk), .Q(new_AGEMA_signal_5396) );
  DFF_X1 new_AGEMA_reg_buffer_3512_s_current_state_reg ( .D(
        new_AGEMA_signal_5399), .CK(clk), .Q(new_AGEMA_signal_5400) );
  DFF_X1 new_AGEMA_reg_buffer_3516_s_current_state_reg ( .D(
        new_AGEMA_signal_5403), .CK(clk), .Q(new_AGEMA_signal_5404) );
  DFF_X1 new_AGEMA_reg_buffer_3520_s_current_state_reg ( .D(
        new_AGEMA_signal_5407), .CK(clk), .Q(new_AGEMA_signal_5408) );
  DFF_X1 new_AGEMA_reg_buffer_3524_s_current_state_reg ( .D(
        new_AGEMA_signal_5411), .CK(clk), .Q(new_AGEMA_signal_5412) );
  DFF_X1 new_AGEMA_reg_buffer_3528_s_current_state_reg ( .D(
        new_AGEMA_signal_5415), .CK(clk), .Q(new_AGEMA_signal_5416) );
  DFF_X1 new_AGEMA_reg_buffer_3532_s_current_state_reg ( .D(
        new_AGEMA_signal_5419), .CK(clk), .Q(new_AGEMA_signal_5420) );
  DFF_X1 new_AGEMA_reg_buffer_3536_s_current_state_reg ( .D(
        new_AGEMA_signal_5423), .CK(clk), .Q(new_AGEMA_signal_5424) );
  DFF_X1 new_AGEMA_reg_buffer_3540_s_current_state_reg ( .D(
        new_AGEMA_signal_5427), .CK(clk), .Q(new_AGEMA_signal_5428) );
  DFF_X1 new_AGEMA_reg_buffer_3544_s_current_state_reg ( .D(
        new_AGEMA_signal_5431), .CK(clk), .Q(new_AGEMA_signal_5432) );
  DFF_X1 new_AGEMA_reg_buffer_3548_s_current_state_reg ( .D(
        new_AGEMA_signal_5435), .CK(clk), .Q(new_AGEMA_signal_5436) );
  DFF_X1 new_AGEMA_reg_buffer_3552_s_current_state_reg ( .D(
        new_AGEMA_signal_5439), .CK(clk), .Q(new_AGEMA_signal_5440) );
  DFF_X1 new_AGEMA_reg_buffer_3556_s_current_state_reg ( .D(
        new_AGEMA_signal_5443), .CK(clk), .Q(new_AGEMA_signal_5444) );
  DFF_X1 new_AGEMA_reg_buffer_3560_s_current_state_reg ( .D(
        new_AGEMA_signal_5447), .CK(clk), .Q(new_AGEMA_signal_5448) );
  DFF_X1 new_AGEMA_reg_buffer_3564_s_current_state_reg ( .D(
        new_AGEMA_signal_5451), .CK(clk), .Q(new_AGEMA_signal_5452) );
  DFF_X1 new_AGEMA_reg_buffer_3568_s_current_state_reg ( .D(
        new_AGEMA_signal_5455), .CK(clk), .Q(new_AGEMA_signal_5456) );
  DFF_X1 new_AGEMA_reg_buffer_3572_s_current_state_reg ( .D(
        new_AGEMA_signal_5459), .CK(clk), .Q(new_AGEMA_signal_5460) );
  DFF_X1 new_AGEMA_reg_buffer_3576_s_current_state_reg ( .D(
        new_AGEMA_signal_5463), .CK(clk), .Q(new_AGEMA_signal_5464) );
  DFF_X1 new_AGEMA_reg_buffer_3580_s_current_state_reg ( .D(
        new_AGEMA_signal_5467), .CK(clk), .Q(new_AGEMA_signal_5468) );
  DFF_X1 new_AGEMA_reg_buffer_3584_s_current_state_reg ( .D(
        new_AGEMA_signal_5471), .CK(clk), .Q(new_AGEMA_signal_5472) );
  DFF_X1 new_AGEMA_reg_buffer_3588_s_current_state_reg ( .D(
        new_AGEMA_signal_5475), .CK(clk), .Q(new_AGEMA_signal_5476) );
  DFF_X1 new_AGEMA_reg_buffer_3592_s_current_state_reg ( .D(
        new_AGEMA_signal_5479), .CK(clk), .Q(new_AGEMA_signal_5480) );
  DFF_X1 new_AGEMA_reg_buffer_3596_s_current_state_reg ( .D(
        new_AGEMA_signal_5483), .CK(clk), .Q(new_AGEMA_signal_5484) );
  DFF_X1 new_AGEMA_reg_buffer_3600_s_current_state_reg ( .D(
        new_AGEMA_signal_5487), .CK(clk), .Q(new_AGEMA_signal_5488) );
  DFF_X1 new_AGEMA_reg_buffer_3604_s_current_state_reg ( .D(
        new_AGEMA_signal_5491), .CK(clk), .Q(new_AGEMA_signal_5492) );
  DFF_X1 new_AGEMA_reg_buffer_3608_s_current_state_reg ( .D(
        new_AGEMA_signal_5495), .CK(clk), .Q(new_AGEMA_signal_5496) );
  DFF_X1 new_AGEMA_reg_buffer_3612_s_current_state_reg ( .D(
        new_AGEMA_signal_5499), .CK(clk), .Q(new_AGEMA_signal_5500) );
  DFF_X1 new_AGEMA_reg_buffer_3616_s_current_state_reg ( .D(
        new_AGEMA_signal_5503), .CK(clk), .Q(new_AGEMA_signal_5504) );
  DFF_X1 new_AGEMA_reg_buffer_3620_s_current_state_reg ( .D(
        new_AGEMA_signal_5507), .CK(clk), .Q(new_AGEMA_signal_5508) );
  DFF_X1 new_AGEMA_reg_buffer_3624_s_current_state_reg ( .D(
        new_AGEMA_signal_5511), .CK(clk), .Q(new_AGEMA_signal_5512) );
  DFF_X1 new_AGEMA_reg_buffer_3628_s_current_state_reg ( .D(
        new_AGEMA_signal_5515), .CK(clk), .Q(new_AGEMA_signal_5516) );
  DFF_X1 new_AGEMA_reg_buffer_3632_s_current_state_reg ( .D(
        new_AGEMA_signal_5519), .CK(clk), .Q(new_AGEMA_signal_5520) );
  DFF_X1 new_AGEMA_reg_buffer_3636_s_current_state_reg ( .D(
        new_AGEMA_signal_5523), .CK(clk), .Q(new_AGEMA_signal_5524) );
  DFF_X1 new_AGEMA_reg_buffer_3640_s_current_state_reg ( .D(
        new_AGEMA_signal_5527), .CK(clk), .Q(new_AGEMA_signal_5528) );
  DFF_X1 new_AGEMA_reg_buffer_3644_s_current_state_reg ( .D(
        new_AGEMA_signal_5531), .CK(clk), .Q(new_AGEMA_signal_5532) );
  DFF_X1 new_AGEMA_reg_buffer_3648_s_current_state_reg ( .D(
        new_AGEMA_signal_5535), .CK(clk), .Q(new_AGEMA_signal_5536) );
  DFF_X1 new_AGEMA_reg_buffer_3652_s_current_state_reg ( .D(
        new_AGEMA_signal_5539), .CK(clk), .Q(new_AGEMA_signal_5540) );
  DFF_X1 new_AGEMA_reg_buffer_3656_s_current_state_reg ( .D(
        new_AGEMA_signal_5543), .CK(clk), .Q(new_AGEMA_signal_5544) );
  DFF_X1 new_AGEMA_reg_buffer_3660_s_current_state_reg ( .D(
        new_AGEMA_signal_5547), .CK(clk), .Q(new_AGEMA_signal_5548) );
  DFF_X1 new_AGEMA_reg_buffer_3664_s_current_state_reg ( .D(
        new_AGEMA_signal_5551), .CK(clk), .Q(new_AGEMA_signal_5552) );
  DFF_X1 new_AGEMA_reg_buffer_3668_s_current_state_reg ( .D(
        new_AGEMA_signal_5555), .CK(clk), .Q(new_AGEMA_signal_5556) );
  DFF_X1 new_AGEMA_reg_buffer_3672_s_current_state_reg ( .D(
        new_AGEMA_signal_5559), .CK(clk), .Q(new_AGEMA_signal_5560) );
  DFF_X1 new_AGEMA_reg_buffer_3676_s_current_state_reg ( .D(
        new_AGEMA_signal_5563), .CK(clk), .Q(new_AGEMA_signal_5564) );
  DFF_X1 new_AGEMA_reg_buffer_3680_s_current_state_reg ( .D(
        new_AGEMA_signal_5567), .CK(clk), .Q(new_AGEMA_signal_5568) );
  DFF_X1 new_AGEMA_reg_buffer_3684_s_current_state_reg ( .D(
        new_AGEMA_signal_5571), .CK(clk), .Q(new_AGEMA_signal_5572) );
  DFF_X1 new_AGEMA_reg_buffer_3688_s_current_state_reg ( .D(
        new_AGEMA_signal_5575), .CK(clk), .Q(new_AGEMA_signal_5576) );
  DFF_X1 new_AGEMA_reg_buffer_3692_s_current_state_reg ( .D(
        new_AGEMA_signal_5579), .CK(clk), .Q(new_AGEMA_signal_5580) );
  DFF_X1 new_AGEMA_reg_buffer_3696_s_current_state_reg ( .D(
        new_AGEMA_signal_5583), .CK(clk), .Q(new_AGEMA_signal_5584) );
  DFF_X1 new_AGEMA_reg_buffer_3700_s_current_state_reg ( .D(
        new_AGEMA_signal_5587), .CK(clk), .Q(new_AGEMA_signal_5588) );
  DFF_X1 new_AGEMA_reg_buffer_3704_s_current_state_reg ( .D(
        new_AGEMA_signal_5591), .CK(clk), .Q(new_AGEMA_signal_5592) );
  DFF_X1 new_AGEMA_reg_buffer_3708_s_current_state_reg ( .D(
        new_AGEMA_signal_5595), .CK(clk), .Q(new_AGEMA_signal_5596) );
  DFF_X1 new_AGEMA_reg_buffer_3712_s_current_state_reg ( .D(
        new_AGEMA_signal_5599), .CK(clk), .Q(new_AGEMA_signal_5600) );
  DFF_X1 new_AGEMA_reg_buffer_3716_s_current_state_reg ( .D(
        new_AGEMA_signal_5603), .CK(clk), .Q(new_AGEMA_signal_5604) );
  DFF_X1 new_AGEMA_reg_buffer_3720_s_current_state_reg ( .D(
        new_AGEMA_signal_5607), .CK(clk), .Q(new_AGEMA_signal_5608) );
  DFF_X1 new_AGEMA_reg_buffer_3724_s_current_state_reg ( .D(
        new_AGEMA_signal_5611), .CK(clk), .Q(new_AGEMA_signal_5612) );
  DFF_X1 new_AGEMA_reg_buffer_3728_s_current_state_reg ( .D(
        new_AGEMA_signal_5615), .CK(clk), .Q(new_AGEMA_signal_5616) );
  DFF_X1 new_AGEMA_reg_buffer_3732_s_current_state_reg ( .D(
        new_AGEMA_signal_5619), .CK(clk), .Q(new_AGEMA_signal_5620) );
  DFF_X1 new_AGEMA_reg_buffer_3736_s_current_state_reg ( .D(
        new_AGEMA_signal_5623), .CK(clk), .Q(new_AGEMA_signal_5624) );
  DFF_X1 new_AGEMA_reg_buffer_3740_s_current_state_reg ( .D(
        new_AGEMA_signal_5627), .CK(clk), .Q(new_AGEMA_signal_5628) );
  DFF_X1 new_AGEMA_reg_buffer_3744_s_current_state_reg ( .D(
        new_AGEMA_signal_5631), .CK(clk), .Q(new_AGEMA_signal_5632) );
  DFF_X1 new_AGEMA_reg_buffer_3748_s_current_state_reg ( .D(
        new_AGEMA_signal_5635), .CK(clk), .Q(new_AGEMA_signal_5636) );
  DFF_X1 new_AGEMA_reg_buffer_3752_s_current_state_reg ( .D(
        new_AGEMA_signal_5639), .CK(clk), .Q(new_AGEMA_signal_5640) );
  DFF_X1 new_AGEMA_reg_buffer_3756_s_current_state_reg ( .D(
        new_AGEMA_signal_5643), .CK(clk), .Q(new_AGEMA_signal_5644) );
  DFF_X1 new_AGEMA_reg_buffer_3760_s_current_state_reg ( .D(
        new_AGEMA_signal_5647), .CK(clk), .Q(new_AGEMA_signal_5648) );
  DFF_X1 new_AGEMA_reg_buffer_3764_s_current_state_reg ( .D(
        new_AGEMA_signal_5651), .CK(clk), .Q(new_AGEMA_signal_5652) );
  DFF_X1 new_AGEMA_reg_buffer_3768_s_current_state_reg ( .D(
        new_AGEMA_signal_5655), .CK(clk), .Q(new_AGEMA_signal_5656) );
  DFF_X1 new_AGEMA_reg_buffer_3772_s_current_state_reg ( .D(
        new_AGEMA_signal_5659), .CK(clk), .Q(new_AGEMA_signal_5660) );
  DFF_X1 new_AGEMA_reg_buffer_3776_s_current_state_reg ( .D(
        new_AGEMA_signal_5663), .CK(clk), .Q(new_AGEMA_signal_5664) );
  DFF_X1 new_AGEMA_reg_buffer_3780_s_current_state_reg ( .D(
        new_AGEMA_signal_5667), .CK(clk), .Q(new_AGEMA_signal_5668) );
  DFF_X1 new_AGEMA_reg_buffer_3784_s_current_state_reg ( .D(
        new_AGEMA_signal_5671), .CK(clk), .Q(new_AGEMA_signal_5672) );
  DFF_X1 new_AGEMA_reg_buffer_3788_s_current_state_reg ( .D(
        new_AGEMA_signal_5675), .CK(clk), .Q(new_AGEMA_signal_5676) );
  DFF_X1 new_AGEMA_reg_buffer_3792_s_current_state_reg ( .D(
        new_AGEMA_signal_5679), .CK(clk), .Q(new_AGEMA_signal_5680) );
  DFF_X1 new_AGEMA_reg_buffer_3796_s_current_state_reg ( .D(
        new_AGEMA_signal_5683), .CK(clk), .Q(new_AGEMA_signal_5684) );
  DFF_X1 new_AGEMA_reg_buffer_3800_s_current_state_reg ( .D(
        new_AGEMA_signal_5687), .CK(clk), .Q(new_AGEMA_signal_5688) );
  DFF_X1 new_AGEMA_reg_buffer_3804_s_current_state_reg ( .D(
        new_AGEMA_signal_5691), .CK(clk), .Q(new_AGEMA_signal_5692) );
  DFF_X1 new_AGEMA_reg_buffer_3808_s_current_state_reg ( .D(
        new_AGEMA_signal_5695), .CK(clk), .Q(new_AGEMA_signal_5696) );
  DFF_X1 new_AGEMA_reg_buffer_3812_s_current_state_reg ( .D(
        new_AGEMA_signal_5699), .CK(clk), .Q(new_AGEMA_signal_5700) );
  DFF_X1 new_AGEMA_reg_buffer_3816_s_current_state_reg ( .D(
        new_AGEMA_signal_5703), .CK(clk), .Q(new_AGEMA_signal_5704) );
  DFF_X1 new_AGEMA_reg_buffer_3820_s_current_state_reg ( .D(
        new_AGEMA_signal_5707), .CK(clk), .Q(new_AGEMA_signal_5708) );
  DFF_X1 new_AGEMA_reg_buffer_3824_s_current_state_reg ( .D(
        new_AGEMA_signal_5711), .CK(clk), .Q(new_AGEMA_signal_5712) );
  DFF_X1 new_AGEMA_reg_buffer_3828_s_current_state_reg ( .D(
        new_AGEMA_signal_5715), .CK(clk), .Q(new_AGEMA_signal_5716) );
  DFF_X1 new_AGEMA_reg_buffer_3832_s_current_state_reg ( .D(
        new_AGEMA_signal_5719), .CK(clk), .Q(new_AGEMA_signal_5720) );
  DFF_X1 new_AGEMA_reg_buffer_3836_s_current_state_reg ( .D(
        new_AGEMA_signal_5723), .CK(clk), .Q(new_AGEMA_signal_5724) );
  DFF_X1 new_AGEMA_reg_buffer_3840_s_current_state_reg ( .D(
        new_AGEMA_signal_5727), .CK(clk), .Q(new_AGEMA_signal_5728) );
  DFF_X1 new_AGEMA_reg_buffer_3844_s_current_state_reg ( .D(
        new_AGEMA_signal_5731), .CK(clk), .Q(new_AGEMA_signal_5732) );
  DFF_X1 new_AGEMA_reg_buffer_3848_s_current_state_reg ( .D(
        new_AGEMA_signal_5735), .CK(clk), .Q(new_AGEMA_signal_5736) );
  DFF_X1 new_AGEMA_reg_buffer_3852_s_current_state_reg ( .D(
        new_AGEMA_signal_5739), .CK(clk), .Q(new_AGEMA_signal_5740) );
  DFF_X1 new_AGEMA_reg_buffer_3856_s_current_state_reg ( .D(
        new_AGEMA_signal_5743), .CK(clk), .Q(new_AGEMA_signal_5744) );
  DFF_X1 new_AGEMA_reg_buffer_3860_s_current_state_reg ( .D(
        new_AGEMA_signal_5747), .CK(clk), .Q(new_AGEMA_signal_5748) );
  DFF_X1 new_AGEMA_reg_buffer_3864_s_current_state_reg ( .D(
        new_AGEMA_signal_5751), .CK(clk), .Q(new_AGEMA_signal_5752) );
  DFF_X1 new_AGEMA_reg_buffer_3868_s_current_state_reg ( .D(
        new_AGEMA_signal_5755), .CK(clk), .Q(new_AGEMA_signal_5756) );
  DFF_X1 new_AGEMA_reg_buffer_3872_s_current_state_reg ( .D(
        new_AGEMA_signal_5759), .CK(clk), .Q(new_AGEMA_signal_5760) );
  DFF_X1 new_AGEMA_reg_buffer_3876_s_current_state_reg ( .D(
        new_AGEMA_signal_5763), .CK(clk), .Q(new_AGEMA_signal_5764) );
  DFF_X1 new_AGEMA_reg_buffer_3880_s_current_state_reg ( .D(
        new_AGEMA_signal_5767), .CK(clk), .Q(new_AGEMA_signal_5768) );
  DFF_X1 new_AGEMA_reg_buffer_3884_s_current_state_reg ( .D(
        new_AGEMA_signal_5771), .CK(clk), .Q(new_AGEMA_signal_5772) );
  DFF_X1 new_AGEMA_reg_buffer_3888_s_current_state_reg ( .D(
        new_AGEMA_signal_5775), .CK(clk), .Q(new_AGEMA_signal_5776) );
  DFF_X1 new_AGEMA_reg_buffer_3892_s_current_state_reg ( .D(
        new_AGEMA_signal_5779), .CK(clk), .Q(new_AGEMA_signal_5780) );
  DFF_X1 new_AGEMA_reg_buffer_3896_s_current_state_reg ( .D(
        new_AGEMA_signal_5783), .CK(clk), .Q(new_AGEMA_signal_5784) );
  DFF_X1 new_AGEMA_reg_buffer_3900_s_current_state_reg ( .D(
        new_AGEMA_signal_5787), .CK(clk), .Q(new_AGEMA_signal_5788) );
  DFF_X1 new_AGEMA_reg_buffer_3904_s_current_state_reg ( .D(
        new_AGEMA_signal_5791), .CK(clk), .Q(new_AGEMA_signal_5792) );
  DFF_X1 new_AGEMA_reg_buffer_3908_s_current_state_reg ( .D(
        new_AGEMA_signal_5795), .CK(clk), .Q(new_AGEMA_signal_5796) );
  DFF_X1 new_AGEMA_reg_buffer_3912_s_current_state_reg ( .D(
        new_AGEMA_signal_5799), .CK(clk), .Q(new_AGEMA_signal_5800) );
  DFF_X1 new_AGEMA_reg_buffer_3916_s_current_state_reg ( .D(
        new_AGEMA_signal_5803), .CK(clk), .Q(new_AGEMA_signal_5804) );
  DFF_X1 new_AGEMA_reg_buffer_3920_s_current_state_reg ( .D(
        new_AGEMA_signal_5807), .CK(clk), .Q(new_AGEMA_signal_5808) );
  DFF_X1 new_AGEMA_reg_buffer_3924_s_current_state_reg ( .D(
        new_AGEMA_signal_5811), .CK(clk), .Q(new_AGEMA_signal_5812) );
  DFF_X1 new_AGEMA_reg_buffer_3928_s_current_state_reg ( .D(
        new_AGEMA_signal_5815), .CK(clk), .Q(new_AGEMA_signal_5816) );
  DFF_X1 new_AGEMA_reg_buffer_3932_s_current_state_reg ( .D(
        new_AGEMA_signal_5819), .CK(clk), .Q(new_AGEMA_signal_5820) );
  DFF_X1 new_AGEMA_reg_buffer_3936_s_current_state_reg ( .D(
        new_AGEMA_signal_5823), .CK(clk), .Q(new_AGEMA_signal_5824) );
  DFF_X1 new_AGEMA_reg_buffer_3940_s_current_state_reg ( .D(
        new_AGEMA_signal_5827), .CK(clk), .Q(new_AGEMA_signal_5828) );
  DFF_X1 new_AGEMA_reg_buffer_3944_s_current_state_reg ( .D(
        new_AGEMA_signal_5831), .CK(clk), .Q(new_AGEMA_signal_5832) );
  DFF_X1 new_AGEMA_reg_buffer_3948_s_current_state_reg ( .D(
        new_AGEMA_signal_5835), .CK(clk), .Q(new_AGEMA_signal_5836) );
  DFF_X1 new_AGEMA_reg_buffer_3952_s_current_state_reg ( .D(
        new_AGEMA_signal_5839), .CK(clk), .Q(new_AGEMA_signal_5840) );
  DFF_X1 new_AGEMA_reg_buffer_3956_s_current_state_reg ( .D(
        new_AGEMA_signal_5843), .CK(clk), .Q(new_AGEMA_signal_5844) );
  DFF_X1 new_AGEMA_reg_buffer_3960_s_current_state_reg ( .D(
        new_AGEMA_signal_5847), .CK(clk), .Q(new_AGEMA_signal_5848) );
  DFF_X1 new_AGEMA_reg_buffer_3964_s_current_state_reg ( .D(
        new_AGEMA_signal_5851), .CK(clk), .Q(new_AGEMA_signal_5852) );
  DFF_X1 new_AGEMA_reg_buffer_3968_s_current_state_reg ( .D(
        new_AGEMA_signal_5855), .CK(clk), .Q(new_AGEMA_signal_5856) );
  DFF_X1 new_AGEMA_reg_buffer_3972_s_current_state_reg ( .D(
        new_AGEMA_signal_5859), .CK(clk), .Q(new_AGEMA_signal_5860) );
  DFF_X1 new_AGEMA_reg_buffer_3976_s_current_state_reg ( .D(
        new_AGEMA_signal_5863), .CK(clk), .Q(new_AGEMA_signal_5864) );
  DFF_X1 new_AGEMA_reg_buffer_3980_s_current_state_reg ( .D(
        new_AGEMA_signal_5867), .CK(clk), .Q(new_AGEMA_signal_5868) );
  DFF_X1 new_AGEMA_reg_buffer_3984_s_current_state_reg ( .D(
        new_AGEMA_signal_5871), .CK(clk), .Q(new_AGEMA_signal_5872) );
  DFF_X1 new_AGEMA_reg_buffer_3988_s_current_state_reg ( .D(
        new_AGEMA_signal_5875), .CK(clk), .Q(new_AGEMA_signal_5876) );
  DFF_X1 new_AGEMA_reg_buffer_3992_s_current_state_reg ( .D(
        new_AGEMA_signal_5879), .CK(clk), .Q(new_AGEMA_signal_5880) );
  DFF_X1 new_AGEMA_reg_buffer_3996_s_current_state_reg ( .D(
        new_AGEMA_signal_5883), .CK(clk), .Q(new_AGEMA_signal_5884) );
  DFF_X1 new_AGEMA_reg_buffer_4000_s_current_state_reg ( .D(
        new_AGEMA_signal_5887), .CK(clk), .Q(new_AGEMA_signal_5888) );
  DFF_X1 new_AGEMA_reg_buffer_4004_s_current_state_reg ( .D(
        new_AGEMA_signal_5891), .CK(clk), .Q(new_AGEMA_signal_5892) );
  DFF_X1 new_AGEMA_reg_buffer_4008_s_current_state_reg ( .D(
        new_AGEMA_signal_5895), .CK(clk), .Q(new_AGEMA_signal_5896) );
  DFF_X1 new_AGEMA_reg_buffer_4012_s_current_state_reg ( .D(
        new_AGEMA_signal_5899), .CK(clk), .Q(new_AGEMA_signal_5900) );
  DFF_X1 new_AGEMA_reg_buffer_4016_s_current_state_reg ( .D(
        new_AGEMA_signal_5903), .CK(clk), .Q(new_AGEMA_signal_5904) );
  DFF_X1 new_AGEMA_reg_buffer_4020_s_current_state_reg ( .D(
        new_AGEMA_signal_5907), .CK(clk), .Q(new_AGEMA_signal_5908) );
  DFF_X1 new_AGEMA_reg_buffer_4024_s_current_state_reg ( .D(
        new_AGEMA_signal_5911), .CK(clk), .Q(new_AGEMA_signal_5912) );
  DFF_X1 new_AGEMA_reg_buffer_4028_s_current_state_reg ( .D(
        new_AGEMA_signal_5915), .CK(clk), .Q(new_AGEMA_signal_5916) );
  DFF_X1 new_AGEMA_reg_buffer_4032_s_current_state_reg ( .D(
        new_AGEMA_signal_5919), .CK(clk), .Q(new_AGEMA_signal_5920) );
  DFF_X1 new_AGEMA_reg_buffer_4036_s_current_state_reg ( .D(
        new_AGEMA_signal_5923), .CK(clk), .Q(new_AGEMA_signal_5924) );
  DFF_X1 new_AGEMA_reg_buffer_4040_s_current_state_reg ( .D(
        new_AGEMA_signal_5927), .CK(clk), .Q(new_AGEMA_signal_5928) );
  DFF_X1 new_AGEMA_reg_buffer_4044_s_current_state_reg ( .D(
        new_AGEMA_signal_5931), .CK(clk), .Q(new_AGEMA_signal_5932) );
  DFF_X1 new_AGEMA_reg_buffer_4048_s_current_state_reg ( .D(
        new_AGEMA_signal_5935), .CK(clk), .Q(new_AGEMA_signal_5936) );
  DFF_X1 new_AGEMA_reg_buffer_4052_s_current_state_reg ( .D(
        new_AGEMA_signal_5939), .CK(clk), .Q(new_AGEMA_signal_5940) );
  DFF_X1 new_AGEMA_reg_buffer_4056_s_current_state_reg ( .D(
        new_AGEMA_signal_5943), .CK(clk), .Q(new_AGEMA_signal_5944) );
  DFF_X1 new_AGEMA_reg_buffer_4060_s_current_state_reg ( .D(
        new_AGEMA_signal_5947), .CK(clk), .Q(new_AGEMA_signal_5948) );
  DFF_X1 new_AGEMA_reg_buffer_4064_s_current_state_reg ( .D(
        new_AGEMA_signal_5951), .CK(clk), .Q(new_AGEMA_signal_5952) );
  DFF_X1 new_AGEMA_reg_buffer_4068_s_current_state_reg ( .D(
        new_AGEMA_signal_5955), .CK(clk), .Q(new_AGEMA_signal_5956) );
  DFF_X1 new_AGEMA_reg_buffer_4072_s_current_state_reg ( .D(
        new_AGEMA_signal_5959), .CK(clk), .Q(new_AGEMA_signal_5960) );
  DFF_X1 new_AGEMA_reg_buffer_4076_s_current_state_reg ( .D(
        new_AGEMA_signal_5963), .CK(clk), .Q(new_AGEMA_signal_5964) );
  DFF_X1 new_AGEMA_reg_buffer_4080_s_current_state_reg ( .D(
        new_AGEMA_signal_5967), .CK(clk), .Q(new_AGEMA_signal_5968) );
  DFF_X1 new_AGEMA_reg_buffer_4084_s_current_state_reg ( .D(
        new_AGEMA_signal_5971), .CK(clk), .Q(new_AGEMA_signal_5972) );
  DFF_X1 new_AGEMA_reg_buffer_4088_s_current_state_reg ( .D(
        new_AGEMA_signal_5975), .CK(clk), .Q(new_AGEMA_signal_5976) );
  DFF_X1 new_AGEMA_reg_buffer_4092_s_current_state_reg ( .D(
        new_AGEMA_signal_5979), .CK(clk), .Q(new_AGEMA_signal_5980) );
  DFF_X1 new_AGEMA_reg_buffer_4096_s_current_state_reg ( .D(
        new_AGEMA_signal_5983), .CK(clk), .Q(new_AGEMA_signal_5984) );
  DFF_X1 new_AGEMA_reg_buffer_4100_s_current_state_reg ( .D(
        new_AGEMA_signal_5987), .CK(clk), .Q(new_AGEMA_signal_5988) );
  DFF_X1 new_AGEMA_reg_buffer_4104_s_current_state_reg ( .D(
        new_AGEMA_signal_5991), .CK(clk), .Q(new_AGEMA_signal_5992) );
  DFF_X1 new_AGEMA_reg_buffer_4108_s_current_state_reg ( .D(
        new_AGEMA_signal_5995), .CK(clk), .Q(new_AGEMA_signal_5996) );
  DFF_X1 new_AGEMA_reg_buffer_4112_s_current_state_reg ( .D(
        new_AGEMA_signal_5999), .CK(clk), .Q(new_AGEMA_signal_6000) );
  DFF_X1 new_AGEMA_reg_buffer_4116_s_current_state_reg ( .D(
        new_AGEMA_signal_6003), .CK(clk), .Q(new_AGEMA_signal_6004) );
  DFF_X1 new_AGEMA_reg_buffer_4120_s_current_state_reg ( .D(
        new_AGEMA_signal_6007), .CK(clk), .Q(new_AGEMA_signal_6008) );
  DFF_X1 new_AGEMA_reg_buffer_4124_s_current_state_reg ( .D(
        new_AGEMA_signal_6011), .CK(clk), .Q(new_AGEMA_signal_6012) );
  DFF_X1 new_AGEMA_reg_buffer_4128_s_current_state_reg ( .D(
        new_AGEMA_signal_6015), .CK(clk), .Q(new_AGEMA_signal_6016) );
  DFF_X1 new_AGEMA_reg_buffer_4132_s_current_state_reg ( .D(
        new_AGEMA_signal_6019), .CK(clk), .Q(new_AGEMA_signal_6020) );
  DFF_X1 new_AGEMA_reg_buffer_4136_s_current_state_reg ( .D(
        new_AGEMA_signal_6023), .CK(clk), .Q(new_AGEMA_signal_6024) );
  DFF_X1 new_AGEMA_reg_buffer_4140_s_current_state_reg ( .D(
        new_AGEMA_signal_6027), .CK(clk), .Q(new_AGEMA_signal_6028) );
  DFF_X1 new_AGEMA_reg_buffer_4144_s_current_state_reg ( .D(
        new_AGEMA_signal_6031), .CK(clk), .Q(new_AGEMA_signal_6032) );
  DFF_X1 new_AGEMA_reg_buffer_4148_s_current_state_reg ( .D(
        new_AGEMA_signal_6035), .CK(clk), .Q(new_AGEMA_signal_6036) );
  DFF_X1 new_AGEMA_reg_buffer_4152_s_current_state_reg ( .D(
        new_AGEMA_signal_6039), .CK(clk), .Q(new_AGEMA_signal_6040) );
  DFF_X1 new_AGEMA_reg_buffer_4156_s_current_state_reg ( .D(
        new_AGEMA_signal_6043), .CK(clk), .Q(new_AGEMA_signal_6044) );
  DFF_X1 new_AGEMA_reg_buffer_4160_s_current_state_reg ( .D(
        new_AGEMA_signal_6047), .CK(clk), .Q(new_AGEMA_signal_6048) );
  DFF_X1 new_AGEMA_reg_buffer_4164_s_current_state_reg ( .D(
        new_AGEMA_signal_6051), .CK(clk), .Q(new_AGEMA_signal_6052) );
  DFF_X1 new_AGEMA_reg_buffer_4168_s_current_state_reg ( .D(
        new_AGEMA_signal_6055), .CK(clk), .Q(new_AGEMA_signal_6056) );
  DFF_X1 new_AGEMA_reg_buffer_4172_s_current_state_reg ( .D(
        new_AGEMA_signal_6059), .CK(clk), .Q(new_AGEMA_signal_6060) );
  DFF_X1 new_AGEMA_reg_buffer_4176_s_current_state_reg ( .D(
        new_AGEMA_signal_6063), .CK(clk), .Q(new_AGEMA_signal_6064) );
  DFF_X1 new_AGEMA_reg_buffer_4180_s_current_state_reg ( .D(
        new_AGEMA_signal_6067), .CK(clk), .Q(new_AGEMA_signal_6068) );
  DFF_X1 new_AGEMA_reg_buffer_4184_s_current_state_reg ( .D(
        new_AGEMA_signal_6071), .CK(clk), .Q(new_AGEMA_signal_6072) );
  DFF_X1 new_AGEMA_reg_buffer_4188_s_current_state_reg ( .D(
        new_AGEMA_signal_6075), .CK(clk), .Q(new_AGEMA_signal_6076) );
  DFF_X1 new_AGEMA_reg_buffer_4192_s_current_state_reg ( .D(
        new_AGEMA_signal_6079), .CK(clk), .Q(new_AGEMA_signal_6080) );
  DFF_X1 new_AGEMA_reg_buffer_4196_s_current_state_reg ( .D(
        new_AGEMA_signal_6083), .CK(clk), .Q(new_AGEMA_signal_6084) );
  DFF_X1 new_AGEMA_reg_buffer_4200_s_current_state_reg ( .D(
        new_AGEMA_signal_6087), .CK(clk), .Q(new_AGEMA_signal_6088) );
  DFF_X1 new_AGEMA_reg_buffer_4204_s_current_state_reg ( .D(
        new_AGEMA_signal_6091), .CK(clk), .Q(new_AGEMA_signal_6092) );
  DFF_X1 new_AGEMA_reg_buffer_4208_s_current_state_reg ( .D(
        new_AGEMA_signal_6095), .CK(clk), .Q(new_AGEMA_signal_6096) );
  DFF_X1 new_AGEMA_reg_buffer_4212_s_current_state_reg ( .D(
        new_AGEMA_signal_6099), .CK(clk), .Q(new_AGEMA_signal_6100) );
  DFF_X1 new_AGEMA_reg_buffer_4216_s_current_state_reg ( .D(
        new_AGEMA_signal_6103), .CK(clk), .Q(new_AGEMA_signal_6104) );
  DFF_X1 new_AGEMA_reg_buffer_4220_s_current_state_reg ( .D(
        new_AGEMA_signal_6107), .CK(clk), .Q(new_AGEMA_signal_6108) );
  DFF_X1 new_AGEMA_reg_buffer_4224_s_current_state_reg ( .D(
        new_AGEMA_signal_6111), .CK(clk), .Q(new_AGEMA_signal_6112) );
  DFF_X1 new_AGEMA_reg_buffer_4228_s_current_state_reg ( .D(
        new_AGEMA_signal_6115), .CK(clk), .Q(new_AGEMA_signal_6116) );
  DFF_X1 new_AGEMA_reg_buffer_4232_s_current_state_reg ( .D(
        new_AGEMA_signal_6119), .CK(clk), .Q(new_AGEMA_signal_6120) );
  DFF_X1 new_AGEMA_reg_buffer_4236_s_current_state_reg ( .D(
        new_AGEMA_signal_6123), .CK(clk), .Q(new_AGEMA_signal_6124) );
  DFF_X1 new_AGEMA_reg_buffer_4240_s_current_state_reg ( .D(
        new_AGEMA_signal_6127), .CK(clk), .Q(new_AGEMA_signal_6128) );
  DFF_X1 new_AGEMA_reg_buffer_4244_s_current_state_reg ( .D(
        new_AGEMA_signal_6131), .CK(clk), .Q(new_AGEMA_signal_6132) );
  DFF_X1 new_AGEMA_reg_buffer_4248_s_current_state_reg ( .D(
        new_AGEMA_signal_6135), .CK(clk), .Q(new_AGEMA_signal_6136) );
  DFF_X1 new_AGEMA_reg_buffer_4252_s_current_state_reg ( .D(
        new_AGEMA_signal_6139), .CK(clk), .Q(new_AGEMA_signal_6140) );
  DFF_X1 new_AGEMA_reg_buffer_4256_s_current_state_reg ( .D(
        new_AGEMA_signal_6143), .CK(clk), .Q(new_AGEMA_signal_6144) );
  DFF_X1 new_AGEMA_reg_buffer_4260_s_current_state_reg ( .D(
        new_AGEMA_signal_6147), .CK(clk), .Q(new_AGEMA_signal_6148) );
  DFF_X1 new_AGEMA_reg_buffer_4264_s_current_state_reg ( .D(
        new_AGEMA_signal_6151), .CK(clk), .Q(new_AGEMA_signal_6152) );
  DFF_X1 new_AGEMA_reg_buffer_4268_s_current_state_reg ( .D(
        new_AGEMA_signal_6155), .CK(clk), .Q(new_AGEMA_signal_6156) );
  DFF_X1 new_AGEMA_reg_buffer_4272_s_current_state_reg ( .D(
        new_AGEMA_signal_6159), .CK(clk), .Q(new_AGEMA_signal_6160) );
  DFF_X1 new_AGEMA_reg_buffer_4276_s_current_state_reg ( .D(
        new_AGEMA_signal_6163), .CK(clk), .Q(new_AGEMA_signal_6164) );
  DFF_X1 new_AGEMA_reg_buffer_4280_s_current_state_reg ( .D(
        new_AGEMA_signal_6167), .CK(clk), .Q(new_AGEMA_signal_6168) );
  DFF_X1 new_AGEMA_reg_buffer_4284_s_current_state_reg ( .D(
        new_AGEMA_signal_6171), .CK(clk), .Q(new_AGEMA_signal_6172) );
  DFF_X1 new_AGEMA_reg_buffer_4288_s_current_state_reg ( .D(
        new_AGEMA_signal_6175), .CK(clk), .Q(new_AGEMA_signal_6176) );
  DFF_X1 new_AGEMA_reg_buffer_4292_s_current_state_reg ( .D(
        new_AGEMA_signal_6179), .CK(clk), .Q(new_AGEMA_signal_6180) );
  DFF_X1 new_AGEMA_reg_buffer_4296_s_current_state_reg ( .D(
        new_AGEMA_signal_6183), .CK(clk), .Q(new_AGEMA_signal_6184) );
  DFF_X1 new_AGEMA_reg_buffer_4300_s_current_state_reg ( .D(
        new_AGEMA_signal_6187), .CK(clk), .Q(new_AGEMA_signal_6188) );
  DFF_X1 new_AGEMA_reg_buffer_4304_s_current_state_reg ( .D(
        new_AGEMA_signal_6191), .CK(clk), .Q(new_AGEMA_signal_6192) );
  DFF_X1 new_AGEMA_reg_buffer_4308_s_current_state_reg ( .D(
        new_AGEMA_signal_6195), .CK(clk), .Q(new_AGEMA_signal_6196) );
  DFF_X1 new_AGEMA_reg_buffer_4312_s_current_state_reg ( .D(
        new_AGEMA_signal_6199), .CK(clk), .Q(new_AGEMA_signal_6200) );
  DFF_X1 new_AGEMA_reg_buffer_4316_s_current_state_reg ( .D(
        new_AGEMA_signal_6203), .CK(clk), .Q(new_AGEMA_signal_6204) );
  DFF_X1 new_AGEMA_reg_buffer_4320_s_current_state_reg ( .D(
        new_AGEMA_signal_6207), .CK(clk), .Q(new_AGEMA_signal_6208) );
  DFF_X1 new_AGEMA_reg_buffer_4324_s_current_state_reg ( .D(
        new_AGEMA_signal_6211), .CK(clk), .Q(new_AGEMA_signal_6212) );
  DFF_X1 new_AGEMA_reg_buffer_4328_s_current_state_reg ( .D(
        new_AGEMA_signal_6215), .CK(clk), .Q(new_AGEMA_signal_6216) );
  DFF_X1 new_AGEMA_reg_buffer_4332_s_current_state_reg ( .D(
        new_AGEMA_signal_6219), .CK(clk), .Q(new_AGEMA_signal_6220) );
  DFF_X1 new_AGEMA_reg_buffer_4336_s_current_state_reg ( .D(
        new_AGEMA_signal_6223), .CK(clk), .Q(new_AGEMA_signal_6224) );
  DFF_X1 new_AGEMA_reg_buffer_4340_s_current_state_reg ( .D(
        new_AGEMA_signal_6227), .CK(clk), .Q(new_AGEMA_signal_6228) );
  NAND2_X1 MUX_StateIn_mux_inst_0_U1_Ins_0_U4 ( .A1(
        MUX_StateIn_mux_inst_0_U1_Ins_0_n8), .A2(
        MUX_StateIn_mux_inst_0_U1_Ins_0_n7), .ZN(StateIn[0]) );
  NAND2_X1 MUX_StateIn_mux_inst_0_U1_Ins_0_U3 ( .A1(SboxOut[0]), .A2(
        MUX_StateIn_mux_inst_0_U1_Ins_0_n6), .ZN(
        MUX_StateIn_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 MUX_StateIn_mux_inst_0_U1_Ins_0_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_0_U1_Ins_0_U1 ( .A1(new_AGEMA_signal_3633),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_0_U1_Ins_1_U4 ( .A1(
        MUX_StateIn_mux_inst_0_U1_Ins_1_n8), .A2(
        MUX_StateIn_mux_inst_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3455) );
  NAND2_X1 MUX_StateIn_mux_inst_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_3456),
        .A2(MUX_StateIn_mux_inst_0_U1_Ins_1_n6), .ZN(
        MUX_StateIn_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 MUX_StateIn_mux_inst_0_U1_Ins_1_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3637),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_1_U1_Ins_0_U4 ( .A1(
        MUX_StateIn_mux_inst_1_U1_Ins_0_n8), .A2(
        MUX_StateIn_mux_inst_1_U1_Ins_0_n7), .ZN(StateIn[1]) );
  NAND2_X1 MUX_StateIn_mux_inst_1_U1_Ins_0_U3 ( .A1(SboxOut[1]), .A2(
        MUX_StateIn_mux_inst_1_U1_Ins_0_n6), .ZN(
        MUX_StateIn_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 MUX_StateIn_mux_inst_1_U1_Ins_0_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_1_U1_Ins_0_U1 ( .A1(new_AGEMA_signal_3641),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_1_U1_Ins_1_U4 ( .A1(
        MUX_StateIn_mux_inst_1_U1_Ins_1_n8), .A2(
        MUX_StateIn_mux_inst_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3464) );
  NAND2_X1 MUX_StateIn_mux_inst_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_3478),
        .A2(MUX_StateIn_mux_inst_1_U1_Ins_1_n6), .ZN(
        MUX_StateIn_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 MUX_StateIn_mux_inst_1_U1_Ins_1_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3645),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_2_U1_Ins_0_U4 ( .A1(
        MUX_StateIn_mux_inst_2_U1_Ins_0_n8), .A2(
        MUX_StateIn_mux_inst_2_U1_Ins_0_n7), .ZN(StateIn[2]) );
  NAND2_X1 MUX_StateIn_mux_inst_2_U1_Ins_0_U3 ( .A1(SboxOut[2]), .A2(
        MUX_StateIn_mux_inst_2_U1_Ins_0_n6), .ZN(
        MUX_StateIn_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 MUX_StateIn_mux_inst_2_U1_Ins_0_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_2_U1_Ins_0_U1 ( .A1(new_AGEMA_signal_3649),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_2_U1_Ins_1_U4 ( .A1(
        MUX_StateIn_mux_inst_2_U1_Ins_1_n8), .A2(
        MUX_StateIn_mux_inst_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3465) );
  NAND2_X1 MUX_StateIn_mux_inst_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_3477),
        .A2(MUX_StateIn_mux_inst_2_U1_Ins_1_n6), .ZN(
        MUX_StateIn_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 MUX_StateIn_mux_inst_2_U1_Ins_1_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3653),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_3_U1_Ins_0_U4 ( .A1(
        MUX_StateIn_mux_inst_3_U1_Ins_0_n8), .A2(
        MUX_StateIn_mux_inst_3_U1_Ins_0_n7), .ZN(StateIn[3]) );
  NAND2_X1 MUX_StateIn_mux_inst_3_U1_Ins_0_U3 ( .A1(SboxOut[3]), .A2(
        MUX_StateIn_mux_inst_3_U1_Ins_0_n6), .ZN(
        MUX_StateIn_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 MUX_StateIn_mux_inst_3_U1_Ins_0_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_3_U1_Ins_0_U1 ( .A1(new_AGEMA_signal_3657),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_3_U1_Ins_1_U4 ( .A1(
        MUX_StateIn_mux_inst_3_U1_Ins_1_n8), .A2(
        MUX_StateIn_mux_inst_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3466) );
  NAND2_X1 MUX_StateIn_mux_inst_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_3476),
        .A2(MUX_StateIn_mux_inst_3_U1_Ins_1_n6), .ZN(
        MUX_StateIn_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 MUX_StateIn_mux_inst_3_U1_Ins_1_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3661),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_4_U1_Ins_0_U4 ( .A1(
        MUX_StateIn_mux_inst_4_U1_Ins_0_n8), .A2(
        MUX_StateIn_mux_inst_4_U1_Ins_0_n7), .ZN(StateIn[4]) );
  NAND2_X1 MUX_StateIn_mux_inst_4_U1_Ins_0_U3 ( .A1(SboxOut[4]), .A2(
        MUX_StateIn_mux_inst_4_U1_Ins_0_n6), .ZN(
        MUX_StateIn_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 MUX_StateIn_mux_inst_4_U1_Ins_0_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_4_U1_Ins_0_U1 ( .A1(new_AGEMA_signal_3665),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_4_U1_Ins_1_U4 ( .A1(
        MUX_StateIn_mux_inst_4_U1_Ins_1_n8), .A2(
        MUX_StateIn_mux_inst_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3467) );
  NAND2_X1 MUX_StateIn_mux_inst_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_3475),
        .A2(MUX_StateIn_mux_inst_4_U1_Ins_1_n6), .ZN(
        MUX_StateIn_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 MUX_StateIn_mux_inst_4_U1_Ins_1_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3669),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_5_U1_Ins_0_U4 ( .A1(
        MUX_StateIn_mux_inst_5_U1_Ins_0_n8), .A2(
        MUX_StateIn_mux_inst_5_U1_Ins_0_n7), .ZN(StateIn[5]) );
  NAND2_X1 MUX_StateIn_mux_inst_5_U1_Ins_0_U3 ( .A1(SboxOut[5]), .A2(
        MUX_StateIn_mux_inst_5_U1_Ins_0_n6), .ZN(
        MUX_StateIn_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 MUX_StateIn_mux_inst_5_U1_Ins_0_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_5_U1_Ins_0_U1 ( .A1(new_AGEMA_signal_3673),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_5_U1_Ins_1_U4 ( .A1(
        MUX_StateIn_mux_inst_5_U1_Ins_1_n8), .A2(
        MUX_StateIn_mux_inst_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3468) );
  NAND2_X1 MUX_StateIn_mux_inst_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_3474),
        .A2(MUX_StateIn_mux_inst_5_U1_Ins_1_n6), .ZN(
        MUX_StateIn_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 MUX_StateIn_mux_inst_5_U1_Ins_1_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3677),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_6_U1_Ins_0_U4 ( .A1(
        MUX_StateIn_mux_inst_6_U1_Ins_0_n8), .A2(
        MUX_StateIn_mux_inst_6_U1_Ins_0_n7), .ZN(StateIn[6]) );
  NAND2_X1 MUX_StateIn_mux_inst_6_U1_Ins_0_U3 ( .A1(SboxOut[6]), .A2(
        MUX_StateIn_mux_inst_6_U1_Ins_0_n6), .ZN(
        MUX_StateIn_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 MUX_StateIn_mux_inst_6_U1_Ins_0_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_6_U1_Ins_0_U1 ( .A1(new_AGEMA_signal_3681),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_6_U1_Ins_1_U4 ( .A1(
        MUX_StateIn_mux_inst_6_U1_Ins_1_n8), .A2(
        MUX_StateIn_mux_inst_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3469) );
  NAND2_X1 MUX_StateIn_mux_inst_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_3473),
        .A2(MUX_StateIn_mux_inst_6_U1_Ins_1_n6), .ZN(
        MUX_StateIn_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 MUX_StateIn_mux_inst_6_U1_Ins_1_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3685),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_7_U1_Ins_0_U4 ( .A1(
        MUX_StateIn_mux_inst_7_U1_Ins_0_n8), .A2(
        MUX_StateIn_mux_inst_7_U1_Ins_0_n7), .ZN(StateIn[7]) );
  NAND2_X1 MUX_StateIn_mux_inst_7_U1_Ins_0_U3 ( .A1(SboxOut[7]), .A2(
        MUX_StateIn_mux_inst_7_U1_Ins_0_n6), .ZN(
        MUX_StateIn_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 MUX_StateIn_mux_inst_7_U1_Ins_0_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_7_U1_Ins_0_U1 ( .A1(new_AGEMA_signal_3689),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 MUX_StateIn_mux_inst_7_U1_Ins_1_U4 ( .A1(
        MUX_StateIn_mux_inst_7_U1_Ins_1_n8), .A2(
        MUX_StateIn_mux_inst_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3470) );
  NAND2_X1 MUX_StateIn_mux_inst_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_3472),
        .A2(MUX_StateIn_mux_inst_7_U1_Ins_1_n6), .ZN(
        MUX_StateIn_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 MUX_StateIn_mux_inst_7_U1_Ins_1_U2 ( .A(n287), .ZN(
        MUX_StateIn_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 MUX_StateIn_mux_inst_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3693),
        .A2(n287), .ZN(MUX_StateIn_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S33reg_gff_1_SFF_0_QD) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS33ser[0]), .A2(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3701), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3497) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3488), .A2(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3705), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S33reg_gff_1_SFF_1_QD) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS33ser[1]), .A2(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3709), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3520) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3499), .A2(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3713), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S33reg_gff_1_SFF_2_QD) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS33ser[2]), .A2(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3717), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3521) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3501), .A2(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3721), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S33reg_gff_1_SFF_3_QD) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS33ser[3]), .A2(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3725), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3522) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3503), .A2(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3729), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S33reg_gff_1_SFF_4_QD) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS33ser[4]), .A2(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3733), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3523) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3505), .A2(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3737), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S33reg_gff_1_SFF_5_QD) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS33ser[5]), .A2(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3741), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3524) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3507), .A2(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3745), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S33reg_gff_1_SFF_6_QD) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS33ser[6]), .A2(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3749), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3525) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3509), .A2(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3753), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        stateArray_S33reg_gff_1_SFF_7_QD) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        stateArray_inS33ser[7]), .A2(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3757), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3526) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3511), .A2(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3761), .A2(n286), .ZN(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_input_MC[0]) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_U3 ( .A1(StateIn[0]),
        .A2(stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3769), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3471) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3455), .A2(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3773), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_input_MC[1]) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_U3 ( .A1(StateIn[1]),
        .A2(stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3777), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3480) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3464), .A2(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3781), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_input_MC[2]) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_U3 ( .A1(StateIn[2]),
        .A2(stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3785), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3481) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3465), .A2(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3789), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_input_MC[3]) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_U3 ( .A1(StateIn[3]),
        .A2(stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3793), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3482) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3466), .A2(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3797), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_input_MC[4]) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_U3 ( .A1(StateIn[4]),
        .A2(stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3801), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3483) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3467), .A2(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3805), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_input_MC[5]) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_U3 ( .A1(StateIn[5]),
        .A2(stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3809), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3484) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3468), .A2(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3813), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_input_MC[6]) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_U3 ( .A1(StateIn[6]),
        .A2(stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3817), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3485) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3469), .A2(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3821), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_input_MC[7]) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_U3 ( .A1(StateIn[7]),
        .A2(stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_U1 ( .A1(
        new_AGEMA_signal_3825), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3486) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3470), .A2(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_n6), .ZN(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_U2 ( .A(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3829), .A2(n285), .ZN(
        stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n7), .ZN(
        stateArray_inS33ser[0]) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_3837), .A2(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_U1 ( .A1(
        stateArray_input_MC[0]), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3488) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3841), .A2(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3471), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n7), .ZN(
        stateArray_inS33ser[1]) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_3845), .A2(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_U1 ( .A1(
        stateArray_input_MC[1]), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3499) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3849), .A2(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3480), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n7), .ZN(
        stateArray_inS33ser[2]) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_3853), .A2(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_U1 ( .A1(
        stateArray_input_MC[2]), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3501) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3857), .A2(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3481), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n7), .ZN(
        stateArray_inS33ser[3]) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_3861), .A2(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_U1 ( .A1(
        stateArray_input_MC[3]), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3503) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3865), .A2(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3482), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n7), .ZN(
        stateArray_inS33ser[4]) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_3869), .A2(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_U1 ( .A1(
        stateArray_input_MC[4]), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3505) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3873), .A2(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3483), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n7), .ZN(
        stateArray_inS33ser[5]) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_3877), .A2(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_U1 ( .A1(
        stateArray_input_MC[5]), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3507) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3881), .A2(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3484), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n7), .ZN(
        stateArray_inS33ser[6]) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_3885), .A2(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_U1 ( .A1(
        stateArray_input_MC[6]), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3509) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3889), .A2(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3485), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n7), .ZN(
        stateArray_inS33ser[7]) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_3893), .A2(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_U1 ( .A1(
        stateArray_input_MC[7]), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_n8) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_U4 ( .A1(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n8), .A2(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3511) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_3897), .A2(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n6), .ZN(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n7) );
  INV_X1 stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_U2 ( .A(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n6) );
  NAND2_X1 stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3486), .A2(n284), .ZN(
        stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_n8) );
  XNOR2_X1 KeyArray_U42_Ins0_U1 ( .A(KeyArray_n55), .B(new_AGEMA_signal_3901),
        .ZN(KeyArray_inS30par[7]) );
  XOR2_X1 KeyArray_U42_Ins_1_U1 ( .A(new_AGEMA_signal_3472), .B(
        new_AGEMA_signal_3905), .Z(new_AGEMA_signal_3489) );
  XNOR2_X1 KeyArray_U41_Ins0_U1 ( .A(new_AGEMA_signal_3909), .B(SboxOut[7]),
        .ZN(KeyArray_n55) );
  XNOR2_X1 KeyArray_U40_Ins0_U1 ( .A(KeyArray_n54), .B(new_AGEMA_signal_3913),
        .ZN(KeyArray_inS30par[6]) );
  XOR2_X1 KeyArray_U40_Ins_1_U1 ( .A(new_AGEMA_signal_3473), .B(
        new_AGEMA_signal_3917), .Z(new_AGEMA_signal_3490) );
  XNOR2_X1 KeyArray_U39_Ins0_U1 ( .A(new_AGEMA_signal_3921), .B(SboxOut[6]),
        .ZN(KeyArray_n54) );
  XNOR2_X1 KeyArray_U38_Ins0_U1 ( .A(KeyArray_n53), .B(new_AGEMA_signal_3925),
        .ZN(KeyArray_inS30par[5]) );
  XOR2_X1 KeyArray_U38_Ins_1_U1 ( .A(new_AGEMA_signal_3474), .B(
        new_AGEMA_signal_3929), .Z(new_AGEMA_signal_3491) );
  XNOR2_X1 KeyArray_U37_Ins0_U1 ( .A(new_AGEMA_signal_3933), .B(SboxOut[5]),
        .ZN(KeyArray_n53) );
  XNOR2_X1 KeyArray_U36_Ins0_U1 ( .A(KeyArray_n52), .B(new_AGEMA_signal_3937),
        .ZN(KeyArray_inS30par[4]) );
  XOR2_X1 KeyArray_U36_Ins_1_U1 ( .A(new_AGEMA_signal_3475), .B(
        new_AGEMA_signal_3941), .Z(new_AGEMA_signal_3492) );
  XNOR2_X1 KeyArray_U35_Ins0_U1 ( .A(new_AGEMA_signal_3945), .B(SboxOut[4]),
        .ZN(KeyArray_n52) );
  XNOR2_X1 KeyArray_U34_Ins0_U1 ( .A(KeyArray_n51), .B(new_AGEMA_signal_3949),
        .ZN(KeyArray_inS30par[3]) );
  XOR2_X1 KeyArray_U34_Ins_1_U1 ( .A(new_AGEMA_signal_3476), .B(
        new_AGEMA_signal_3953), .Z(new_AGEMA_signal_3493) );
  XNOR2_X1 KeyArray_U33_Ins0_U1 ( .A(new_AGEMA_signal_3957), .B(SboxOut[3]),
        .ZN(KeyArray_n51) );
  XNOR2_X1 KeyArray_U32_Ins0_U1 ( .A(KeyArray_n50), .B(new_AGEMA_signal_3961),
        .ZN(KeyArray_inS30par[2]) );
  XOR2_X1 KeyArray_U32_Ins_1_U1 ( .A(new_AGEMA_signal_3477), .B(
        new_AGEMA_signal_3965), .Z(new_AGEMA_signal_3494) );
  XNOR2_X1 KeyArray_U31_Ins0_U1 ( .A(new_AGEMA_signal_3969), .B(SboxOut[2]),
        .ZN(KeyArray_n50) );
  XNOR2_X1 KeyArray_U30_Ins0_U1 ( .A(KeyArray_n49), .B(new_AGEMA_signal_3973),
        .ZN(KeyArray_inS30par[1]) );
  XOR2_X1 KeyArray_U30_Ins_1_U1 ( .A(new_AGEMA_signal_3478), .B(
        new_AGEMA_signal_3977), .Z(new_AGEMA_signal_3495) );
  XNOR2_X1 KeyArray_U29_Ins0_U1 ( .A(new_AGEMA_signal_3981), .B(SboxOut[1]),
        .ZN(KeyArray_n49) );
  XNOR2_X1 KeyArray_U28_Ins0_U1 ( .A(KeyArray_n48), .B(new_AGEMA_signal_3985),
        .ZN(KeyArray_inS30par[0]) );
  XOR2_X1 KeyArray_U28_Ins_1_U1 ( .A(new_AGEMA_signal_3456), .B(
        new_AGEMA_signal_3989), .Z(new_AGEMA_signal_3479) );
  XNOR2_X1 KeyArray_U27_Ins0_U1 ( .A(new_AGEMA_signal_3993), .B(SboxOut[0]),
        .ZN(KeyArray_n48) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_n5) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_U3 ( .A1(new_AGEMA_signal_4001), .A2(KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A1(
        KeyArray_S30reg_gff_1_SFF_0_QD), .A2(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3512)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_4005), .A2(KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3496), .A2(n283), .ZN(KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_QD) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_4013), .A2(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_inS30par[0]), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3496) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_4017), .A2(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3479), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_n5) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_U3 ( .A1(new_AGEMA_signal_4021), .A2(KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A1(
        KeyArray_S30reg_gff_1_SFF_1_QD), .A2(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3527)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_4025), .A2(KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3513), .A2(n283), .ZN(KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_QD) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_4029), .A2(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_inS30par[1]), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3513) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_4033), .A2(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3495), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_n5) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_U3 ( .A1(new_AGEMA_signal_4037), .A2(KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A1(
        KeyArray_S30reg_gff_1_SFF_2_QD), .A2(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3528)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_4041), .A2(KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3514), .A2(n283), .ZN(KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_QD) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_4045), .A2(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_inS30par[2]), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3514) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_4049), .A2(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3494), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_n5) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_U3 ( .A1(new_AGEMA_signal_4053), .A2(KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A1(
        KeyArray_S30reg_gff_1_SFF_3_QD), .A2(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3529)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_4057), .A2(KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3515), .A2(n283), .ZN(KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_QD) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_4061), .A2(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_inS30par[3]), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3515) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_4065), .A2(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3493), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_n5) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_U3 ( .A1(new_AGEMA_signal_4069), .A2(KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A1(
        KeyArray_S30reg_gff_1_SFF_4_QD), .A2(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3530)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_4073), .A2(KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3516), .A2(n283), .ZN(KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_QD) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_4077), .A2(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_inS30par[4]), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3516) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_4081), .A2(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3492), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_n5) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_U3 ( .A1(new_AGEMA_signal_4085), .A2(KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A1(
        KeyArray_S30reg_gff_1_SFF_5_QD), .A2(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3531)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_4089), .A2(KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3517), .A2(n283), .ZN(KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_QD) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_4093), .A2(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_inS30par[5]), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3517) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_4097), .A2(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3491), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_n5) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_U3 ( .A1(new_AGEMA_signal_4101), .A2(KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A1(
        KeyArray_S30reg_gff_1_SFF_6_QD), .A2(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3532)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_4105), .A2(KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3518), .A2(n283), .ZN(KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_QD) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_4109), .A2(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_inS30par[6]), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3518) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_4113), .A2(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3490), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_n5) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_U3 ( .A1(new_AGEMA_signal_4117), .A2(KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A1(
        KeyArray_S30reg_gff_1_SFF_7_QD), .A2(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_n7), .ZN(new_AGEMA_signal_3533)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_U3 ( .A1(new_AGEMA_signal_4121), .A2(KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_U2 ( .A(n283), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A1(new_AGEMA_signal_3519), .A2(n283), .ZN(KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_QD) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U3 ( .A1(
        new_AGEMA_signal_4125), .A2(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A1(
        KeyArray_inS30par[7]), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_n8) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U4 ( .A1(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8), .A2(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7), .ZN(
        new_AGEMA_signal_3519) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U3 ( .A1(
        new_AGEMA_signal_4129), .A2(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n7) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U2 ( .A(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n6) );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A1(
        new_AGEMA_signal_3489), .A2(n282), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_n8) );
  XOR2_X1 Inst_bSbox_AND_M46_U1_U16 ( .A(Fresh[32]), .B(
        Inst_bSbox_AND_M46_U1_n23), .Z(Inst_bSbox_AND_M46_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M46_U1_U15 ( .A1(new_AGEMA_signal_3404), .A2(
        Inst_bSbox_AND_M46_U1_n22), .ZN(Inst_bSbox_AND_M46_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M46_U1_U14 ( .A(Fresh[32]), .B(
        Inst_bSbox_AND_M46_U1_n21), .Z(Inst_bSbox_AND_M46_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M46_U1_U13 ( .A1(Inst_bSbox_M44), .A2(
        Inst_bSbox_AND_M46_U1_n22), .ZN(Inst_bSbox_AND_M46_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M46_U1_U12 ( .A(Inst_bSbox_AND_M46_U1_n20), .B(
        Inst_bSbox_AND_M46_U1_n19), .ZN(Inst_bSbox_M46) );
  NAND2_X1 Inst_bSbox_AND_M46_U1_U11 ( .A1(Inst_bSbox_AND_M46_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M46_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M46_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M46_U1_U10 ( .A(Inst_bSbox_AND_M46_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M46_U1_z[0]), .Z(Inst_bSbox_AND_M46_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M46_U1_U9 ( .A(Inst_bSbox_AND_M46_U1_n18), .B(
        Inst_bSbox_AND_M46_U1_n17), .ZN(new_AGEMA_signal_3414) );
  NAND2_X1 Inst_bSbox_AND_M46_U1_U8 ( .A1(Inst_bSbox_AND_M46_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M46_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M46_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M46_U1_U7 ( .A(Inst_bSbox_AND_M46_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M46_U1_z[1]), .Z(Inst_bSbox_AND_M46_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M46_U1_U6 ( .A(new_AGEMA_signal_4135), .B(
        Inst_bSbox_AND_M46_U1_n22), .ZN(Inst_bSbox_AND_M46_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M46_U1_U5 ( .A(new_AGEMA_signal_4132), .B(
        Inst_bSbox_AND_M46_U1_n22), .ZN(Inst_bSbox_AND_M46_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M46_U1_U4 ( .A(Fresh[33]), .ZN(
        Inst_bSbox_AND_M46_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M46_U1_U3 ( .A1(new_AGEMA_signal_3404), .A2(
        new_AGEMA_signal_4135), .ZN(Inst_bSbox_AND_M46_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M46_U1_U2 ( .A1(Inst_bSbox_M44), .A2(
        new_AGEMA_signal_4132), .ZN(Inst_bSbox_AND_M46_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M46_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M46_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M46_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M44),
        .CK(clk), .Q(Inst_bSbox_AND_M46_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M46_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M46_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M46_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M46_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M46_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M46_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M46_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3404), .CK(clk), .Q(Inst_bSbox_AND_M46_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M46_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M46_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M46_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M46_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M47_U1_U16 ( .A(Fresh[34]), .B(
        Inst_bSbox_AND_M47_U1_n23), .Z(Inst_bSbox_AND_M47_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M47_U1_U15 ( .A1(new_AGEMA_signal_3400), .A2(
        Inst_bSbox_AND_M47_U1_n22), .ZN(Inst_bSbox_AND_M47_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M47_U1_U14 ( .A(Fresh[34]), .B(
        Inst_bSbox_AND_M47_U1_n21), .Z(Inst_bSbox_AND_M47_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M47_U1_U13 ( .A1(Inst_bSbox_M40), .A2(
        Inst_bSbox_AND_M47_U1_n22), .ZN(Inst_bSbox_AND_M47_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M47_U1_U12 ( .A(Inst_bSbox_AND_M47_U1_n20), .B(
        Inst_bSbox_AND_M47_U1_n19), .ZN(Inst_bSbox_M47) );
  NAND2_X1 Inst_bSbox_AND_M47_U1_U11 ( .A1(Inst_bSbox_AND_M47_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M47_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M47_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M47_U1_U10 ( .A(Inst_bSbox_AND_M47_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M47_U1_z[0]), .Z(Inst_bSbox_AND_M47_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M47_U1_U9 ( .A(Inst_bSbox_AND_M47_U1_n18), .B(
        Inst_bSbox_AND_M47_U1_n17), .ZN(new_AGEMA_signal_3405) );
  NAND2_X1 Inst_bSbox_AND_M47_U1_U8 ( .A1(Inst_bSbox_AND_M47_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M47_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M47_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M47_U1_U7 ( .A(Inst_bSbox_AND_M47_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M47_U1_z[1]), .Z(Inst_bSbox_AND_M47_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M47_U1_U6 ( .A(new_AGEMA_signal_4141), .B(
        Inst_bSbox_AND_M47_U1_n22), .ZN(Inst_bSbox_AND_M47_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M47_U1_U5 ( .A(new_AGEMA_signal_4138), .B(
        Inst_bSbox_AND_M47_U1_n22), .ZN(Inst_bSbox_AND_M47_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M47_U1_U4 ( .A(Fresh[35]), .ZN(
        Inst_bSbox_AND_M47_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M47_U1_U3 ( .A1(Inst_bSbox_M40), .A2(
        new_AGEMA_signal_4138), .ZN(Inst_bSbox_AND_M47_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M47_U1_U2 ( .A1(new_AGEMA_signal_3400), .A2(
        new_AGEMA_signal_4141), .ZN(Inst_bSbox_AND_M47_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M47_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M47_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M47_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M40),
        .CK(clk), .Q(Inst_bSbox_AND_M47_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M47_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M47_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M47_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M47_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M47_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M47_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M47_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3400), .CK(clk), .Q(Inst_bSbox_AND_M47_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M47_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M47_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M47_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M47_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M48_U1_U16 ( .A(Fresh[36]), .B(
        Inst_bSbox_AND_M48_U1_n23), .Z(Inst_bSbox_AND_M48_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M48_U1_U15 ( .A1(new_AGEMA_signal_3399), .A2(
        Inst_bSbox_AND_M48_U1_n22), .ZN(Inst_bSbox_AND_M48_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M48_U1_U14 ( .A(Fresh[36]), .B(
        Inst_bSbox_AND_M48_U1_n21), .Z(Inst_bSbox_AND_M48_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M48_U1_U13 ( .A1(Inst_bSbox_M39), .A2(
        Inst_bSbox_AND_M48_U1_n22), .ZN(Inst_bSbox_AND_M48_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M48_U1_U12 ( .A(Inst_bSbox_AND_M48_U1_n20), .B(
        Inst_bSbox_AND_M48_U1_n19), .ZN(Inst_bSbox_M48) );
  NAND2_X1 Inst_bSbox_AND_M48_U1_U11 ( .A1(Inst_bSbox_AND_M48_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M48_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M48_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M48_U1_U10 ( .A(Inst_bSbox_AND_M48_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M48_U1_z[0]), .Z(Inst_bSbox_AND_M48_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M48_U1_U9 ( .A(Inst_bSbox_AND_M48_U1_n18), .B(
        Inst_bSbox_AND_M48_U1_n17), .ZN(new_AGEMA_signal_3406) );
  NAND2_X1 Inst_bSbox_AND_M48_U1_U8 ( .A1(Inst_bSbox_AND_M48_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M48_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M48_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M48_U1_U7 ( .A(Inst_bSbox_AND_M48_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M48_U1_z[1]), .Z(Inst_bSbox_AND_M48_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M48_U1_U6 ( .A(new_AGEMA_signal_4147), .B(
        Inst_bSbox_AND_M48_U1_n22), .ZN(Inst_bSbox_AND_M48_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M48_U1_U5 ( .A(new_AGEMA_signal_4144), .B(
        Inst_bSbox_AND_M48_U1_n22), .ZN(Inst_bSbox_AND_M48_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M48_U1_U4 ( .A(Fresh[37]), .ZN(
        Inst_bSbox_AND_M48_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M48_U1_U3 ( .A1(Inst_bSbox_M39), .A2(
        new_AGEMA_signal_4144), .ZN(Inst_bSbox_AND_M48_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M48_U1_U2 ( .A1(new_AGEMA_signal_3399), .A2(
        new_AGEMA_signal_4147), .ZN(Inst_bSbox_AND_M48_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M48_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M48_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M48_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M39),
        .CK(clk), .Q(Inst_bSbox_AND_M48_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M48_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M48_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M48_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M48_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M48_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M48_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M48_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3399), .CK(clk), .Q(Inst_bSbox_AND_M48_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M48_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M48_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M48_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M48_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M49_U1_U16 ( .A(Fresh[38]), .B(
        Inst_bSbox_AND_M49_U1_n23), .Z(Inst_bSbox_AND_M49_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M49_U1_U15 ( .A1(new_AGEMA_signal_3403), .A2(
        Inst_bSbox_AND_M49_U1_n22), .ZN(Inst_bSbox_AND_M49_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M49_U1_U14 ( .A(Fresh[38]), .B(
        Inst_bSbox_AND_M49_U1_n21), .Z(Inst_bSbox_AND_M49_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M49_U1_U13 ( .A1(Inst_bSbox_M43), .A2(
        Inst_bSbox_AND_M49_U1_n22), .ZN(Inst_bSbox_AND_M49_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M49_U1_U12 ( .A(Inst_bSbox_AND_M49_U1_n20), .B(
        Inst_bSbox_AND_M49_U1_n19), .ZN(Inst_bSbox_M49) );
  NAND2_X1 Inst_bSbox_AND_M49_U1_U11 ( .A1(Inst_bSbox_AND_M49_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M49_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M49_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M49_U1_U10 ( .A(Inst_bSbox_AND_M49_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M49_U1_z[0]), .Z(Inst_bSbox_AND_M49_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M49_U1_U9 ( .A(Inst_bSbox_AND_M49_U1_n18), .B(
        Inst_bSbox_AND_M49_U1_n17), .ZN(new_AGEMA_signal_3415) );
  NAND2_X1 Inst_bSbox_AND_M49_U1_U8 ( .A1(Inst_bSbox_AND_M49_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M49_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M49_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M49_U1_U7 ( .A(Inst_bSbox_AND_M49_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M49_U1_z[1]), .Z(Inst_bSbox_AND_M49_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M49_U1_U6 ( .A(new_AGEMA_signal_4153), .B(
        Inst_bSbox_AND_M49_U1_n22), .ZN(Inst_bSbox_AND_M49_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M49_U1_U5 ( .A(new_AGEMA_signal_4150), .B(
        Inst_bSbox_AND_M49_U1_n22), .ZN(Inst_bSbox_AND_M49_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M49_U1_U4 ( .A(Fresh[39]), .ZN(
        Inst_bSbox_AND_M49_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M49_U1_U3 ( .A1(Inst_bSbox_M43), .A2(
        new_AGEMA_signal_4150), .ZN(Inst_bSbox_AND_M49_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M49_U1_U2 ( .A1(new_AGEMA_signal_3403), .A2(
        new_AGEMA_signal_4153), .ZN(Inst_bSbox_AND_M49_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M49_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M49_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M49_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M43),
        .CK(clk), .Q(Inst_bSbox_AND_M49_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M49_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M49_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M49_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M49_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M49_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M49_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M49_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3403), .CK(clk), .Q(Inst_bSbox_AND_M49_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M49_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M49_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M49_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M49_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M50_U1_U16 ( .A(Fresh[40]), .B(
        Inst_bSbox_AND_M50_U1_n23), .Z(Inst_bSbox_AND_M50_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M50_U1_U15 ( .A1(new_AGEMA_signal_3398), .A2(
        Inst_bSbox_AND_M50_U1_n22), .ZN(Inst_bSbox_AND_M50_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M50_U1_U14 ( .A(Fresh[40]), .B(
        Inst_bSbox_AND_M50_U1_n21), .Z(Inst_bSbox_AND_M50_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M50_U1_U13 ( .A1(Inst_bSbox_M38), .A2(
        Inst_bSbox_AND_M50_U1_n22), .ZN(Inst_bSbox_AND_M50_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M50_U1_U12 ( .A(Inst_bSbox_AND_M50_U1_n20), .B(
        Inst_bSbox_AND_M50_U1_n19), .ZN(Inst_bSbox_M50) );
  NAND2_X1 Inst_bSbox_AND_M50_U1_U11 ( .A1(Inst_bSbox_AND_M50_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M50_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M50_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M50_U1_U10 ( .A(Inst_bSbox_AND_M50_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M50_U1_z[0]), .Z(Inst_bSbox_AND_M50_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M50_U1_U9 ( .A(Inst_bSbox_AND_M50_U1_n18), .B(
        Inst_bSbox_AND_M50_U1_n17), .ZN(new_AGEMA_signal_3407) );
  NAND2_X1 Inst_bSbox_AND_M50_U1_U8 ( .A1(Inst_bSbox_AND_M50_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M50_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M50_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M50_U1_U7 ( .A(Inst_bSbox_AND_M50_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M50_U1_z[1]), .Z(Inst_bSbox_AND_M50_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M50_U1_U6 ( .A(new_AGEMA_signal_4159), .B(
        Inst_bSbox_AND_M50_U1_n22), .ZN(Inst_bSbox_AND_M50_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M50_U1_U5 ( .A(new_AGEMA_signal_4156), .B(
        Inst_bSbox_AND_M50_U1_n22), .ZN(Inst_bSbox_AND_M50_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M50_U1_U4 ( .A(Fresh[41]), .ZN(
        Inst_bSbox_AND_M50_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M50_U1_U3 ( .A1(new_AGEMA_signal_3398), .A2(
        new_AGEMA_signal_4159), .ZN(Inst_bSbox_AND_M50_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M50_U1_U2 ( .A1(Inst_bSbox_M38), .A2(
        new_AGEMA_signal_4156), .ZN(Inst_bSbox_AND_M50_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M50_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M50_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M50_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M38),
        .CK(clk), .Q(Inst_bSbox_AND_M50_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M50_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M50_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M50_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M50_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M50_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M50_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M50_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3398), .CK(clk), .Q(Inst_bSbox_AND_M50_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M50_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M50_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M50_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M50_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M51_U1_U16 ( .A(Fresh[42]), .B(
        Inst_bSbox_AND_M51_U1_n23), .Z(Inst_bSbox_AND_M51_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M51_U1_U15 ( .A1(new_AGEMA_signal_3397), .A2(
        Inst_bSbox_AND_M51_U1_n22), .ZN(Inst_bSbox_AND_M51_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M51_U1_U14 ( .A(Fresh[42]), .B(
        Inst_bSbox_AND_M51_U1_n21), .Z(Inst_bSbox_AND_M51_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M51_U1_U13 ( .A1(Inst_bSbox_M37), .A2(
        Inst_bSbox_AND_M51_U1_n22), .ZN(Inst_bSbox_AND_M51_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M51_U1_U12 ( .A(Inst_bSbox_AND_M51_U1_n20), .B(
        Inst_bSbox_AND_M51_U1_n19), .ZN(Inst_bSbox_M51) );
  NAND2_X1 Inst_bSbox_AND_M51_U1_U11 ( .A1(Inst_bSbox_AND_M51_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M51_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M51_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M51_U1_U10 ( .A(Inst_bSbox_AND_M51_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M51_U1_z[0]), .Z(Inst_bSbox_AND_M51_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M51_U1_U9 ( .A(Inst_bSbox_AND_M51_U1_n18), .B(
        Inst_bSbox_AND_M51_U1_n17), .ZN(new_AGEMA_signal_3408) );
  NAND2_X1 Inst_bSbox_AND_M51_U1_U8 ( .A1(Inst_bSbox_AND_M51_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M51_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M51_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M51_U1_U7 ( .A(Inst_bSbox_AND_M51_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M51_U1_z[1]), .Z(Inst_bSbox_AND_M51_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M51_U1_U6 ( .A(new_AGEMA_signal_4165), .B(
        Inst_bSbox_AND_M51_U1_n22), .ZN(Inst_bSbox_AND_M51_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M51_U1_U5 ( .A(new_AGEMA_signal_4162), .B(
        Inst_bSbox_AND_M51_U1_n22), .ZN(Inst_bSbox_AND_M51_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M51_U1_U4 ( .A(Fresh[43]), .ZN(
        Inst_bSbox_AND_M51_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M51_U1_U3 ( .A1(Inst_bSbox_M37), .A2(
        new_AGEMA_signal_4162), .ZN(Inst_bSbox_AND_M51_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M51_U1_U2 ( .A1(new_AGEMA_signal_3397), .A2(
        new_AGEMA_signal_4165), .ZN(Inst_bSbox_AND_M51_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M51_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M51_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M51_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M37),
        .CK(clk), .Q(Inst_bSbox_AND_M51_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M51_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M51_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M51_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M51_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M51_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M51_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M51_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3397), .CK(clk), .Q(Inst_bSbox_AND_M51_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M51_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M51_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M51_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M51_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M52_U1_U16 ( .A(Fresh[44]), .B(
        Inst_bSbox_AND_M52_U1_n23), .Z(Inst_bSbox_AND_M52_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M52_U1_U15 ( .A1(new_AGEMA_signal_3402), .A2(
        Inst_bSbox_AND_M52_U1_n22), .ZN(Inst_bSbox_AND_M52_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M52_U1_U14 ( .A(Fresh[44]), .B(
        Inst_bSbox_AND_M52_U1_n21), .Z(Inst_bSbox_AND_M52_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M52_U1_U13 ( .A1(Inst_bSbox_M42), .A2(
        Inst_bSbox_AND_M52_U1_n22), .ZN(Inst_bSbox_AND_M52_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M52_U1_U12 ( .A(Inst_bSbox_AND_M52_U1_n20), .B(
        Inst_bSbox_AND_M52_U1_n19), .ZN(Inst_bSbox_M52) );
  NAND2_X1 Inst_bSbox_AND_M52_U1_U11 ( .A1(Inst_bSbox_AND_M52_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M52_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M52_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M52_U1_U10 ( .A(Inst_bSbox_AND_M52_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M52_U1_z[0]), .Z(Inst_bSbox_AND_M52_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M52_U1_U9 ( .A(Inst_bSbox_AND_M52_U1_n18), .B(
        Inst_bSbox_AND_M52_U1_n17), .ZN(new_AGEMA_signal_3416) );
  NAND2_X1 Inst_bSbox_AND_M52_U1_U8 ( .A1(Inst_bSbox_AND_M52_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M52_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M52_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M52_U1_U7 ( .A(Inst_bSbox_AND_M52_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M52_U1_z[1]), .Z(Inst_bSbox_AND_M52_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M52_U1_U6 ( .A(new_AGEMA_signal_4171), .B(
        Inst_bSbox_AND_M52_U1_n22), .ZN(Inst_bSbox_AND_M52_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M52_U1_U5 ( .A(new_AGEMA_signal_4168), .B(
        Inst_bSbox_AND_M52_U1_n22), .ZN(Inst_bSbox_AND_M52_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M52_U1_U4 ( .A(Fresh[45]), .ZN(
        Inst_bSbox_AND_M52_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M52_U1_U3 ( .A1(new_AGEMA_signal_3402), .A2(
        new_AGEMA_signal_4171), .ZN(Inst_bSbox_AND_M52_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M52_U1_U2 ( .A1(Inst_bSbox_M42), .A2(
        new_AGEMA_signal_4168), .ZN(Inst_bSbox_AND_M52_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M52_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M52_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M52_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M42),
        .CK(clk), .Q(Inst_bSbox_AND_M52_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M52_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M52_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M52_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M52_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M52_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M52_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M52_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3402), .CK(clk), .Q(Inst_bSbox_AND_M52_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M52_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M52_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M52_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M52_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M53_U1_U16 ( .A(Fresh[46]), .B(
        Inst_bSbox_AND_M53_U1_n23), .Z(Inst_bSbox_AND_M53_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M53_U1_U15 ( .A1(new_AGEMA_signal_3413), .A2(
        Inst_bSbox_AND_M53_U1_n22), .ZN(Inst_bSbox_AND_M53_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M53_U1_U14 ( .A(Fresh[46]), .B(
        Inst_bSbox_AND_M53_U1_n21), .Z(Inst_bSbox_AND_M53_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M53_U1_U13 ( .A1(Inst_bSbox_M45), .A2(
        Inst_bSbox_AND_M53_U1_n22), .ZN(Inst_bSbox_AND_M53_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M53_U1_U12 ( .A(Inst_bSbox_AND_M53_U1_n20), .B(
        Inst_bSbox_AND_M53_U1_n19), .ZN(Inst_bSbox_M53) );
  NAND2_X1 Inst_bSbox_AND_M53_U1_U11 ( .A1(Inst_bSbox_AND_M53_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M53_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M53_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M53_U1_U10 ( .A(Inst_bSbox_AND_M53_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M53_U1_z[0]), .Z(Inst_bSbox_AND_M53_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M53_U1_U9 ( .A(Inst_bSbox_AND_M53_U1_n18), .B(
        Inst_bSbox_AND_M53_U1_n17), .ZN(new_AGEMA_signal_3425) );
  NAND2_X1 Inst_bSbox_AND_M53_U1_U8 ( .A1(Inst_bSbox_AND_M53_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M53_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M53_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M53_U1_U7 ( .A(Inst_bSbox_AND_M53_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M53_U1_z[1]), .Z(Inst_bSbox_AND_M53_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M53_U1_U6 ( .A(new_AGEMA_signal_4177), .B(
        Inst_bSbox_AND_M53_U1_n22), .ZN(Inst_bSbox_AND_M53_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M53_U1_U5 ( .A(new_AGEMA_signal_4174), .B(
        Inst_bSbox_AND_M53_U1_n22), .ZN(Inst_bSbox_AND_M53_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M53_U1_U4 ( .A(Fresh[47]), .ZN(
        Inst_bSbox_AND_M53_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M53_U1_U3 ( .A1(new_AGEMA_signal_3413), .A2(
        new_AGEMA_signal_4177), .ZN(Inst_bSbox_AND_M53_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M53_U1_U2 ( .A1(Inst_bSbox_M45), .A2(
        new_AGEMA_signal_4174), .ZN(Inst_bSbox_AND_M53_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M53_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M53_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M53_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M45),
        .CK(clk), .Q(Inst_bSbox_AND_M53_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M53_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M53_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M53_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M53_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M53_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M53_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M53_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3413), .CK(clk), .Q(Inst_bSbox_AND_M53_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M53_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M53_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M53_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M53_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M54_U1_U16 ( .A(Fresh[48]), .B(
        Inst_bSbox_AND_M54_U1_n23), .Z(Inst_bSbox_AND_M54_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M54_U1_U15 ( .A1(new_AGEMA_signal_3401), .A2(
        Inst_bSbox_AND_M54_U1_n22), .ZN(Inst_bSbox_AND_M54_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M54_U1_U14 ( .A(Fresh[48]), .B(
        Inst_bSbox_AND_M54_U1_n21), .Z(Inst_bSbox_AND_M54_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M54_U1_U13 ( .A1(Inst_bSbox_M41), .A2(
        Inst_bSbox_AND_M54_U1_n22), .ZN(Inst_bSbox_AND_M54_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M54_U1_U12 ( .A(Inst_bSbox_AND_M54_U1_n20), .B(
        Inst_bSbox_AND_M54_U1_n19), .ZN(Inst_bSbox_M54) );
  NAND2_X1 Inst_bSbox_AND_M54_U1_U11 ( .A1(Inst_bSbox_AND_M54_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M54_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M54_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M54_U1_U10 ( .A(Inst_bSbox_AND_M54_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M54_U1_z[0]), .Z(Inst_bSbox_AND_M54_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M54_U1_U9 ( .A(Inst_bSbox_AND_M54_U1_n18), .B(
        Inst_bSbox_AND_M54_U1_n17), .ZN(new_AGEMA_signal_3417) );
  NAND2_X1 Inst_bSbox_AND_M54_U1_U8 ( .A1(Inst_bSbox_AND_M54_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M54_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M54_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M54_U1_U7 ( .A(Inst_bSbox_AND_M54_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M54_U1_z[1]), .Z(Inst_bSbox_AND_M54_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M54_U1_U6 ( .A(new_AGEMA_signal_4183), .B(
        Inst_bSbox_AND_M54_U1_n22), .ZN(Inst_bSbox_AND_M54_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M54_U1_U5 ( .A(new_AGEMA_signal_4180), .B(
        Inst_bSbox_AND_M54_U1_n22), .ZN(Inst_bSbox_AND_M54_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M54_U1_U4 ( .A(Fresh[49]), .ZN(
        Inst_bSbox_AND_M54_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M54_U1_U3 ( .A1(Inst_bSbox_M41), .A2(
        new_AGEMA_signal_4180), .ZN(Inst_bSbox_AND_M54_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M54_U1_U2 ( .A1(new_AGEMA_signal_3401), .A2(
        new_AGEMA_signal_4183), .ZN(Inst_bSbox_AND_M54_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M54_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M54_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M54_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M41),
        .CK(clk), .Q(Inst_bSbox_AND_M54_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M54_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M54_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M54_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M54_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M54_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M54_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M54_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3401), .CK(clk), .Q(Inst_bSbox_AND_M54_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M54_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M54_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M54_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M54_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M55_U1_U16 ( .A(Fresh[50]), .B(
        Inst_bSbox_AND_M55_U1_n23), .Z(Inst_bSbox_AND_M55_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M55_U1_U15 ( .A1(new_AGEMA_signal_3404), .A2(
        Inst_bSbox_AND_M55_U1_n22), .ZN(Inst_bSbox_AND_M55_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M55_U1_U14 ( .A(Fresh[50]), .B(
        Inst_bSbox_AND_M55_U1_n21), .Z(Inst_bSbox_AND_M55_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M55_U1_U13 ( .A1(Inst_bSbox_M44), .A2(
        Inst_bSbox_AND_M55_U1_n22), .ZN(Inst_bSbox_AND_M55_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M55_U1_U12 ( .A(Inst_bSbox_AND_M55_U1_n20), .B(
        Inst_bSbox_AND_M55_U1_n19), .ZN(Inst_bSbox_M55) );
  NAND2_X1 Inst_bSbox_AND_M55_U1_U11 ( .A1(Inst_bSbox_AND_M55_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M55_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M55_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M55_U1_U10 ( .A(Inst_bSbox_AND_M55_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M55_U1_z[0]), .Z(Inst_bSbox_AND_M55_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M55_U1_U9 ( .A(Inst_bSbox_AND_M55_U1_n18), .B(
        Inst_bSbox_AND_M55_U1_n17), .ZN(new_AGEMA_signal_3418) );
  NAND2_X1 Inst_bSbox_AND_M55_U1_U8 ( .A1(Inst_bSbox_AND_M55_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M55_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M55_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M55_U1_U7 ( .A(Inst_bSbox_AND_M55_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M55_U1_z[1]), .Z(Inst_bSbox_AND_M55_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M55_U1_U6 ( .A(new_AGEMA_signal_4189), .B(
        Inst_bSbox_AND_M55_U1_n22), .ZN(Inst_bSbox_AND_M55_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M55_U1_U5 ( .A(new_AGEMA_signal_4186), .B(
        Inst_bSbox_AND_M55_U1_n22), .ZN(Inst_bSbox_AND_M55_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M55_U1_U4 ( .A(Fresh[51]), .ZN(
        Inst_bSbox_AND_M55_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M55_U1_U3 ( .A1(Inst_bSbox_M44), .A2(
        new_AGEMA_signal_4186), .ZN(Inst_bSbox_AND_M55_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M55_U1_U2 ( .A1(new_AGEMA_signal_3404), .A2(
        new_AGEMA_signal_4189), .ZN(Inst_bSbox_AND_M55_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M55_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M55_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M55_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M44),
        .CK(clk), .Q(Inst_bSbox_AND_M55_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M55_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M55_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M55_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M55_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M55_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M55_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M55_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3404), .CK(clk), .Q(Inst_bSbox_AND_M55_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M55_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M55_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M55_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M55_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M56_U1_U16 ( .A(Fresh[52]), .B(
        Inst_bSbox_AND_M56_U1_n23), .Z(Inst_bSbox_AND_M56_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M56_U1_U15 ( .A1(new_AGEMA_signal_3400), .A2(
        Inst_bSbox_AND_M56_U1_n22), .ZN(Inst_bSbox_AND_M56_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M56_U1_U14 ( .A(Fresh[52]), .B(
        Inst_bSbox_AND_M56_U1_n21), .Z(Inst_bSbox_AND_M56_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M56_U1_U13 ( .A1(Inst_bSbox_M40), .A2(
        Inst_bSbox_AND_M56_U1_n22), .ZN(Inst_bSbox_AND_M56_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M56_U1_U12 ( .A(Inst_bSbox_AND_M56_U1_n20), .B(
        Inst_bSbox_AND_M56_U1_n19), .ZN(Inst_bSbox_M56) );
  NAND2_X1 Inst_bSbox_AND_M56_U1_U11 ( .A1(Inst_bSbox_AND_M56_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M56_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M56_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M56_U1_U10 ( .A(Inst_bSbox_AND_M56_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M56_U1_z[0]), .Z(Inst_bSbox_AND_M56_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M56_U1_U9 ( .A(Inst_bSbox_AND_M56_U1_n18), .B(
        Inst_bSbox_AND_M56_U1_n17), .ZN(new_AGEMA_signal_3409) );
  NAND2_X1 Inst_bSbox_AND_M56_U1_U8 ( .A1(Inst_bSbox_AND_M56_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M56_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M56_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M56_U1_U7 ( .A(Inst_bSbox_AND_M56_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M56_U1_z[1]), .Z(Inst_bSbox_AND_M56_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M56_U1_U6 ( .A(new_AGEMA_signal_4195), .B(
        Inst_bSbox_AND_M56_U1_n22), .ZN(Inst_bSbox_AND_M56_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M56_U1_U5 ( .A(new_AGEMA_signal_4192), .B(
        Inst_bSbox_AND_M56_U1_n22), .ZN(Inst_bSbox_AND_M56_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M56_U1_U4 ( .A(Fresh[53]), .ZN(
        Inst_bSbox_AND_M56_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M56_U1_U3 ( .A1(new_AGEMA_signal_3400), .A2(
        new_AGEMA_signal_4195), .ZN(Inst_bSbox_AND_M56_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M56_U1_U2 ( .A1(Inst_bSbox_M40), .A2(
        new_AGEMA_signal_4192), .ZN(Inst_bSbox_AND_M56_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M56_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M56_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M56_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M40),
        .CK(clk), .Q(Inst_bSbox_AND_M56_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M56_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M56_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M56_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M56_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M56_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M56_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M56_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3400), .CK(clk), .Q(Inst_bSbox_AND_M56_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M56_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M56_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M56_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M56_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M57_U1_U16 ( .A(Fresh[54]), .B(
        Inst_bSbox_AND_M57_U1_n23), .Z(Inst_bSbox_AND_M57_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M57_U1_U15 ( .A1(new_AGEMA_signal_3399), .A2(
        Inst_bSbox_AND_M57_U1_n22), .ZN(Inst_bSbox_AND_M57_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M57_U1_U14 ( .A(Fresh[54]), .B(
        Inst_bSbox_AND_M57_U1_n21), .Z(Inst_bSbox_AND_M57_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M57_U1_U13 ( .A1(Inst_bSbox_M39), .A2(
        Inst_bSbox_AND_M57_U1_n22), .ZN(Inst_bSbox_AND_M57_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M57_U1_U12 ( .A(Inst_bSbox_AND_M57_U1_n20), .B(
        Inst_bSbox_AND_M57_U1_n19), .ZN(Inst_bSbox_M57) );
  NAND2_X1 Inst_bSbox_AND_M57_U1_U11 ( .A1(Inst_bSbox_AND_M57_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M57_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M57_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M57_U1_U10 ( .A(Inst_bSbox_AND_M57_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M57_U1_z[0]), .Z(Inst_bSbox_AND_M57_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M57_U1_U9 ( .A(Inst_bSbox_AND_M57_U1_n18), .B(
        Inst_bSbox_AND_M57_U1_n17), .ZN(new_AGEMA_signal_3410) );
  NAND2_X1 Inst_bSbox_AND_M57_U1_U8 ( .A1(Inst_bSbox_AND_M57_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M57_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M57_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M57_U1_U7 ( .A(Inst_bSbox_AND_M57_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M57_U1_z[1]), .Z(Inst_bSbox_AND_M57_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M57_U1_U6 ( .A(new_AGEMA_signal_4201), .B(
        Inst_bSbox_AND_M57_U1_n22), .ZN(Inst_bSbox_AND_M57_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M57_U1_U5 ( .A(new_AGEMA_signal_4198), .B(
        Inst_bSbox_AND_M57_U1_n22), .ZN(Inst_bSbox_AND_M57_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M57_U1_U4 ( .A(Fresh[55]), .ZN(
        Inst_bSbox_AND_M57_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M57_U1_U3 ( .A1(new_AGEMA_signal_3399), .A2(
        new_AGEMA_signal_4201), .ZN(Inst_bSbox_AND_M57_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M57_U1_U2 ( .A1(Inst_bSbox_M39), .A2(
        new_AGEMA_signal_4198), .ZN(Inst_bSbox_AND_M57_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M57_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M57_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M57_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M39),
        .CK(clk), .Q(Inst_bSbox_AND_M57_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M57_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M57_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M57_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M57_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M57_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M57_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M57_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3399), .CK(clk), .Q(Inst_bSbox_AND_M57_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M57_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M57_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M57_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M57_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M58_U1_U16 ( .A(Fresh[56]), .B(
        Inst_bSbox_AND_M58_U1_n23), .Z(Inst_bSbox_AND_M58_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M58_U1_U15 ( .A1(new_AGEMA_signal_3403), .A2(
        Inst_bSbox_AND_M58_U1_n22), .ZN(Inst_bSbox_AND_M58_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M58_U1_U14 ( .A(Fresh[56]), .B(
        Inst_bSbox_AND_M58_U1_n21), .Z(Inst_bSbox_AND_M58_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M58_U1_U13 ( .A1(Inst_bSbox_M43), .A2(
        Inst_bSbox_AND_M58_U1_n22), .ZN(Inst_bSbox_AND_M58_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M58_U1_U12 ( .A(Inst_bSbox_AND_M58_U1_n20), .B(
        Inst_bSbox_AND_M58_U1_n19), .ZN(Inst_bSbox_M58) );
  NAND2_X1 Inst_bSbox_AND_M58_U1_U11 ( .A1(Inst_bSbox_AND_M58_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M58_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M58_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M58_U1_U10 ( .A(Inst_bSbox_AND_M58_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M58_U1_z[0]), .Z(Inst_bSbox_AND_M58_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M58_U1_U9 ( .A(Inst_bSbox_AND_M58_U1_n18), .B(
        Inst_bSbox_AND_M58_U1_n17), .ZN(new_AGEMA_signal_3419) );
  NAND2_X1 Inst_bSbox_AND_M58_U1_U8 ( .A1(Inst_bSbox_AND_M58_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M58_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M58_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M58_U1_U7 ( .A(Inst_bSbox_AND_M58_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M58_U1_z[1]), .Z(Inst_bSbox_AND_M58_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M58_U1_U6 ( .A(new_AGEMA_signal_4207), .B(
        Inst_bSbox_AND_M58_U1_n22), .ZN(Inst_bSbox_AND_M58_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M58_U1_U5 ( .A(new_AGEMA_signal_4204), .B(
        Inst_bSbox_AND_M58_U1_n22), .ZN(Inst_bSbox_AND_M58_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M58_U1_U4 ( .A(Fresh[57]), .ZN(
        Inst_bSbox_AND_M58_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M58_U1_U3 ( .A1(new_AGEMA_signal_3403), .A2(
        new_AGEMA_signal_4207), .ZN(Inst_bSbox_AND_M58_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M58_U1_U2 ( .A1(Inst_bSbox_M43), .A2(
        new_AGEMA_signal_4204), .ZN(Inst_bSbox_AND_M58_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M58_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M58_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M58_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M43),
        .CK(clk), .Q(Inst_bSbox_AND_M58_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M58_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M58_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M58_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M58_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M58_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M58_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M58_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3403), .CK(clk), .Q(Inst_bSbox_AND_M58_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M58_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M58_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M58_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M58_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M59_U1_U16 ( .A(Fresh[58]), .B(
        Inst_bSbox_AND_M59_U1_n23), .Z(Inst_bSbox_AND_M59_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M59_U1_U15 ( .A1(new_AGEMA_signal_3398), .A2(
        Inst_bSbox_AND_M59_U1_n22), .ZN(Inst_bSbox_AND_M59_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M59_U1_U14 ( .A(Fresh[58]), .B(
        Inst_bSbox_AND_M59_U1_n21), .Z(Inst_bSbox_AND_M59_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M59_U1_U13 ( .A1(Inst_bSbox_M38), .A2(
        Inst_bSbox_AND_M59_U1_n22), .ZN(Inst_bSbox_AND_M59_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M59_U1_U12 ( .A(Inst_bSbox_AND_M59_U1_n20), .B(
        Inst_bSbox_AND_M59_U1_n19), .ZN(Inst_bSbox_M59) );
  NAND2_X1 Inst_bSbox_AND_M59_U1_U11 ( .A1(Inst_bSbox_AND_M59_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M59_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M59_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M59_U1_U10 ( .A(Inst_bSbox_AND_M59_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M59_U1_z[0]), .Z(Inst_bSbox_AND_M59_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M59_U1_U9 ( .A(Inst_bSbox_AND_M59_U1_n18), .B(
        Inst_bSbox_AND_M59_U1_n17), .ZN(new_AGEMA_signal_3411) );
  NAND2_X1 Inst_bSbox_AND_M59_U1_U8 ( .A1(Inst_bSbox_AND_M59_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M59_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M59_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M59_U1_U7 ( .A(Inst_bSbox_AND_M59_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M59_U1_z[1]), .Z(Inst_bSbox_AND_M59_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M59_U1_U6 ( .A(new_AGEMA_signal_4213), .B(
        Inst_bSbox_AND_M59_U1_n22), .ZN(Inst_bSbox_AND_M59_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M59_U1_U5 ( .A(new_AGEMA_signal_4210), .B(
        Inst_bSbox_AND_M59_U1_n22), .ZN(Inst_bSbox_AND_M59_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M59_U1_U4 ( .A(Fresh[59]), .ZN(
        Inst_bSbox_AND_M59_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M59_U1_U3 ( .A1(Inst_bSbox_M38), .A2(
        new_AGEMA_signal_4210), .ZN(Inst_bSbox_AND_M59_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M59_U1_U2 ( .A1(new_AGEMA_signal_3398), .A2(
        new_AGEMA_signal_4213), .ZN(Inst_bSbox_AND_M59_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M59_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M59_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M59_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M38),
        .CK(clk), .Q(Inst_bSbox_AND_M59_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M59_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M59_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M59_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M59_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M59_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M59_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M59_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3398), .CK(clk), .Q(Inst_bSbox_AND_M59_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M59_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M59_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M59_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M59_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M60_U1_U16 ( .A(Fresh[60]), .B(
        Inst_bSbox_AND_M60_U1_n23), .Z(Inst_bSbox_AND_M60_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M60_U1_U15 ( .A1(new_AGEMA_signal_3397), .A2(
        Inst_bSbox_AND_M60_U1_n22), .ZN(Inst_bSbox_AND_M60_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M60_U1_U14 ( .A(Fresh[60]), .B(
        Inst_bSbox_AND_M60_U1_n21), .Z(Inst_bSbox_AND_M60_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M60_U1_U13 ( .A1(Inst_bSbox_M37), .A2(
        Inst_bSbox_AND_M60_U1_n22), .ZN(Inst_bSbox_AND_M60_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M60_U1_U12 ( .A(Inst_bSbox_AND_M60_U1_n20), .B(
        Inst_bSbox_AND_M60_U1_n19), .ZN(Inst_bSbox_M60) );
  NAND2_X1 Inst_bSbox_AND_M60_U1_U11 ( .A1(Inst_bSbox_AND_M60_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M60_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M60_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M60_U1_U10 ( .A(Inst_bSbox_AND_M60_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M60_U1_z[0]), .Z(Inst_bSbox_AND_M60_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M60_U1_U9 ( .A(Inst_bSbox_AND_M60_U1_n18), .B(
        Inst_bSbox_AND_M60_U1_n17), .ZN(new_AGEMA_signal_3412) );
  NAND2_X1 Inst_bSbox_AND_M60_U1_U8 ( .A1(Inst_bSbox_AND_M60_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M60_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M60_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M60_U1_U7 ( .A(Inst_bSbox_AND_M60_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M60_U1_z[1]), .Z(Inst_bSbox_AND_M60_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M60_U1_U6 ( .A(new_AGEMA_signal_4219), .B(
        Inst_bSbox_AND_M60_U1_n22), .ZN(Inst_bSbox_AND_M60_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M60_U1_U5 ( .A(new_AGEMA_signal_4216), .B(
        Inst_bSbox_AND_M60_U1_n22), .ZN(Inst_bSbox_AND_M60_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M60_U1_U4 ( .A(Fresh[61]), .ZN(
        Inst_bSbox_AND_M60_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M60_U1_U3 ( .A1(Inst_bSbox_M37), .A2(
        new_AGEMA_signal_4216), .ZN(Inst_bSbox_AND_M60_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M60_U1_U2 ( .A1(new_AGEMA_signal_3397), .A2(
        new_AGEMA_signal_4219), .ZN(Inst_bSbox_AND_M60_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M60_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M60_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M60_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M37),
        .CK(clk), .Q(Inst_bSbox_AND_M60_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M60_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M60_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M60_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M60_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M60_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M60_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M60_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3397), .CK(clk), .Q(Inst_bSbox_AND_M60_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M60_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M60_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M60_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M60_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M61_U1_U16 ( .A(Fresh[62]), .B(
        Inst_bSbox_AND_M61_U1_n23), .Z(Inst_bSbox_AND_M61_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M61_U1_U15 ( .A1(new_AGEMA_signal_3402), .A2(
        Inst_bSbox_AND_M61_U1_n22), .ZN(Inst_bSbox_AND_M61_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M61_U1_U14 ( .A(Fresh[62]), .B(
        Inst_bSbox_AND_M61_U1_n21), .Z(Inst_bSbox_AND_M61_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M61_U1_U13 ( .A1(Inst_bSbox_M42), .A2(
        Inst_bSbox_AND_M61_U1_n22), .ZN(Inst_bSbox_AND_M61_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M61_U1_U12 ( .A(Inst_bSbox_AND_M61_U1_n20), .B(
        Inst_bSbox_AND_M61_U1_n19), .ZN(Inst_bSbox_M61) );
  NAND2_X1 Inst_bSbox_AND_M61_U1_U11 ( .A1(Inst_bSbox_AND_M61_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M61_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M61_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M61_U1_U10 ( .A(Inst_bSbox_AND_M61_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M61_U1_z[0]), .Z(Inst_bSbox_AND_M61_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M61_U1_U9 ( .A(Inst_bSbox_AND_M61_U1_n18), .B(
        Inst_bSbox_AND_M61_U1_n17), .ZN(new_AGEMA_signal_3420) );
  NAND2_X1 Inst_bSbox_AND_M61_U1_U8 ( .A1(Inst_bSbox_AND_M61_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M61_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M61_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M61_U1_U7 ( .A(Inst_bSbox_AND_M61_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M61_U1_z[1]), .Z(Inst_bSbox_AND_M61_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M61_U1_U6 ( .A(new_AGEMA_signal_4225), .B(
        Inst_bSbox_AND_M61_U1_n22), .ZN(Inst_bSbox_AND_M61_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M61_U1_U5 ( .A(new_AGEMA_signal_4222), .B(
        Inst_bSbox_AND_M61_U1_n22), .ZN(Inst_bSbox_AND_M61_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M61_U1_U4 ( .A(Fresh[63]), .ZN(
        Inst_bSbox_AND_M61_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M61_U1_U3 ( .A1(Inst_bSbox_M42), .A2(
        new_AGEMA_signal_4222), .ZN(Inst_bSbox_AND_M61_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M61_U1_U2 ( .A1(new_AGEMA_signal_3402), .A2(
        new_AGEMA_signal_4225), .ZN(Inst_bSbox_AND_M61_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M61_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M61_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M61_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M42),
        .CK(clk), .Q(Inst_bSbox_AND_M61_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M61_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M61_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M61_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M61_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M61_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M61_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M61_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3402), .CK(clk), .Q(Inst_bSbox_AND_M61_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M61_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M61_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M61_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M61_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M62_U1_U16 ( .A(Fresh[64]), .B(
        Inst_bSbox_AND_M62_U1_n23), .Z(Inst_bSbox_AND_M62_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M62_U1_U15 ( .A1(new_AGEMA_signal_3413), .A2(
        Inst_bSbox_AND_M62_U1_n22), .ZN(Inst_bSbox_AND_M62_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M62_U1_U14 ( .A(Fresh[64]), .B(
        Inst_bSbox_AND_M62_U1_n21), .Z(Inst_bSbox_AND_M62_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M62_U1_U13 ( .A1(Inst_bSbox_M45), .A2(
        Inst_bSbox_AND_M62_U1_n22), .ZN(Inst_bSbox_AND_M62_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M62_U1_U12 ( .A(Inst_bSbox_AND_M62_U1_n20), .B(
        Inst_bSbox_AND_M62_U1_n19), .ZN(Inst_bSbox_M62) );
  NAND2_X1 Inst_bSbox_AND_M62_U1_U11 ( .A1(Inst_bSbox_AND_M62_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M62_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M62_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M62_U1_U10 ( .A(Inst_bSbox_AND_M62_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M62_U1_z[0]), .Z(Inst_bSbox_AND_M62_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M62_U1_U9 ( .A(Inst_bSbox_AND_M62_U1_n18), .B(
        Inst_bSbox_AND_M62_U1_n17), .ZN(new_AGEMA_signal_3426) );
  NAND2_X1 Inst_bSbox_AND_M62_U1_U8 ( .A1(Inst_bSbox_AND_M62_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M62_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M62_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M62_U1_U7 ( .A(Inst_bSbox_AND_M62_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M62_U1_z[1]), .Z(Inst_bSbox_AND_M62_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M62_U1_U6 ( .A(new_AGEMA_signal_4231), .B(
        Inst_bSbox_AND_M62_U1_n22), .ZN(Inst_bSbox_AND_M62_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M62_U1_U5 ( .A(new_AGEMA_signal_4228), .B(
        Inst_bSbox_AND_M62_U1_n22), .ZN(Inst_bSbox_AND_M62_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M62_U1_U4 ( .A(Fresh[65]), .ZN(
        Inst_bSbox_AND_M62_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M62_U1_U3 ( .A1(new_AGEMA_signal_3413), .A2(
        new_AGEMA_signal_4231), .ZN(Inst_bSbox_AND_M62_U1_mul[1]) );
  AND2_X1 Inst_bSbox_AND_M62_U1_U2 ( .A1(Inst_bSbox_M45), .A2(
        new_AGEMA_signal_4228), .ZN(Inst_bSbox_AND_M62_U1_mul[0]) );
  DFF_X1 Inst_bSbox_AND_M62_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M62_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M62_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M45),
        .CK(clk), .Q(Inst_bSbox_AND_M62_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M62_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M62_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M62_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M62_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M62_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M62_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M62_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3413), .CK(clk), .Q(Inst_bSbox_AND_M62_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M62_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M62_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M62_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M62_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_AND_M63_U1_U16 ( .A(Fresh[66]), .B(
        Inst_bSbox_AND_M63_U1_n23), .Z(Inst_bSbox_AND_M63_U1_p_0_in_1__0_) );
  NOR2_X1 Inst_bSbox_AND_M63_U1_U15 ( .A1(new_AGEMA_signal_3401), .A2(
        Inst_bSbox_AND_M63_U1_n22), .ZN(Inst_bSbox_AND_M63_U1_n23) );
  XOR2_X1 Inst_bSbox_AND_M63_U1_U14 ( .A(Fresh[66]), .B(
        Inst_bSbox_AND_M63_U1_n21), .Z(Inst_bSbox_AND_M63_U1_p_0_in_0__1_) );
  NOR2_X1 Inst_bSbox_AND_M63_U1_U13 ( .A1(Inst_bSbox_M41), .A2(
        Inst_bSbox_AND_M63_U1_n22), .ZN(Inst_bSbox_AND_M63_U1_n21) );
  XNOR2_X1 Inst_bSbox_AND_M63_U1_U12 ( .A(Inst_bSbox_AND_M63_U1_n20), .B(
        Inst_bSbox_AND_M63_U1_n19), .ZN(Inst_bSbox_M63) );
  NAND2_X1 Inst_bSbox_AND_M63_U1_U11 ( .A1(Inst_bSbox_AND_M63_U1_a_reg[0]),
        .A2(Inst_bSbox_AND_M63_U1_s_out_0__1_), .ZN(Inst_bSbox_AND_M63_U1_n19)
         );
  XOR2_X1 Inst_bSbox_AND_M63_U1_U10 ( .A(Inst_bSbox_AND_M63_U1_p_0_out_0__1_),
        .B(Inst_bSbox_AND_M63_U1_z[0]), .Z(Inst_bSbox_AND_M63_U1_n20) );
  XNOR2_X1 Inst_bSbox_AND_M63_U1_U9 ( .A(Inst_bSbox_AND_M63_U1_n18), .B(
        Inst_bSbox_AND_M63_U1_n17), .ZN(new_AGEMA_signal_3421) );
  NAND2_X1 Inst_bSbox_AND_M63_U1_U8 ( .A1(Inst_bSbox_AND_M63_U1_a_reg[1]),
        .A2(Inst_bSbox_AND_M63_U1_s_out_1__0_), .ZN(Inst_bSbox_AND_M63_U1_n17)
         );
  XOR2_X1 Inst_bSbox_AND_M63_U1_U7 ( .A(Inst_bSbox_AND_M63_U1_p_0_out_1__0_),
        .B(Inst_bSbox_AND_M63_U1_z[1]), .Z(Inst_bSbox_AND_M63_U1_n18) );
  XNOR2_X1 Inst_bSbox_AND_M63_U1_U6 ( .A(new_AGEMA_signal_4237), .B(
        Inst_bSbox_AND_M63_U1_n22), .ZN(Inst_bSbox_AND_M63_U1_s_in_0__1_) );
  XNOR2_X1 Inst_bSbox_AND_M63_U1_U5 ( .A(new_AGEMA_signal_4234), .B(
        Inst_bSbox_AND_M63_U1_n22), .ZN(Inst_bSbox_AND_M63_U1_s_in_1__0_) );
  INV_X1 Inst_bSbox_AND_M63_U1_U4 ( .A(Fresh[67]), .ZN(
        Inst_bSbox_AND_M63_U1_n22) );
  AND2_X1 Inst_bSbox_AND_M63_U1_U3 ( .A1(Inst_bSbox_M41), .A2(
        new_AGEMA_signal_4234), .ZN(Inst_bSbox_AND_M63_U1_mul[0]) );
  AND2_X1 Inst_bSbox_AND_M63_U1_U2 ( .A1(new_AGEMA_signal_3401), .A2(
        new_AGEMA_signal_4237), .ZN(Inst_bSbox_AND_M63_U1_mul[1]) );
  DFF_X1 Inst_bSbox_AND_M63_U1_mul_pipe_s1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_mul[0]), .CK(clk), .Q(Inst_bSbox_AND_M63_U1_z[0]) );
  DFF_X1 Inst_bSbox_AND_M63_U1_a_i_0_s_current_state_reg ( .D(Inst_bSbox_M41),
        .CK(clk), .Q(Inst_bSbox_AND_M63_U1_a_reg[0]) );
  DFF_X1 Inst_bSbox_AND_M63_U1_s_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_s_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M63_U1_s_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M63_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_p_0_in_0__1_), .CK(clk), .Q(
        Inst_bSbox_AND_M63_U1_p_0_out_0__1_) );
  DFF_X1 Inst_bSbox_AND_M63_U1_mul_pipe_s1_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_mul[1]), .CK(clk), .Q(Inst_bSbox_AND_M63_U1_z[1]) );
  DFF_X1 Inst_bSbox_AND_M63_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3401), .CK(clk), .Q(Inst_bSbox_AND_M63_U1_a_reg[1])
         );
  DFF_X1 Inst_bSbox_AND_M63_U1_s_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_s_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M63_U1_s_out_1__0_) );
  DFF_X1 Inst_bSbox_AND_M63_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_p_0_in_1__0_), .CK(clk), .Q(
        Inst_bSbox_AND_M63_U1_p_0_out_1__0_) );
  XOR2_X1 Inst_bSbox_XOR_L0_U1_Ins_0_U1 ( .A(Inst_bSbox_M61), .B(
        Inst_bSbox_M62), .Z(Inst_bSbox_L0) );
  XOR2_X1 Inst_bSbox_XOR_L0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3420), .B(
        new_AGEMA_signal_3426), .Z(new_AGEMA_signal_3435) );
  XOR2_X1 Inst_bSbox_XOR_L1_U1_Ins_0_U1 ( .A(Inst_bSbox_M50), .B(
        Inst_bSbox_M56), .Z(Inst_bSbox_L1) );
  XOR2_X1 Inst_bSbox_XOR_L1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3407), .B(
        new_AGEMA_signal_3409), .Z(new_AGEMA_signal_3422) );
  XOR2_X1 Inst_bSbox_XOR_L2_U1_Ins_0_U1 ( .A(Inst_bSbox_M46), .B(
        Inst_bSbox_M48), .Z(Inst_bSbox_L2) );
  XOR2_X1 Inst_bSbox_XOR_L2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3414), .B(
        new_AGEMA_signal_3406), .Z(new_AGEMA_signal_3427) );
  XOR2_X1 Inst_bSbox_XOR_L3_U1_Ins_0_U1 ( .A(Inst_bSbox_M47), .B(
        Inst_bSbox_M55), .Z(Inst_bSbox_L3) );
  XOR2_X1 Inst_bSbox_XOR_L3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3405), .B(
        new_AGEMA_signal_3418), .Z(new_AGEMA_signal_3428) );
  XOR2_X1 Inst_bSbox_XOR_L4_U1_Ins_0_U1 ( .A(Inst_bSbox_M54), .B(
        Inst_bSbox_M58), .Z(Inst_bSbox_L4) );
  XOR2_X1 Inst_bSbox_XOR_L4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3417), .B(
        new_AGEMA_signal_3419), .Z(new_AGEMA_signal_3429) );
  XOR2_X1 Inst_bSbox_XOR_L5_U1_Ins_0_U1 ( .A(Inst_bSbox_M49), .B(
        Inst_bSbox_M61), .Z(Inst_bSbox_L5) );
  XOR2_X1 Inst_bSbox_XOR_L5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3415), .B(
        new_AGEMA_signal_3420), .Z(new_AGEMA_signal_3430) );
  XOR2_X1 Inst_bSbox_XOR_L6_U1_Ins_0_U1 ( .A(Inst_bSbox_M62), .B(Inst_bSbox_L5), .Z(Inst_bSbox_L6) );
  XOR2_X1 Inst_bSbox_XOR_L6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3426), .B(
        new_AGEMA_signal_3430), .Z(new_AGEMA_signal_3436) );
  XOR2_X1 Inst_bSbox_XOR_L7_U1_Ins_0_U1 ( .A(Inst_bSbox_M46), .B(Inst_bSbox_L3), .Z(Inst_bSbox_L7) );
  XOR2_X1 Inst_bSbox_XOR_L7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3414), .B(
        new_AGEMA_signal_3428), .Z(new_AGEMA_signal_3437) );
  XOR2_X1 Inst_bSbox_XOR_L8_U1_Ins_0_U1 ( .A(Inst_bSbox_M51), .B(
        Inst_bSbox_M59), .Z(Inst_bSbox_L8) );
  XOR2_X1 Inst_bSbox_XOR_L8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3408), .B(
        new_AGEMA_signal_3411), .Z(new_AGEMA_signal_3423) );
  XOR2_X1 Inst_bSbox_XOR_L9_U1_Ins_0_U1 ( .A(Inst_bSbox_M52), .B(
        Inst_bSbox_M53), .Z(Inst_bSbox_L9) );
  XOR2_X1 Inst_bSbox_XOR_L9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3416), .B(
        new_AGEMA_signal_3425), .Z(new_AGEMA_signal_3438) );
  XOR2_X1 Inst_bSbox_XOR_L10_U1_Ins_0_U1 ( .A(Inst_bSbox_M53), .B(
        Inst_bSbox_L4), .Z(Inst_bSbox_L10) );
  XOR2_X1 Inst_bSbox_XOR_L10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3425), .B(
        new_AGEMA_signal_3429), .Z(new_AGEMA_signal_3439) );
  XOR2_X1 Inst_bSbox_XOR_L11_U1_Ins_0_U1 ( .A(Inst_bSbox_M60), .B(
        Inst_bSbox_L2), .Z(Inst_bSbox_L11) );
  XOR2_X1 Inst_bSbox_XOR_L11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3412), .B(
        new_AGEMA_signal_3427), .Z(new_AGEMA_signal_3440) );
  XOR2_X1 Inst_bSbox_XOR_L12_U1_Ins_0_U1 ( .A(Inst_bSbox_M48), .B(
        Inst_bSbox_M51), .Z(Inst_bSbox_L12) );
  XOR2_X1 Inst_bSbox_XOR_L12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3406), .B(
        new_AGEMA_signal_3408), .Z(new_AGEMA_signal_3424) );
  XOR2_X1 Inst_bSbox_XOR_L13_U1_Ins_0_U1 ( .A(Inst_bSbox_M50), .B(
        Inst_bSbox_L0), .Z(Inst_bSbox_L13) );
  XOR2_X1 Inst_bSbox_XOR_L13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3407), .B(
        new_AGEMA_signal_3435), .Z(new_AGEMA_signal_3444) );
  XOR2_X1 Inst_bSbox_XOR_L14_U1_Ins_0_U1 ( .A(Inst_bSbox_M52), .B(
        Inst_bSbox_M61), .Z(Inst_bSbox_L14) );
  XOR2_X1 Inst_bSbox_XOR_L14_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3416), .B(
        new_AGEMA_signal_3420), .Z(new_AGEMA_signal_3431) );
  XOR2_X1 Inst_bSbox_XOR_L15_U1_Ins_0_U1 ( .A(Inst_bSbox_M55), .B(
        Inst_bSbox_L1), .Z(Inst_bSbox_L15) );
  XOR2_X1 Inst_bSbox_XOR_L15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3418), .B(
        new_AGEMA_signal_3422), .Z(new_AGEMA_signal_3432) );
  XOR2_X1 Inst_bSbox_XOR_L16_U1_Ins_0_U1 ( .A(Inst_bSbox_M56), .B(
        Inst_bSbox_L0), .Z(Inst_bSbox_L16) );
  XOR2_X1 Inst_bSbox_XOR_L16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3409), .B(
        new_AGEMA_signal_3435), .Z(new_AGEMA_signal_3445) );
  XOR2_X1 Inst_bSbox_XOR_L17_U1_Ins_0_U1 ( .A(Inst_bSbox_M57), .B(
        Inst_bSbox_L1), .Z(Inst_bSbox_L17) );
  XOR2_X1 Inst_bSbox_XOR_L17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3410), .B(
        new_AGEMA_signal_3422), .Z(new_AGEMA_signal_3433) );
  XOR2_X1 Inst_bSbox_XOR_L18_U1_Ins_0_U1 ( .A(Inst_bSbox_M58), .B(
        Inst_bSbox_L8), .Z(Inst_bSbox_L18) );
  XOR2_X1 Inst_bSbox_XOR_L18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3419), .B(
        new_AGEMA_signal_3423), .Z(new_AGEMA_signal_3434) );
  XOR2_X1 Inst_bSbox_XOR_L19_U1_Ins_0_U1 ( .A(Inst_bSbox_M63), .B(
        Inst_bSbox_L4), .Z(Inst_bSbox_L19) );
  XOR2_X1 Inst_bSbox_XOR_L19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3421), .B(
        new_AGEMA_signal_3429), .Z(new_AGEMA_signal_3441) );
  XOR2_X1 Inst_bSbox_XOR_L20_U1_Ins_0_U1 ( .A(Inst_bSbox_L0), .B(Inst_bSbox_L1), .Z(Inst_bSbox_L20) );
  XOR2_X1 Inst_bSbox_XOR_L20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3435), .B(
        new_AGEMA_signal_3422), .Z(new_AGEMA_signal_3446) );
  XOR2_X1 Inst_bSbox_XOR_L21_U1_Ins_0_U1 ( .A(Inst_bSbox_L1), .B(Inst_bSbox_L7), .Z(Inst_bSbox_L21) );
  XOR2_X1 Inst_bSbox_XOR_L21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3422), .B(
        new_AGEMA_signal_3437), .Z(new_AGEMA_signal_3447) );
  XOR2_X1 Inst_bSbox_XOR_L22_U1_Ins_0_U1 ( .A(Inst_bSbox_L3), .B(
        Inst_bSbox_L12), .Z(Inst_bSbox_L22) );
  XOR2_X1 Inst_bSbox_XOR_L22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3428), .B(
        new_AGEMA_signal_3424), .Z(new_AGEMA_signal_3442) );
  XOR2_X1 Inst_bSbox_XOR_L23_U1_Ins_0_U1 ( .A(Inst_bSbox_L18), .B(
        Inst_bSbox_L2), .Z(Inst_bSbox_L23) );
  XOR2_X1 Inst_bSbox_XOR_L23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3434), .B(
        new_AGEMA_signal_3427), .Z(new_AGEMA_signal_3443) );
  XOR2_X1 Inst_bSbox_XOR_L24_U1_Ins_0_U1 ( .A(Inst_bSbox_L15), .B(
        Inst_bSbox_L9), .Z(Inst_bSbox_L24) );
  XOR2_X1 Inst_bSbox_XOR_L24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3432), .B(
        new_AGEMA_signal_3438), .Z(new_AGEMA_signal_3448) );
  XOR2_X1 Inst_bSbox_XOR_L25_U1_Ins_0_U1 ( .A(Inst_bSbox_L6), .B(
        Inst_bSbox_L10), .Z(Inst_bSbox_L25) );
  XOR2_X1 Inst_bSbox_XOR_L25_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3436), .B(
        new_AGEMA_signal_3439), .Z(new_AGEMA_signal_3449) );
  XOR2_X1 Inst_bSbox_XOR_L26_U1_Ins_0_U1 ( .A(Inst_bSbox_L7), .B(Inst_bSbox_L9), .Z(Inst_bSbox_L26) );
  XOR2_X1 Inst_bSbox_XOR_L26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3437), .B(
        new_AGEMA_signal_3438), .Z(new_AGEMA_signal_3450) );
  XOR2_X1 Inst_bSbox_XOR_L27_U1_Ins_0_U1 ( .A(Inst_bSbox_L8), .B(
        Inst_bSbox_L10), .Z(Inst_bSbox_L27) );
  XOR2_X1 Inst_bSbox_XOR_L27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3423), .B(
        new_AGEMA_signal_3439), .Z(new_AGEMA_signal_3451) );
  XOR2_X1 Inst_bSbox_XOR_L28_U1_Ins_0_U1 ( .A(Inst_bSbox_L11), .B(
        Inst_bSbox_L14), .Z(Inst_bSbox_L28) );
  XOR2_X1 Inst_bSbox_XOR_L28_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3440), .B(
        new_AGEMA_signal_3431), .Z(new_AGEMA_signal_3452) );
  XOR2_X1 Inst_bSbox_XOR_L29_U1_Ins_0_U1 ( .A(Inst_bSbox_L11), .B(
        Inst_bSbox_L17), .Z(Inst_bSbox_L29) );
  XOR2_X1 Inst_bSbox_XOR_L29_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3440), .B(
        new_AGEMA_signal_3433), .Z(new_AGEMA_signal_3453) );
  XOR2_X1 Inst_bSbox_XOR_S0_U1_Ins_0_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L24), .Z(SboxOut[7]) );
  XOR2_X1 Inst_bSbox_XOR_S0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3436), .B(
        new_AGEMA_signal_3448), .Z(new_AGEMA_signal_3472) );
  XNOR2_X1 Inst_bSbox_XOR_S1_U1_Ins0_U1 ( .A(Inst_bSbox_L16), .B(
        Inst_bSbox_L26), .ZN(SboxOut[6]) );
  XOR2_X1 Inst_bSbox_XOR_S1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3445), .B(
        new_AGEMA_signal_3450), .Z(new_AGEMA_signal_3473) );
  XNOR2_X1 Inst_bSbox_XOR_S2_U1_Ins0_U1 ( .A(Inst_bSbox_L19), .B(
        Inst_bSbox_L28), .ZN(SboxOut[5]) );
  XOR2_X1 Inst_bSbox_XOR_S2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3441), .B(
        new_AGEMA_signal_3452), .Z(new_AGEMA_signal_3474) );
  XOR2_X1 Inst_bSbox_XOR_S3_U1_Ins_0_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L21), .Z(SboxOut[4]) );
  XOR2_X1 Inst_bSbox_XOR_S3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3436), .B(
        new_AGEMA_signal_3447), .Z(new_AGEMA_signal_3475) );
  XOR2_X1 Inst_bSbox_XOR_S4_U1_Ins_0_U1 ( .A(Inst_bSbox_L20), .B(
        Inst_bSbox_L22), .Z(SboxOut[3]) );
  XOR2_X1 Inst_bSbox_XOR_S4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3446), .B(
        new_AGEMA_signal_3442), .Z(new_AGEMA_signal_3476) );
  XOR2_X1 Inst_bSbox_XOR_S5_U1_Ins_0_U1 ( .A(Inst_bSbox_L25), .B(
        Inst_bSbox_L29), .Z(SboxOut[2]) );
  XOR2_X1 Inst_bSbox_XOR_S5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3449), .B(
        new_AGEMA_signal_3453), .Z(new_AGEMA_signal_3477) );
  XNOR2_X1 Inst_bSbox_XOR_S6_U1_Ins0_U1 ( .A(Inst_bSbox_L13), .B(
        Inst_bSbox_L27), .ZN(SboxOut[1]) );
  XOR2_X1 Inst_bSbox_XOR_S6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3444), .B(
        new_AGEMA_signal_3451), .Z(new_AGEMA_signal_3478) );
  XNOR2_X1 Inst_bSbox_XOR_S7_U1_Ins0_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L23), .ZN(SboxOut[0]) );
  XOR2_X1 Inst_bSbox_XOR_S7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3436), .B(
        new_AGEMA_signal_3443), .Z(new_AGEMA_signal_3456) );
  DFF_X1 new_AGEMA_reg_buffer_1741_s_current_state_reg ( .D(
        new_AGEMA_signal_3628), .CK(clk), .Q(new_AGEMA_signal_3629) );
  DFF_X1 new_AGEMA_reg_buffer_1745_s_current_state_reg ( .D(
        new_AGEMA_signal_3632), .CK(clk), .Q(new_AGEMA_signal_3633) );
  DFF_X1 new_AGEMA_reg_buffer_1749_s_current_state_reg ( .D(
        new_AGEMA_signal_3636), .CK(clk), .Q(new_AGEMA_signal_3637) );
  DFF_X1 new_AGEMA_reg_buffer_1753_s_current_state_reg ( .D(
        new_AGEMA_signal_3640), .CK(clk), .Q(new_AGEMA_signal_3641) );
  DFF_X1 new_AGEMA_reg_buffer_1757_s_current_state_reg ( .D(
        new_AGEMA_signal_3644), .CK(clk), .Q(new_AGEMA_signal_3645) );
  DFF_X1 new_AGEMA_reg_buffer_1761_s_current_state_reg ( .D(
        new_AGEMA_signal_3648), .CK(clk), .Q(new_AGEMA_signal_3649) );
  DFF_X1 new_AGEMA_reg_buffer_1765_s_current_state_reg ( .D(
        new_AGEMA_signal_3652), .CK(clk), .Q(new_AGEMA_signal_3653) );
  DFF_X1 new_AGEMA_reg_buffer_1769_s_current_state_reg ( .D(
        new_AGEMA_signal_3656), .CK(clk), .Q(new_AGEMA_signal_3657) );
  DFF_X1 new_AGEMA_reg_buffer_1773_s_current_state_reg ( .D(
        new_AGEMA_signal_3660), .CK(clk), .Q(new_AGEMA_signal_3661) );
  DFF_X1 new_AGEMA_reg_buffer_1777_s_current_state_reg ( .D(
        new_AGEMA_signal_3664), .CK(clk), .Q(new_AGEMA_signal_3665) );
  DFF_X1 new_AGEMA_reg_buffer_1781_s_current_state_reg ( .D(
        new_AGEMA_signal_3668), .CK(clk), .Q(new_AGEMA_signal_3669) );
  DFF_X1 new_AGEMA_reg_buffer_1785_s_current_state_reg ( .D(
        new_AGEMA_signal_3672), .CK(clk), .Q(new_AGEMA_signal_3673) );
  DFF_X1 new_AGEMA_reg_buffer_1789_s_current_state_reg ( .D(
        new_AGEMA_signal_3676), .CK(clk), .Q(new_AGEMA_signal_3677) );
  DFF_X1 new_AGEMA_reg_buffer_1793_s_current_state_reg ( .D(
        new_AGEMA_signal_3680), .CK(clk), .Q(new_AGEMA_signal_3681) );
  DFF_X1 new_AGEMA_reg_buffer_1797_s_current_state_reg ( .D(
        new_AGEMA_signal_3684), .CK(clk), .Q(new_AGEMA_signal_3685) );
  DFF_X1 new_AGEMA_reg_buffer_1801_s_current_state_reg ( .D(
        new_AGEMA_signal_3688), .CK(clk), .Q(new_AGEMA_signal_3689) );
  DFF_X1 new_AGEMA_reg_buffer_1805_s_current_state_reg ( .D(
        new_AGEMA_signal_3692), .CK(clk), .Q(new_AGEMA_signal_3693) );
  DFF_X1 new_AGEMA_reg_buffer_1809_s_current_state_reg ( .D(
        new_AGEMA_signal_3696), .CK(clk), .Q(new_AGEMA_signal_3697) );
  DFF_X1 new_AGEMA_reg_buffer_1813_s_current_state_reg ( .D(
        new_AGEMA_signal_3700), .CK(clk), .Q(new_AGEMA_signal_3701) );
  DFF_X1 new_AGEMA_reg_buffer_1817_s_current_state_reg ( .D(
        new_AGEMA_signal_3704), .CK(clk), .Q(new_AGEMA_signal_3705) );
  DFF_X1 new_AGEMA_reg_buffer_1821_s_current_state_reg ( .D(
        new_AGEMA_signal_3708), .CK(clk), .Q(new_AGEMA_signal_3709) );
  DFF_X1 new_AGEMA_reg_buffer_1825_s_current_state_reg ( .D(
        new_AGEMA_signal_3712), .CK(clk), .Q(new_AGEMA_signal_3713) );
  DFF_X1 new_AGEMA_reg_buffer_1829_s_current_state_reg ( .D(
        new_AGEMA_signal_3716), .CK(clk), .Q(new_AGEMA_signal_3717) );
  DFF_X1 new_AGEMA_reg_buffer_1833_s_current_state_reg ( .D(
        new_AGEMA_signal_3720), .CK(clk), .Q(new_AGEMA_signal_3721) );
  DFF_X1 new_AGEMA_reg_buffer_1837_s_current_state_reg ( .D(
        new_AGEMA_signal_3724), .CK(clk), .Q(new_AGEMA_signal_3725) );
  DFF_X1 new_AGEMA_reg_buffer_1841_s_current_state_reg ( .D(
        new_AGEMA_signal_3728), .CK(clk), .Q(new_AGEMA_signal_3729) );
  DFF_X1 new_AGEMA_reg_buffer_1845_s_current_state_reg ( .D(
        new_AGEMA_signal_3732), .CK(clk), .Q(new_AGEMA_signal_3733) );
  DFF_X1 new_AGEMA_reg_buffer_1849_s_current_state_reg ( .D(
        new_AGEMA_signal_3736), .CK(clk), .Q(new_AGEMA_signal_3737) );
  DFF_X1 new_AGEMA_reg_buffer_1853_s_current_state_reg ( .D(
        new_AGEMA_signal_3740), .CK(clk), .Q(new_AGEMA_signal_3741) );
  DFF_X1 new_AGEMA_reg_buffer_1857_s_current_state_reg ( .D(
        new_AGEMA_signal_3744), .CK(clk), .Q(new_AGEMA_signal_3745) );
  DFF_X1 new_AGEMA_reg_buffer_1861_s_current_state_reg ( .D(
        new_AGEMA_signal_3748), .CK(clk), .Q(new_AGEMA_signal_3749) );
  DFF_X1 new_AGEMA_reg_buffer_1865_s_current_state_reg ( .D(
        new_AGEMA_signal_3752), .CK(clk), .Q(new_AGEMA_signal_3753) );
  DFF_X1 new_AGEMA_reg_buffer_1869_s_current_state_reg ( .D(
        new_AGEMA_signal_3756), .CK(clk), .Q(new_AGEMA_signal_3757) );
  DFF_X1 new_AGEMA_reg_buffer_1873_s_current_state_reg ( .D(
        new_AGEMA_signal_3760), .CK(clk), .Q(new_AGEMA_signal_3761) );
  DFF_X1 new_AGEMA_reg_buffer_1877_s_current_state_reg ( .D(
        new_AGEMA_signal_3764), .CK(clk), .Q(new_AGEMA_signal_3765) );
  DFF_X1 new_AGEMA_reg_buffer_1881_s_current_state_reg ( .D(
        new_AGEMA_signal_3768), .CK(clk), .Q(new_AGEMA_signal_3769) );
  DFF_X1 new_AGEMA_reg_buffer_1885_s_current_state_reg ( .D(
        new_AGEMA_signal_3772), .CK(clk), .Q(new_AGEMA_signal_3773) );
  DFF_X1 new_AGEMA_reg_buffer_1889_s_current_state_reg ( .D(
        new_AGEMA_signal_3776), .CK(clk), .Q(new_AGEMA_signal_3777) );
  DFF_X1 new_AGEMA_reg_buffer_1893_s_current_state_reg ( .D(
        new_AGEMA_signal_3780), .CK(clk), .Q(new_AGEMA_signal_3781) );
  DFF_X1 new_AGEMA_reg_buffer_1897_s_current_state_reg ( .D(
        new_AGEMA_signal_3784), .CK(clk), .Q(new_AGEMA_signal_3785) );
  DFF_X1 new_AGEMA_reg_buffer_1901_s_current_state_reg ( .D(
        new_AGEMA_signal_3788), .CK(clk), .Q(new_AGEMA_signal_3789) );
  DFF_X1 new_AGEMA_reg_buffer_1905_s_current_state_reg ( .D(
        new_AGEMA_signal_3792), .CK(clk), .Q(new_AGEMA_signal_3793) );
  DFF_X1 new_AGEMA_reg_buffer_1909_s_current_state_reg ( .D(
        new_AGEMA_signal_3796), .CK(clk), .Q(new_AGEMA_signal_3797) );
  DFF_X1 new_AGEMA_reg_buffer_1913_s_current_state_reg ( .D(
        new_AGEMA_signal_3800), .CK(clk), .Q(new_AGEMA_signal_3801) );
  DFF_X1 new_AGEMA_reg_buffer_1917_s_current_state_reg ( .D(
        new_AGEMA_signal_3804), .CK(clk), .Q(new_AGEMA_signal_3805) );
  DFF_X1 new_AGEMA_reg_buffer_1921_s_current_state_reg ( .D(
        new_AGEMA_signal_3808), .CK(clk), .Q(new_AGEMA_signal_3809) );
  DFF_X1 new_AGEMA_reg_buffer_1925_s_current_state_reg ( .D(
        new_AGEMA_signal_3812), .CK(clk), .Q(new_AGEMA_signal_3813) );
  DFF_X1 new_AGEMA_reg_buffer_1929_s_current_state_reg ( .D(
        new_AGEMA_signal_3816), .CK(clk), .Q(new_AGEMA_signal_3817) );
  DFF_X1 new_AGEMA_reg_buffer_1933_s_current_state_reg ( .D(
        new_AGEMA_signal_3820), .CK(clk), .Q(new_AGEMA_signal_3821) );
  DFF_X1 new_AGEMA_reg_buffer_1937_s_current_state_reg ( .D(
        new_AGEMA_signal_3824), .CK(clk), .Q(new_AGEMA_signal_3825) );
  DFF_X1 new_AGEMA_reg_buffer_1941_s_current_state_reg ( .D(
        new_AGEMA_signal_3828), .CK(clk), .Q(new_AGEMA_signal_3829) );
  DFF_X1 new_AGEMA_reg_buffer_1945_s_current_state_reg ( .D(
        new_AGEMA_signal_3832), .CK(clk), .Q(new_AGEMA_signal_3833) );
  DFF_X1 new_AGEMA_reg_buffer_1949_s_current_state_reg ( .D(
        new_AGEMA_signal_3836), .CK(clk), .Q(new_AGEMA_signal_3837) );
  DFF_X1 new_AGEMA_reg_buffer_1953_s_current_state_reg ( .D(
        new_AGEMA_signal_3840), .CK(clk), .Q(new_AGEMA_signal_3841) );
  DFF_X1 new_AGEMA_reg_buffer_1957_s_current_state_reg ( .D(
        new_AGEMA_signal_3844), .CK(clk), .Q(new_AGEMA_signal_3845) );
  DFF_X1 new_AGEMA_reg_buffer_1961_s_current_state_reg ( .D(
        new_AGEMA_signal_3848), .CK(clk), .Q(new_AGEMA_signal_3849) );
  DFF_X1 new_AGEMA_reg_buffer_1965_s_current_state_reg ( .D(
        new_AGEMA_signal_3852), .CK(clk), .Q(new_AGEMA_signal_3853) );
  DFF_X1 new_AGEMA_reg_buffer_1969_s_current_state_reg ( .D(
        new_AGEMA_signal_3856), .CK(clk), .Q(new_AGEMA_signal_3857) );
  DFF_X1 new_AGEMA_reg_buffer_1973_s_current_state_reg ( .D(
        new_AGEMA_signal_3860), .CK(clk), .Q(new_AGEMA_signal_3861) );
  DFF_X1 new_AGEMA_reg_buffer_1977_s_current_state_reg ( .D(
        new_AGEMA_signal_3864), .CK(clk), .Q(new_AGEMA_signal_3865) );
  DFF_X1 new_AGEMA_reg_buffer_1981_s_current_state_reg ( .D(
        new_AGEMA_signal_3868), .CK(clk), .Q(new_AGEMA_signal_3869) );
  DFF_X1 new_AGEMA_reg_buffer_1985_s_current_state_reg ( .D(
        new_AGEMA_signal_3872), .CK(clk), .Q(new_AGEMA_signal_3873) );
  DFF_X1 new_AGEMA_reg_buffer_1989_s_current_state_reg ( .D(
        new_AGEMA_signal_3876), .CK(clk), .Q(new_AGEMA_signal_3877) );
  DFF_X1 new_AGEMA_reg_buffer_1993_s_current_state_reg ( .D(
        new_AGEMA_signal_3880), .CK(clk), .Q(new_AGEMA_signal_3881) );
  DFF_X1 new_AGEMA_reg_buffer_1997_s_current_state_reg ( .D(
        new_AGEMA_signal_3884), .CK(clk), .Q(new_AGEMA_signal_3885) );
  DFF_X1 new_AGEMA_reg_buffer_2001_s_current_state_reg ( .D(
        new_AGEMA_signal_3888), .CK(clk), .Q(new_AGEMA_signal_3889) );
  DFF_X1 new_AGEMA_reg_buffer_2005_s_current_state_reg ( .D(
        new_AGEMA_signal_3892), .CK(clk), .Q(new_AGEMA_signal_3893) );
  DFF_X1 new_AGEMA_reg_buffer_2009_s_current_state_reg ( .D(
        new_AGEMA_signal_3896), .CK(clk), .Q(new_AGEMA_signal_3897) );
  DFF_X1 new_AGEMA_reg_buffer_2013_s_current_state_reg ( .D(
        new_AGEMA_signal_3900), .CK(clk), .Q(new_AGEMA_signal_3901) );
  DFF_X1 new_AGEMA_reg_buffer_2017_s_current_state_reg ( .D(
        new_AGEMA_signal_3904), .CK(clk), .Q(new_AGEMA_signal_3905) );
  DFF_X1 new_AGEMA_reg_buffer_2021_s_current_state_reg ( .D(
        new_AGEMA_signal_3908), .CK(clk), .Q(new_AGEMA_signal_3909) );
  DFF_X1 new_AGEMA_reg_buffer_2025_s_current_state_reg ( .D(
        new_AGEMA_signal_3912), .CK(clk), .Q(new_AGEMA_signal_3913) );
  DFF_X1 new_AGEMA_reg_buffer_2029_s_current_state_reg ( .D(
        new_AGEMA_signal_3916), .CK(clk), .Q(new_AGEMA_signal_3917) );
  DFF_X1 new_AGEMA_reg_buffer_2033_s_current_state_reg ( .D(
        new_AGEMA_signal_3920), .CK(clk), .Q(new_AGEMA_signal_3921) );
  DFF_X1 new_AGEMA_reg_buffer_2037_s_current_state_reg ( .D(
        new_AGEMA_signal_3924), .CK(clk), .Q(new_AGEMA_signal_3925) );
  DFF_X1 new_AGEMA_reg_buffer_2041_s_current_state_reg ( .D(
        new_AGEMA_signal_3928), .CK(clk), .Q(new_AGEMA_signal_3929) );
  DFF_X1 new_AGEMA_reg_buffer_2045_s_current_state_reg ( .D(
        new_AGEMA_signal_3932), .CK(clk), .Q(new_AGEMA_signal_3933) );
  DFF_X1 new_AGEMA_reg_buffer_2049_s_current_state_reg ( .D(
        new_AGEMA_signal_3936), .CK(clk), .Q(new_AGEMA_signal_3937) );
  DFF_X1 new_AGEMA_reg_buffer_2053_s_current_state_reg ( .D(
        new_AGEMA_signal_3940), .CK(clk), .Q(new_AGEMA_signal_3941) );
  DFF_X1 new_AGEMA_reg_buffer_2057_s_current_state_reg ( .D(
        new_AGEMA_signal_3944), .CK(clk), .Q(new_AGEMA_signal_3945) );
  DFF_X1 new_AGEMA_reg_buffer_2061_s_current_state_reg ( .D(
        new_AGEMA_signal_3948), .CK(clk), .Q(new_AGEMA_signal_3949) );
  DFF_X1 new_AGEMA_reg_buffer_2065_s_current_state_reg ( .D(
        new_AGEMA_signal_3952), .CK(clk), .Q(new_AGEMA_signal_3953) );
  DFF_X1 new_AGEMA_reg_buffer_2069_s_current_state_reg ( .D(
        new_AGEMA_signal_3956), .CK(clk), .Q(new_AGEMA_signal_3957) );
  DFF_X1 new_AGEMA_reg_buffer_2073_s_current_state_reg ( .D(
        new_AGEMA_signal_3960), .CK(clk), .Q(new_AGEMA_signal_3961) );
  DFF_X1 new_AGEMA_reg_buffer_2077_s_current_state_reg ( .D(
        new_AGEMA_signal_3964), .CK(clk), .Q(new_AGEMA_signal_3965) );
  DFF_X1 new_AGEMA_reg_buffer_2081_s_current_state_reg ( .D(
        new_AGEMA_signal_3968), .CK(clk), .Q(new_AGEMA_signal_3969) );
  DFF_X1 new_AGEMA_reg_buffer_2085_s_current_state_reg ( .D(
        new_AGEMA_signal_3972), .CK(clk), .Q(new_AGEMA_signal_3973) );
  DFF_X1 new_AGEMA_reg_buffer_2089_s_current_state_reg ( .D(
        new_AGEMA_signal_3976), .CK(clk), .Q(new_AGEMA_signal_3977) );
  DFF_X1 new_AGEMA_reg_buffer_2093_s_current_state_reg ( .D(
        new_AGEMA_signal_3980), .CK(clk), .Q(new_AGEMA_signal_3981) );
  DFF_X1 new_AGEMA_reg_buffer_2097_s_current_state_reg ( .D(
        new_AGEMA_signal_3984), .CK(clk), .Q(new_AGEMA_signal_3985) );
  DFF_X1 new_AGEMA_reg_buffer_2101_s_current_state_reg ( .D(
        new_AGEMA_signal_3988), .CK(clk), .Q(new_AGEMA_signal_3989) );
  DFF_X1 new_AGEMA_reg_buffer_2105_s_current_state_reg ( .D(
        new_AGEMA_signal_3992), .CK(clk), .Q(new_AGEMA_signal_3993) );
  DFF_X1 new_AGEMA_reg_buffer_2109_s_current_state_reg ( .D(
        new_AGEMA_signal_3996), .CK(clk), .Q(new_AGEMA_signal_3997) );
  DFF_X1 new_AGEMA_reg_buffer_2113_s_current_state_reg ( .D(
        new_AGEMA_signal_4000), .CK(clk), .Q(new_AGEMA_signal_4001) );
  DFF_X1 new_AGEMA_reg_buffer_2117_s_current_state_reg ( .D(
        new_AGEMA_signal_4004), .CK(clk), .Q(new_AGEMA_signal_4005) );
  DFF_X1 new_AGEMA_reg_buffer_2121_s_current_state_reg ( .D(
        new_AGEMA_signal_4008), .CK(clk), .Q(new_AGEMA_signal_4009) );
  DFF_X1 new_AGEMA_reg_buffer_2125_s_current_state_reg ( .D(
        new_AGEMA_signal_4012), .CK(clk), .Q(new_AGEMA_signal_4013) );
  DFF_X1 new_AGEMA_reg_buffer_2129_s_current_state_reg ( .D(
        new_AGEMA_signal_4016), .CK(clk), .Q(new_AGEMA_signal_4017) );
  DFF_X1 new_AGEMA_reg_buffer_2133_s_current_state_reg ( .D(
        new_AGEMA_signal_4020), .CK(clk), .Q(new_AGEMA_signal_4021) );
  DFF_X1 new_AGEMA_reg_buffer_2137_s_current_state_reg ( .D(
        new_AGEMA_signal_4024), .CK(clk), .Q(new_AGEMA_signal_4025) );
  DFF_X1 new_AGEMA_reg_buffer_2141_s_current_state_reg ( .D(
        new_AGEMA_signal_4028), .CK(clk), .Q(new_AGEMA_signal_4029) );
  DFF_X1 new_AGEMA_reg_buffer_2145_s_current_state_reg ( .D(
        new_AGEMA_signal_4032), .CK(clk), .Q(new_AGEMA_signal_4033) );
  DFF_X1 new_AGEMA_reg_buffer_2149_s_current_state_reg ( .D(
        new_AGEMA_signal_4036), .CK(clk), .Q(new_AGEMA_signal_4037) );
  DFF_X1 new_AGEMA_reg_buffer_2153_s_current_state_reg ( .D(
        new_AGEMA_signal_4040), .CK(clk), .Q(new_AGEMA_signal_4041) );
  DFF_X1 new_AGEMA_reg_buffer_2157_s_current_state_reg ( .D(
        new_AGEMA_signal_4044), .CK(clk), .Q(new_AGEMA_signal_4045) );
  DFF_X1 new_AGEMA_reg_buffer_2161_s_current_state_reg ( .D(
        new_AGEMA_signal_4048), .CK(clk), .Q(new_AGEMA_signal_4049) );
  DFF_X1 new_AGEMA_reg_buffer_2165_s_current_state_reg ( .D(
        new_AGEMA_signal_4052), .CK(clk), .Q(new_AGEMA_signal_4053) );
  DFF_X1 new_AGEMA_reg_buffer_2169_s_current_state_reg ( .D(
        new_AGEMA_signal_4056), .CK(clk), .Q(new_AGEMA_signal_4057) );
  DFF_X1 new_AGEMA_reg_buffer_2173_s_current_state_reg ( .D(
        new_AGEMA_signal_4060), .CK(clk), .Q(new_AGEMA_signal_4061) );
  DFF_X1 new_AGEMA_reg_buffer_2177_s_current_state_reg ( .D(
        new_AGEMA_signal_4064), .CK(clk), .Q(new_AGEMA_signal_4065) );
  DFF_X1 new_AGEMA_reg_buffer_2181_s_current_state_reg ( .D(
        new_AGEMA_signal_4068), .CK(clk), .Q(new_AGEMA_signal_4069) );
  DFF_X1 new_AGEMA_reg_buffer_2185_s_current_state_reg ( .D(
        new_AGEMA_signal_4072), .CK(clk), .Q(new_AGEMA_signal_4073) );
  DFF_X1 new_AGEMA_reg_buffer_2189_s_current_state_reg ( .D(
        new_AGEMA_signal_4076), .CK(clk), .Q(new_AGEMA_signal_4077) );
  DFF_X1 new_AGEMA_reg_buffer_2193_s_current_state_reg ( .D(
        new_AGEMA_signal_4080), .CK(clk), .Q(new_AGEMA_signal_4081) );
  DFF_X1 new_AGEMA_reg_buffer_2197_s_current_state_reg ( .D(
        new_AGEMA_signal_4084), .CK(clk), .Q(new_AGEMA_signal_4085) );
  DFF_X1 new_AGEMA_reg_buffer_2201_s_current_state_reg ( .D(
        new_AGEMA_signal_4088), .CK(clk), .Q(new_AGEMA_signal_4089) );
  DFF_X1 new_AGEMA_reg_buffer_2205_s_current_state_reg ( .D(
        new_AGEMA_signal_4092), .CK(clk), .Q(new_AGEMA_signal_4093) );
  DFF_X1 new_AGEMA_reg_buffer_2209_s_current_state_reg ( .D(
        new_AGEMA_signal_4096), .CK(clk), .Q(new_AGEMA_signal_4097) );
  DFF_X1 new_AGEMA_reg_buffer_2213_s_current_state_reg ( .D(
        new_AGEMA_signal_4100), .CK(clk), .Q(new_AGEMA_signal_4101) );
  DFF_X1 new_AGEMA_reg_buffer_2217_s_current_state_reg ( .D(
        new_AGEMA_signal_4104), .CK(clk), .Q(new_AGEMA_signal_4105) );
  DFF_X1 new_AGEMA_reg_buffer_2221_s_current_state_reg ( .D(
        new_AGEMA_signal_4108), .CK(clk), .Q(new_AGEMA_signal_4109) );
  DFF_X1 new_AGEMA_reg_buffer_2225_s_current_state_reg ( .D(
        new_AGEMA_signal_4112), .CK(clk), .Q(new_AGEMA_signal_4113) );
  DFF_X1 new_AGEMA_reg_buffer_2229_s_current_state_reg ( .D(
        new_AGEMA_signal_4116), .CK(clk), .Q(new_AGEMA_signal_4117) );
  DFF_X1 new_AGEMA_reg_buffer_2233_s_current_state_reg ( .D(
        new_AGEMA_signal_4120), .CK(clk), .Q(new_AGEMA_signal_4121) );
  DFF_X1 new_AGEMA_reg_buffer_2237_s_current_state_reg ( .D(
        new_AGEMA_signal_4124), .CK(clk), .Q(new_AGEMA_signal_4125) );
  DFF_X1 new_AGEMA_reg_buffer_2241_s_current_state_reg ( .D(
        new_AGEMA_signal_4128), .CK(clk), .Q(new_AGEMA_signal_4129) );
  DFF_X1 new_AGEMA_reg_buffer_2353_s_current_state_reg ( .D(
        new_AGEMA_signal_4240), .CK(clk), .Q(new_AGEMA_signal_4241) );
  DFF_X1 new_AGEMA_reg_buffer_2357_s_current_state_reg ( .D(
        new_AGEMA_signal_4244), .CK(clk), .Q(new_AGEMA_signal_4245) );
  DFF_X1 new_AGEMA_reg_buffer_2361_s_current_state_reg ( .D(
        new_AGEMA_signal_4248), .CK(clk), .Q(new_AGEMA_signal_4249) );
  DFF_X1 new_AGEMA_reg_buffer_2365_s_current_state_reg ( .D(
        new_AGEMA_signal_4252), .CK(clk), .Q(new_AGEMA_signal_4253) );
  DFF_X1 new_AGEMA_reg_buffer_2369_s_current_state_reg ( .D(
        new_AGEMA_signal_4256), .CK(clk), .Q(new_AGEMA_signal_4257) );
  DFF_X1 new_AGEMA_reg_buffer_2373_s_current_state_reg ( .D(
        new_AGEMA_signal_4260), .CK(clk), .Q(new_AGEMA_signal_4261) );
  DFF_X1 new_AGEMA_reg_buffer_2377_s_current_state_reg ( .D(
        new_AGEMA_signal_4264), .CK(clk), .Q(new_AGEMA_signal_4265) );
  DFF_X1 new_AGEMA_reg_buffer_2381_s_current_state_reg ( .D(
        new_AGEMA_signal_4268), .CK(clk), .Q(new_AGEMA_signal_4269) );
  DFF_X1 new_AGEMA_reg_buffer_2385_s_current_state_reg ( .D(
        new_AGEMA_signal_4272), .CK(clk), .Q(new_AGEMA_signal_4273) );
  DFF_X1 new_AGEMA_reg_buffer_2389_s_current_state_reg ( .D(
        new_AGEMA_signal_4276), .CK(clk), .Q(new_AGEMA_signal_4277) );
  DFF_X1 new_AGEMA_reg_buffer_2393_s_current_state_reg ( .D(
        new_AGEMA_signal_4280), .CK(clk), .Q(new_AGEMA_signal_4281) );
  DFF_X1 new_AGEMA_reg_buffer_2397_s_current_state_reg ( .D(
        new_AGEMA_signal_4284), .CK(clk), .Q(new_AGEMA_signal_4285) );
  DFF_X1 new_AGEMA_reg_buffer_2401_s_current_state_reg ( .D(
        new_AGEMA_signal_4288), .CK(clk), .Q(new_AGEMA_signal_4289) );
  DFF_X1 new_AGEMA_reg_buffer_2405_s_current_state_reg ( .D(
        new_AGEMA_signal_4292), .CK(clk), .Q(new_AGEMA_signal_4293) );
  DFF_X1 new_AGEMA_reg_buffer_2409_s_current_state_reg ( .D(
        new_AGEMA_signal_4296), .CK(clk), .Q(new_AGEMA_signal_4297) );
  DFF_X1 new_AGEMA_reg_buffer_2413_s_current_state_reg ( .D(
        new_AGEMA_signal_4300), .CK(clk), .Q(new_AGEMA_signal_4301) );
  DFF_X1 new_AGEMA_reg_buffer_2417_s_current_state_reg ( .D(
        new_AGEMA_signal_4304), .CK(clk), .Q(new_AGEMA_signal_4305) );
  DFF_X1 new_AGEMA_reg_buffer_2421_s_current_state_reg ( .D(
        new_AGEMA_signal_4308), .CK(clk), .Q(new_AGEMA_signal_4309) );
  DFF_X1 new_AGEMA_reg_buffer_2425_s_current_state_reg ( .D(
        new_AGEMA_signal_4312), .CK(clk), .Q(new_AGEMA_signal_4313) );
  DFF_X1 new_AGEMA_reg_buffer_2429_s_current_state_reg ( .D(
        new_AGEMA_signal_4316), .CK(clk), .Q(new_AGEMA_signal_4317) );
  DFF_X1 new_AGEMA_reg_buffer_2433_s_current_state_reg ( .D(
        new_AGEMA_signal_4320), .CK(clk), .Q(new_AGEMA_signal_4321) );
  DFF_X1 new_AGEMA_reg_buffer_2437_s_current_state_reg ( .D(
        new_AGEMA_signal_4324), .CK(clk), .Q(new_AGEMA_signal_4325) );
  DFF_X1 new_AGEMA_reg_buffer_2441_s_current_state_reg ( .D(
        new_AGEMA_signal_4328), .CK(clk), .Q(new_AGEMA_signal_4329) );
  DFF_X1 new_AGEMA_reg_buffer_2445_s_current_state_reg ( .D(
        new_AGEMA_signal_4332), .CK(clk), .Q(new_AGEMA_signal_4333) );
  DFF_X1 new_AGEMA_reg_buffer_2449_s_current_state_reg ( .D(
        new_AGEMA_signal_4336), .CK(clk), .Q(new_AGEMA_signal_4337) );
  DFF_X1 new_AGEMA_reg_buffer_2453_s_current_state_reg ( .D(
        new_AGEMA_signal_4340), .CK(clk), .Q(new_AGEMA_signal_4341) );
  DFF_X1 new_AGEMA_reg_buffer_2457_s_current_state_reg ( .D(
        new_AGEMA_signal_4344), .CK(clk), .Q(new_AGEMA_signal_4345) );
  DFF_X1 new_AGEMA_reg_buffer_2461_s_current_state_reg ( .D(
        new_AGEMA_signal_4348), .CK(clk), .Q(new_AGEMA_signal_4349) );
  DFF_X1 new_AGEMA_reg_buffer_2465_s_current_state_reg ( .D(
        new_AGEMA_signal_4352), .CK(clk), .Q(new_AGEMA_signal_4353) );
  DFF_X1 new_AGEMA_reg_buffer_2469_s_current_state_reg ( .D(
        new_AGEMA_signal_4356), .CK(clk), .Q(new_AGEMA_signal_4357) );
  DFF_X1 new_AGEMA_reg_buffer_2473_s_current_state_reg ( .D(
        new_AGEMA_signal_4360), .CK(clk), .Q(new_AGEMA_signal_4361) );
  DFF_X1 new_AGEMA_reg_buffer_2477_s_current_state_reg ( .D(
        new_AGEMA_signal_4364), .CK(clk), .Q(new_AGEMA_signal_4365) );
  DFF_X1 new_AGEMA_reg_buffer_2481_s_current_state_reg ( .D(
        new_AGEMA_signal_4368), .CK(clk), .Q(new_AGEMA_signal_4369) );
  DFF_X1 new_AGEMA_reg_buffer_2485_s_current_state_reg ( .D(
        new_AGEMA_signal_4372), .CK(clk), .Q(new_AGEMA_signal_4373) );
  DFF_X1 new_AGEMA_reg_buffer_2489_s_current_state_reg ( .D(
        new_AGEMA_signal_4376), .CK(clk), .Q(new_AGEMA_signal_4377) );
  DFF_X1 new_AGEMA_reg_buffer_2493_s_current_state_reg ( .D(
        new_AGEMA_signal_4380), .CK(clk), .Q(new_AGEMA_signal_4381) );
  DFF_X1 new_AGEMA_reg_buffer_2497_s_current_state_reg ( .D(
        new_AGEMA_signal_4384), .CK(clk), .Q(new_AGEMA_signal_4385) );
  DFF_X1 new_AGEMA_reg_buffer_2501_s_current_state_reg ( .D(
        new_AGEMA_signal_4388), .CK(clk), .Q(new_AGEMA_signal_4389) );
  DFF_X1 new_AGEMA_reg_buffer_2505_s_current_state_reg ( .D(
        new_AGEMA_signal_4392), .CK(clk), .Q(new_AGEMA_signal_4393) );
  DFF_X1 new_AGEMA_reg_buffer_2509_s_current_state_reg ( .D(
        new_AGEMA_signal_4396), .CK(clk), .Q(new_AGEMA_signal_4397) );
  DFF_X1 new_AGEMA_reg_buffer_2513_s_current_state_reg ( .D(
        new_AGEMA_signal_4400), .CK(clk), .Q(new_AGEMA_signal_4401) );
  DFF_X1 new_AGEMA_reg_buffer_2517_s_current_state_reg ( .D(
        new_AGEMA_signal_4404), .CK(clk), .Q(new_AGEMA_signal_4405) );
  DFF_X1 new_AGEMA_reg_buffer_2521_s_current_state_reg ( .D(
        new_AGEMA_signal_4408), .CK(clk), .Q(new_AGEMA_signal_4409) );
  DFF_X1 new_AGEMA_reg_buffer_2525_s_current_state_reg ( .D(
        new_AGEMA_signal_4412), .CK(clk), .Q(new_AGEMA_signal_4413) );
  DFF_X1 new_AGEMA_reg_buffer_2529_s_current_state_reg ( .D(
        new_AGEMA_signal_4416), .CK(clk), .Q(new_AGEMA_signal_4417) );
  DFF_X1 new_AGEMA_reg_buffer_2533_s_current_state_reg ( .D(
        new_AGEMA_signal_4420), .CK(clk), .Q(new_AGEMA_signal_4421) );
  DFF_X1 new_AGEMA_reg_buffer_2537_s_current_state_reg ( .D(
        new_AGEMA_signal_4424), .CK(clk), .Q(new_AGEMA_signal_4425) );
  DFF_X1 new_AGEMA_reg_buffer_2541_s_current_state_reg ( .D(
        new_AGEMA_signal_4428), .CK(clk), .Q(new_AGEMA_signal_4429) );
  DFF_X1 new_AGEMA_reg_buffer_2545_s_current_state_reg ( .D(
        new_AGEMA_signal_4432), .CK(clk), .Q(new_AGEMA_signal_4433) );
  DFF_X1 new_AGEMA_reg_buffer_2549_s_current_state_reg ( .D(
        new_AGEMA_signal_4436), .CK(clk), .Q(new_AGEMA_signal_4437) );
  DFF_X1 new_AGEMA_reg_buffer_2553_s_current_state_reg ( .D(
        new_AGEMA_signal_4440), .CK(clk), .Q(new_AGEMA_signal_4441) );
  DFF_X1 new_AGEMA_reg_buffer_2557_s_current_state_reg ( .D(
        new_AGEMA_signal_4444), .CK(clk), .Q(new_AGEMA_signal_4445) );
  DFF_X1 new_AGEMA_reg_buffer_2561_s_current_state_reg ( .D(
        new_AGEMA_signal_4448), .CK(clk), .Q(new_AGEMA_signal_4449) );
  DFF_X1 new_AGEMA_reg_buffer_2565_s_current_state_reg ( .D(
        new_AGEMA_signal_4452), .CK(clk), .Q(new_AGEMA_signal_4453) );
  DFF_X1 new_AGEMA_reg_buffer_2569_s_current_state_reg ( .D(
        new_AGEMA_signal_4456), .CK(clk), .Q(new_AGEMA_signal_4457) );
  DFF_X1 new_AGEMA_reg_buffer_2573_s_current_state_reg ( .D(
        new_AGEMA_signal_4460), .CK(clk), .Q(new_AGEMA_signal_4461) );
  DFF_X1 new_AGEMA_reg_buffer_2577_s_current_state_reg ( .D(
        new_AGEMA_signal_4464), .CK(clk), .Q(new_AGEMA_signal_4465) );
  DFF_X1 new_AGEMA_reg_buffer_2581_s_current_state_reg ( .D(
        new_AGEMA_signal_4468), .CK(clk), .Q(new_AGEMA_signal_4469) );
  DFF_X1 new_AGEMA_reg_buffer_2585_s_current_state_reg ( .D(
        new_AGEMA_signal_4472), .CK(clk), .Q(new_AGEMA_signal_4473) );
  DFF_X1 new_AGEMA_reg_buffer_2589_s_current_state_reg ( .D(
        new_AGEMA_signal_4476), .CK(clk), .Q(new_AGEMA_signal_4477) );
  DFF_X1 new_AGEMA_reg_buffer_2593_s_current_state_reg ( .D(
        new_AGEMA_signal_4480), .CK(clk), .Q(new_AGEMA_signal_4481) );
  DFF_X1 new_AGEMA_reg_buffer_2597_s_current_state_reg ( .D(
        new_AGEMA_signal_4484), .CK(clk), .Q(new_AGEMA_signal_4485) );
  DFF_X1 new_AGEMA_reg_buffer_2601_s_current_state_reg ( .D(
        new_AGEMA_signal_4488), .CK(clk), .Q(new_AGEMA_signal_4489) );
  DFF_X1 new_AGEMA_reg_buffer_2605_s_current_state_reg ( .D(
        new_AGEMA_signal_4492), .CK(clk), .Q(new_AGEMA_signal_4493) );
  DFF_X1 new_AGEMA_reg_buffer_2609_s_current_state_reg ( .D(
        new_AGEMA_signal_4496), .CK(clk), .Q(new_AGEMA_signal_4497) );
  DFF_X1 new_AGEMA_reg_buffer_2613_s_current_state_reg ( .D(
        new_AGEMA_signal_4500), .CK(clk), .Q(new_AGEMA_signal_4501) );
  DFF_X1 new_AGEMA_reg_buffer_2617_s_current_state_reg ( .D(
        new_AGEMA_signal_4504), .CK(clk), .Q(new_AGEMA_signal_4505) );
  DFF_X1 new_AGEMA_reg_buffer_2621_s_current_state_reg ( .D(
        new_AGEMA_signal_4508), .CK(clk), .Q(new_AGEMA_signal_4509) );
  DFF_X1 new_AGEMA_reg_buffer_2625_s_current_state_reg ( .D(
        new_AGEMA_signal_4512), .CK(clk), .Q(new_AGEMA_signal_4513) );
  DFF_X1 new_AGEMA_reg_buffer_2629_s_current_state_reg ( .D(
        new_AGEMA_signal_4516), .CK(clk), .Q(new_AGEMA_signal_4517) );
  DFF_X1 new_AGEMA_reg_buffer_2633_s_current_state_reg ( .D(
        new_AGEMA_signal_4520), .CK(clk), .Q(new_AGEMA_signal_4521) );
  DFF_X1 new_AGEMA_reg_buffer_2637_s_current_state_reg ( .D(
        new_AGEMA_signal_4524), .CK(clk), .Q(new_AGEMA_signal_4525) );
  DFF_X1 new_AGEMA_reg_buffer_2641_s_current_state_reg ( .D(
        new_AGEMA_signal_4528), .CK(clk), .Q(new_AGEMA_signal_4529) );
  DFF_X1 new_AGEMA_reg_buffer_2645_s_current_state_reg ( .D(
        new_AGEMA_signal_4532), .CK(clk), .Q(new_AGEMA_signal_4533) );
  DFF_X1 new_AGEMA_reg_buffer_2649_s_current_state_reg ( .D(
        new_AGEMA_signal_4536), .CK(clk), .Q(new_AGEMA_signal_4537) );
  DFF_X1 new_AGEMA_reg_buffer_2653_s_current_state_reg ( .D(
        new_AGEMA_signal_4540), .CK(clk), .Q(new_AGEMA_signal_4541) );
  DFF_X1 new_AGEMA_reg_buffer_2657_s_current_state_reg ( .D(
        new_AGEMA_signal_4544), .CK(clk), .Q(new_AGEMA_signal_4545) );
  DFF_X1 new_AGEMA_reg_buffer_2661_s_current_state_reg ( .D(
        new_AGEMA_signal_4548), .CK(clk), .Q(new_AGEMA_signal_4549) );
  DFF_X1 new_AGEMA_reg_buffer_2665_s_current_state_reg ( .D(
        new_AGEMA_signal_4552), .CK(clk), .Q(new_AGEMA_signal_4553) );
  DFF_X1 new_AGEMA_reg_buffer_2669_s_current_state_reg ( .D(
        new_AGEMA_signal_4556), .CK(clk), .Q(new_AGEMA_signal_4557) );
  DFF_X1 new_AGEMA_reg_buffer_2673_s_current_state_reg ( .D(
        new_AGEMA_signal_4560), .CK(clk), .Q(new_AGEMA_signal_4561) );
  DFF_X1 new_AGEMA_reg_buffer_2677_s_current_state_reg ( .D(
        new_AGEMA_signal_4564), .CK(clk), .Q(new_AGEMA_signal_4565) );
  DFF_X1 new_AGEMA_reg_buffer_2681_s_current_state_reg ( .D(
        new_AGEMA_signal_4568), .CK(clk), .Q(new_AGEMA_signal_4569) );
  DFF_X1 new_AGEMA_reg_buffer_2685_s_current_state_reg ( .D(
        new_AGEMA_signal_4572), .CK(clk), .Q(new_AGEMA_signal_4573) );
  DFF_X1 new_AGEMA_reg_buffer_2689_s_current_state_reg ( .D(
        new_AGEMA_signal_4576), .CK(clk), .Q(new_AGEMA_signal_4577) );
  DFF_X1 new_AGEMA_reg_buffer_2693_s_current_state_reg ( .D(
        new_AGEMA_signal_4580), .CK(clk), .Q(new_AGEMA_signal_4581) );
  DFF_X1 new_AGEMA_reg_buffer_2697_s_current_state_reg ( .D(
        new_AGEMA_signal_4584), .CK(clk), .Q(new_AGEMA_signal_4585) );
  DFF_X1 new_AGEMA_reg_buffer_2701_s_current_state_reg ( .D(
        new_AGEMA_signal_4588), .CK(clk), .Q(new_AGEMA_signal_4589) );
  DFF_X1 new_AGEMA_reg_buffer_2705_s_current_state_reg ( .D(
        new_AGEMA_signal_4592), .CK(clk), .Q(new_AGEMA_signal_4593) );
  DFF_X1 new_AGEMA_reg_buffer_2709_s_current_state_reg ( .D(
        new_AGEMA_signal_4596), .CK(clk), .Q(new_AGEMA_signal_4597) );
  DFF_X1 new_AGEMA_reg_buffer_2713_s_current_state_reg ( .D(
        new_AGEMA_signal_4600), .CK(clk), .Q(new_AGEMA_signal_4601) );
  DFF_X1 new_AGEMA_reg_buffer_2717_s_current_state_reg ( .D(
        new_AGEMA_signal_4604), .CK(clk), .Q(new_AGEMA_signal_4605) );
  DFF_X1 new_AGEMA_reg_buffer_2721_s_current_state_reg ( .D(
        new_AGEMA_signal_4608), .CK(clk), .Q(new_AGEMA_signal_4609) );
  DFF_X1 new_AGEMA_reg_buffer_2725_s_current_state_reg ( .D(
        new_AGEMA_signal_4612), .CK(clk), .Q(new_AGEMA_signal_4613) );
  DFF_X1 new_AGEMA_reg_buffer_2729_s_current_state_reg ( .D(
        new_AGEMA_signal_4616), .CK(clk), .Q(new_AGEMA_signal_4617) );
  DFF_X1 new_AGEMA_reg_buffer_2733_s_current_state_reg ( .D(
        new_AGEMA_signal_4620), .CK(clk), .Q(new_AGEMA_signal_4621) );
  DFF_X1 new_AGEMA_reg_buffer_2737_s_current_state_reg ( .D(
        new_AGEMA_signal_4624), .CK(clk), .Q(new_AGEMA_signal_4625) );
  DFF_X1 new_AGEMA_reg_buffer_2741_s_current_state_reg ( .D(
        new_AGEMA_signal_4628), .CK(clk), .Q(new_AGEMA_signal_4629) );
  DFF_X1 new_AGEMA_reg_buffer_2745_s_current_state_reg ( .D(
        new_AGEMA_signal_4632), .CK(clk), .Q(new_AGEMA_signal_4633) );
  DFF_X1 new_AGEMA_reg_buffer_2749_s_current_state_reg ( .D(
        new_AGEMA_signal_4636), .CK(clk), .Q(new_AGEMA_signal_4637) );
  DFF_X1 new_AGEMA_reg_buffer_2753_s_current_state_reg ( .D(
        new_AGEMA_signal_4640), .CK(clk), .Q(new_AGEMA_signal_4641) );
  DFF_X1 new_AGEMA_reg_buffer_2757_s_current_state_reg ( .D(
        new_AGEMA_signal_4644), .CK(clk), .Q(new_AGEMA_signal_4645) );
  DFF_X1 new_AGEMA_reg_buffer_2761_s_current_state_reg ( .D(
        new_AGEMA_signal_4648), .CK(clk), .Q(new_AGEMA_signal_4649) );
  DFF_X1 new_AGEMA_reg_buffer_2765_s_current_state_reg ( .D(
        new_AGEMA_signal_4652), .CK(clk), .Q(new_AGEMA_signal_4653) );
  DFF_X1 new_AGEMA_reg_buffer_2769_s_current_state_reg ( .D(
        new_AGEMA_signal_4656), .CK(clk), .Q(new_AGEMA_signal_4657) );
  DFF_X1 new_AGEMA_reg_buffer_2773_s_current_state_reg ( .D(
        new_AGEMA_signal_4660), .CK(clk), .Q(new_AGEMA_signal_4661) );
  DFF_X1 new_AGEMA_reg_buffer_2777_s_current_state_reg ( .D(
        new_AGEMA_signal_4664), .CK(clk), .Q(new_AGEMA_signal_4665) );
  DFF_X1 new_AGEMA_reg_buffer_2781_s_current_state_reg ( .D(
        new_AGEMA_signal_4668), .CK(clk), .Q(new_AGEMA_signal_4669) );
  DFF_X1 new_AGEMA_reg_buffer_2785_s_current_state_reg ( .D(
        new_AGEMA_signal_4672), .CK(clk), .Q(new_AGEMA_signal_4673) );
  DFF_X1 new_AGEMA_reg_buffer_2789_s_current_state_reg ( .D(
        new_AGEMA_signal_4676), .CK(clk), .Q(new_AGEMA_signal_4677) );
  DFF_X1 new_AGEMA_reg_buffer_2793_s_current_state_reg ( .D(
        new_AGEMA_signal_4680), .CK(clk), .Q(new_AGEMA_signal_4681) );
  DFF_X1 new_AGEMA_reg_buffer_2797_s_current_state_reg ( .D(
        new_AGEMA_signal_4684), .CK(clk), .Q(new_AGEMA_signal_4685) );
  DFF_X1 new_AGEMA_reg_buffer_2801_s_current_state_reg ( .D(
        new_AGEMA_signal_4688), .CK(clk), .Q(new_AGEMA_signal_4689) );
  DFF_X1 new_AGEMA_reg_buffer_2805_s_current_state_reg ( .D(
        new_AGEMA_signal_4692), .CK(clk), .Q(new_AGEMA_signal_4693) );
  DFF_X1 new_AGEMA_reg_buffer_2809_s_current_state_reg ( .D(
        new_AGEMA_signal_4696), .CK(clk), .Q(new_AGEMA_signal_4697) );
  DFF_X1 new_AGEMA_reg_buffer_2813_s_current_state_reg ( .D(
        new_AGEMA_signal_4700), .CK(clk), .Q(new_AGEMA_signal_4701) );
  DFF_X1 new_AGEMA_reg_buffer_2817_s_current_state_reg ( .D(
        new_AGEMA_signal_4704), .CK(clk), .Q(new_AGEMA_signal_4705) );
  DFF_X1 new_AGEMA_reg_buffer_2821_s_current_state_reg ( .D(
        new_AGEMA_signal_4708), .CK(clk), .Q(new_AGEMA_signal_4709) );
  DFF_X1 new_AGEMA_reg_buffer_2825_s_current_state_reg ( .D(
        new_AGEMA_signal_4712), .CK(clk), .Q(new_AGEMA_signal_4713) );
  DFF_X1 new_AGEMA_reg_buffer_2829_s_current_state_reg ( .D(
        new_AGEMA_signal_4716), .CK(clk), .Q(new_AGEMA_signal_4717) );
  DFF_X1 new_AGEMA_reg_buffer_2833_s_current_state_reg ( .D(
        new_AGEMA_signal_4720), .CK(clk), .Q(new_AGEMA_signal_4721) );
  DFF_X1 new_AGEMA_reg_buffer_2837_s_current_state_reg ( .D(
        new_AGEMA_signal_4724), .CK(clk), .Q(new_AGEMA_signal_4725) );
  DFF_X1 new_AGEMA_reg_buffer_2841_s_current_state_reg ( .D(
        new_AGEMA_signal_4728), .CK(clk), .Q(new_AGEMA_signal_4729) );
  DFF_X1 new_AGEMA_reg_buffer_2845_s_current_state_reg ( .D(
        new_AGEMA_signal_4732), .CK(clk), .Q(new_AGEMA_signal_4733) );
  DFF_X1 new_AGEMA_reg_buffer_2849_s_current_state_reg ( .D(
        new_AGEMA_signal_4736), .CK(clk), .Q(new_AGEMA_signal_4737) );
  DFF_X1 new_AGEMA_reg_buffer_2853_s_current_state_reg ( .D(
        new_AGEMA_signal_4740), .CK(clk), .Q(new_AGEMA_signal_4741) );
  DFF_X1 new_AGEMA_reg_buffer_2857_s_current_state_reg ( .D(
        new_AGEMA_signal_4744), .CK(clk), .Q(new_AGEMA_signal_4745) );
  DFF_X1 new_AGEMA_reg_buffer_2861_s_current_state_reg ( .D(
        new_AGEMA_signal_4748), .CK(clk), .Q(new_AGEMA_signal_4749) );
  DFF_X1 new_AGEMA_reg_buffer_2865_s_current_state_reg ( .D(
        new_AGEMA_signal_4752), .CK(clk), .Q(new_AGEMA_signal_4753) );
  DFF_X1 new_AGEMA_reg_buffer_2869_s_current_state_reg ( .D(
        new_AGEMA_signal_4756), .CK(clk), .Q(new_AGEMA_signal_4757) );
  DFF_X1 new_AGEMA_reg_buffer_2873_s_current_state_reg ( .D(
        new_AGEMA_signal_4760), .CK(clk), .Q(new_AGEMA_signal_4761) );
  DFF_X1 new_AGEMA_reg_buffer_2877_s_current_state_reg ( .D(
        new_AGEMA_signal_4764), .CK(clk), .Q(new_AGEMA_signal_4765) );
  DFF_X1 new_AGEMA_reg_buffer_2881_s_current_state_reg ( .D(
        new_AGEMA_signal_4768), .CK(clk), .Q(new_AGEMA_signal_4769) );
  DFF_X1 new_AGEMA_reg_buffer_2885_s_current_state_reg ( .D(
        new_AGEMA_signal_4772), .CK(clk), .Q(new_AGEMA_signal_4773) );
  DFF_X1 new_AGEMA_reg_buffer_2889_s_current_state_reg ( .D(
        new_AGEMA_signal_4776), .CK(clk), .Q(new_AGEMA_signal_4777) );
  DFF_X1 new_AGEMA_reg_buffer_2893_s_current_state_reg ( .D(
        new_AGEMA_signal_4780), .CK(clk), .Q(new_AGEMA_signal_4781) );
  DFF_X1 new_AGEMA_reg_buffer_2897_s_current_state_reg ( .D(
        new_AGEMA_signal_4784), .CK(clk), .Q(new_AGEMA_signal_4785) );
  DFF_X1 new_AGEMA_reg_buffer_2901_s_current_state_reg ( .D(
        new_AGEMA_signal_4788), .CK(clk), .Q(new_AGEMA_signal_4789) );
  DFF_X1 new_AGEMA_reg_buffer_2905_s_current_state_reg ( .D(
        new_AGEMA_signal_4792), .CK(clk), .Q(new_AGEMA_signal_4793) );
  DFF_X1 new_AGEMA_reg_buffer_2909_s_current_state_reg ( .D(
        new_AGEMA_signal_4796), .CK(clk), .Q(new_AGEMA_signal_4797) );
  DFF_X1 new_AGEMA_reg_buffer_2913_s_current_state_reg ( .D(
        new_AGEMA_signal_4800), .CK(clk), .Q(new_AGEMA_signal_4801) );
  DFF_X1 new_AGEMA_reg_buffer_2917_s_current_state_reg ( .D(
        new_AGEMA_signal_4804), .CK(clk), .Q(new_AGEMA_signal_4805) );
  DFF_X1 new_AGEMA_reg_buffer_2921_s_current_state_reg ( .D(
        new_AGEMA_signal_4808), .CK(clk), .Q(new_AGEMA_signal_4809) );
  DFF_X1 new_AGEMA_reg_buffer_2925_s_current_state_reg ( .D(
        new_AGEMA_signal_4812), .CK(clk), .Q(new_AGEMA_signal_4813) );
  DFF_X1 new_AGEMA_reg_buffer_2929_s_current_state_reg ( .D(
        new_AGEMA_signal_4816), .CK(clk), .Q(new_AGEMA_signal_4817) );
  DFF_X1 new_AGEMA_reg_buffer_2933_s_current_state_reg ( .D(
        new_AGEMA_signal_4820), .CK(clk), .Q(new_AGEMA_signal_4821) );
  DFF_X1 new_AGEMA_reg_buffer_2937_s_current_state_reg ( .D(
        new_AGEMA_signal_4824), .CK(clk), .Q(new_AGEMA_signal_4825) );
  DFF_X1 new_AGEMA_reg_buffer_2941_s_current_state_reg ( .D(
        new_AGEMA_signal_4828), .CK(clk), .Q(new_AGEMA_signal_4829) );
  DFF_X1 new_AGEMA_reg_buffer_2945_s_current_state_reg ( .D(
        new_AGEMA_signal_4832), .CK(clk), .Q(new_AGEMA_signal_4833) );
  DFF_X1 new_AGEMA_reg_buffer_2949_s_current_state_reg ( .D(
        new_AGEMA_signal_4836), .CK(clk), .Q(new_AGEMA_signal_4837) );
  DFF_X1 new_AGEMA_reg_buffer_2953_s_current_state_reg ( .D(
        new_AGEMA_signal_4840), .CK(clk), .Q(new_AGEMA_signal_4841) );
  DFF_X1 new_AGEMA_reg_buffer_2957_s_current_state_reg ( .D(
        new_AGEMA_signal_4844), .CK(clk), .Q(new_AGEMA_signal_4845) );
  DFF_X1 new_AGEMA_reg_buffer_2961_s_current_state_reg ( .D(
        new_AGEMA_signal_4848), .CK(clk), .Q(new_AGEMA_signal_4849) );
  DFF_X1 new_AGEMA_reg_buffer_2965_s_current_state_reg ( .D(
        new_AGEMA_signal_4852), .CK(clk), .Q(new_AGEMA_signal_4853) );
  DFF_X1 new_AGEMA_reg_buffer_2969_s_current_state_reg ( .D(
        new_AGEMA_signal_4856), .CK(clk), .Q(new_AGEMA_signal_4857) );
  DFF_X1 new_AGEMA_reg_buffer_2973_s_current_state_reg ( .D(
        new_AGEMA_signal_4860), .CK(clk), .Q(new_AGEMA_signal_4861) );
  DFF_X1 new_AGEMA_reg_buffer_2977_s_current_state_reg ( .D(
        new_AGEMA_signal_4864), .CK(clk), .Q(new_AGEMA_signal_4865) );
  DFF_X1 new_AGEMA_reg_buffer_2981_s_current_state_reg ( .D(
        new_AGEMA_signal_4868), .CK(clk), .Q(new_AGEMA_signal_4869) );
  DFF_X1 new_AGEMA_reg_buffer_2985_s_current_state_reg ( .D(
        new_AGEMA_signal_4872), .CK(clk), .Q(new_AGEMA_signal_4873) );
  DFF_X1 new_AGEMA_reg_buffer_2989_s_current_state_reg ( .D(
        new_AGEMA_signal_4876), .CK(clk), .Q(new_AGEMA_signal_4877) );
  DFF_X1 new_AGEMA_reg_buffer_2993_s_current_state_reg ( .D(
        new_AGEMA_signal_4880), .CK(clk), .Q(new_AGEMA_signal_4881) );
  DFF_X1 new_AGEMA_reg_buffer_2997_s_current_state_reg ( .D(
        new_AGEMA_signal_4884), .CK(clk), .Q(new_AGEMA_signal_4885) );
  DFF_X1 new_AGEMA_reg_buffer_3001_s_current_state_reg ( .D(
        new_AGEMA_signal_4888), .CK(clk), .Q(new_AGEMA_signal_4889) );
  DFF_X1 new_AGEMA_reg_buffer_3005_s_current_state_reg ( .D(
        new_AGEMA_signal_4892), .CK(clk), .Q(new_AGEMA_signal_4893) );
  DFF_X1 new_AGEMA_reg_buffer_3009_s_current_state_reg ( .D(
        new_AGEMA_signal_4896), .CK(clk), .Q(new_AGEMA_signal_4897) );
  DFF_X1 new_AGEMA_reg_buffer_3013_s_current_state_reg ( .D(
        new_AGEMA_signal_4900), .CK(clk), .Q(new_AGEMA_signal_4901) );
  DFF_X1 new_AGEMA_reg_buffer_3017_s_current_state_reg ( .D(
        new_AGEMA_signal_4904), .CK(clk), .Q(new_AGEMA_signal_4905) );
  DFF_X1 new_AGEMA_reg_buffer_3021_s_current_state_reg ( .D(
        new_AGEMA_signal_4908), .CK(clk), .Q(new_AGEMA_signal_4909) );
  DFF_X1 new_AGEMA_reg_buffer_3025_s_current_state_reg ( .D(
        new_AGEMA_signal_4912), .CK(clk), .Q(new_AGEMA_signal_4913) );
  DFF_X1 new_AGEMA_reg_buffer_3029_s_current_state_reg ( .D(
        new_AGEMA_signal_4916), .CK(clk), .Q(new_AGEMA_signal_4917) );
  DFF_X1 new_AGEMA_reg_buffer_3033_s_current_state_reg ( .D(
        new_AGEMA_signal_4920), .CK(clk), .Q(new_AGEMA_signal_4921) );
  DFF_X1 new_AGEMA_reg_buffer_3037_s_current_state_reg ( .D(
        new_AGEMA_signal_4924), .CK(clk), .Q(new_AGEMA_signal_4925) );
  DFF_X1 new_AGEMA_reg_buffer_3041_s_current_state_reg ( .D(
        new_AGEMA_signal_4928), .CK(clk), .Q(new_AGEMA_signal_4929) );
  DFF_X1 new_AGEMA_reg_buffer_3045_s_current_state_reg ( .D(
        new_AGEMA_signal_4932), .CK(clk), .Q(new_AGEMA_signal_4933) );
  DFF_X1 new_AGEMA_reg_buffer_3049_s_current_state_reg ( .D(
        new_AGEMA_signal_4936), .CK(clk), .Q(new_AGEMA_signal_4937) );
  DFF_X1 new_AGEMA_reg_buffer_3053_s_current_state_reg ( .D(
        new_AGEMA_signal_4940), .CK(clk), .Q(new_AGEMA_signal_4941) );
  DFF_X1 new_AGEMA_reg_buffer_3057_s_current_state_reg ( .D(
        new_AGEMA_signal_4944), .CK(clk), .Q(new_AGEMA_signal_4945) );
  DFF_X1 new_AGEMA_reg_buffer_3061_s_current_state_reg ( .D(
        new_AGEMA_signal_4948), .CK(clk), .Q(new_AGEMA_signal_4949) );
  DFF_X1 new_AGEMA_reg_buffer_3065_s_current_state_reg ( .D(
        new_AGEMA_signal_4952), .CK(clk), .Q(new_AGEMA_signal_4953) );
  DFF_X1 new_AGEMA_reg_buffer_3069_s_current_state_reg ( .D(
        new_AGEMA_signal_4956), .CK(clk), .Q(new_AGEMA_signal_4957) );
  DFF_X1 new_AGEMA_reg_buffer_3073_s_current_state_reg ( .D(
        new_AGEMA_signal_4960), .CK(clk), .Q(new_AGEMA_signal_4961) );
  DFF_X1 new_AGEMA_reg_buffer_3077_s_current_state_reg ( .D(
        new_AGEMA_signal_4964), .CK(clk), .Q(new_AGEMA_signal_4965) );
  DFF_X1 new_AGEMA_reg_buffer_3081_s_current_state_reg ( .D(
        new_AGEMA_signal_4968), .CK(clk), .Q(new_AGEMA_signal_4969) );
  DFF_X1 new_AGEMA_reg_buffer_3085_s_current_state_reg ( .D(
        new_AGEMA_signal_4972), .CK(clk), .Q(new_AGEMA_signal_4973) );
  DFF_X1 new_AGEMA_reg_buffer_3089_s_current_state_reg ( .D(
        new_AGEMA_signal_4976), .CK(clk), .Q(new_AGEMA_signal_4977) );
  DFF_X1 new_AGEMA_reg_buffer_3093_s_current_state_reg ( .D(
        new_AGEMA_signal_4980), .CK(clk), .Q(new_AGEMA_signal_4981) );
  DFF_X1 new_AGEMA_reg_buffer_3097_s_current_state_reg ( .D(
        new_AGEMA_signal_4984), .CK(clk), .Q(new_AGEMA_signal_4985) );
  DFF_X1 new_AGEMA_reg_buffer_3101_s_current_state_reg ( .D(
        new_AGEMA_signal_4988), .CK(clk), .Q(new_AGEMA_signal_4989) );
  DFF_X1 new_AGEMA_reg_buffer_3105_s_current_state_reg ( .D(
        new_AGEMA_signal_4992), .CK(clk), .Q(new_AGEMA_signal_4993) );
  DFF_X1 new_AGEMA_reg_buffer_3109_s_current_state_reg ( .D(
        new_AGEMA_signal_4996), .CK(clk), .Q(new_AGEMA_signal_4997) );
  DFF_X1 new_AGEMA_reg_buffer_3113_s_current_state_reg ( .D(
        new_AGEMA_signal_5000), .CK(clk), .Q(new_AGEMA_signal_5001) );
  DFF_X1 new_AGEMA_reg_buffer_3117_s_current_state_reg ( .D(
        new_AGEMA_signal_5004), .CK(clk), .Q(new_AGEMA_signal_5005) );
  DFF_X1 new_AGEMA_reg_buffer_3121_s_current_state_reg ( .D(
        new_AGEMA_signal_5008), .CK(clk), .Q(new_AGEMA_signal_5009) );
  DFF_X1 new_AGEMA_reg_buffer_3125_s_current_state_reg ( .D(
        new_AGEMA_signal_5012), .CK(clk), .Q(new_AGEMA_signal_5013) );
  DFF_X1 new_AGEMA_reg_buffer_3129_s_current_state_reg ( .D(
        new_AGEMA_signal_5016), .CK(clk), .Q(new_AGEMA_signal_5017) );
  DFF_X1 new_AGEMA_reg_buffer_3133_s_current_state_reg ( .D(
        new_AGEMA_signal_5020), .CK(clk), .Q(new_AGEMA_signal_5021) );
  DFF_X1 new_AGEMA_reg_buffer_3137_s_current_state_reg ( .D(
        new_AGEMA_signal_5024), .CK(clk), .Q(new_AGEMA_signal_5025) );
  DFF_X1 new_AGEMA_reg_buffer_3141_s_current_state_reg ( .D(
        new_AGEMA_signal_5028), .CK(clk), .Q(new_AGEMA_signal_5029) );
  DFF_X1 new_AGEMA_reg_buffer_3145_s_current_state_reg ( .D(
        new_AGEMA_signal_5032), .CK(clk), .Q(new_AGEMA_signal_5033) );
  DFF_X1 new_AGEMA_reg_buffer_3149_s_current_state_reg ( .D(
        new_AGEMA_signal_5036), .CK(clk), .Q(new_AGEMA_signal_5037) );
  DFF_X1 new_AGEMA_reg_buffer_3153_s_current_state_reg ( .D(
        new_AGEMA_signal_5040), .CK(clk), .Q(new_AGEMA_signal_5041) );
  DFF_X1 new_AGEMA_reg_buffer_3157_s_current_state_reg ( .D(
        new_AGEMA_signal_5044), .CK(clk), .Q(new_AGEMA_signal_5045) );
  DFF_X1 new_AGEMA_reg_buffer_3161_s_current_state_reg ( .D(
        new_AGEMA_signal_5048), .CK(clk), .Q(new_AGEMA_signal_5049) );
  DFF_X1 new_AGEMA_reg_buffer_3165_s_current_state_reg ( .D(
        new_AGEMA_signal_5052), .CK(clk), .Q(new_AGEMA_signal_5053) );
  DFF_X1 new_AGEMA_reg_buffer_3169_s_current_state_reg ( .D(
        new_AGEMA_signal_5056), .CK(clk), .Q(new_AGEMA_signal_5057) );
  DFF_X1 new_AGEMA_reg_buffer_3173_s_current_state_reg ( .D(
        new_AGEMA_signal_5060), .CK(clk), .Q(new_AGEMA_signal_5061) );
  DFF_X1 new_AGEMA_reg_buffer_3177_s_current_state_reg ( .D(
        new_AGEMA_signal_5064), .CK(clk), .Q(new_AGEMA_signal_5065) );
  DFF_X1 new_AGEMA_reg_buffer_3181_s_current_state_reg ( .D(
        new_AGEMA_signal_5068), .CK(clk), .Q(new_AGEMA_signal_5069) );
  DFF_X1 new_AGEMA_reg_buffer_3185_s_current_state_reg ( .D(
        new_AGEMA_signal_5072), .CK(clk), .Q(new_AGEMA_signal_5073) );
  DFF_X1 new_AGEMA_reg_buffer_3189_s_current_state_reg ( .D(
        new_AGEMA_signal_5076), .CK(clk), .Q(new_AGEMA_signal_5077) );
  DFF_X1 new_AGEMA_reg_buffer_3193_s_current_state_reg ( .D(
        new_AGEMA_signal_5080), .CK(clk), .Q(new_AGEMA_signal_5081) );
  DFF_X1 new_AGEMA_reg_buffer_3197_s_current_state_reg ( .D(
        new_AGEMA_signal_5084), .CK(clk), .Q(new_AGEMA_signal_5085) );
  DFF_X1 new_AGEMA_reg_buffer_3201_s_current_state_reg ( .D(
        new_AGEMA_signal_5088), .CK(clk), .Q(new_AGEMA_signal_5089) );
  DFF_X1 new_AGEMA_reg_buffer_3205_s_current_state_reg ( .D(
        new_AGEMA_signal_5092), .CK(clk), .Q(new_AGEMA_signal_5093) );
  DFF_X1 new_AGEMA_reg_buffer_3209_s_current_state_reg ( .D(
        new_AGEMA_signal_5096), .CK(clk), .Q(new_AGEMA_signal_5097) );
  DFF_X1 new_AGEMA_reg_buffer_3213_s_current_state_reg ( .D(
        new_AGEMA_signal_5100), .CK(clk), .Q(new_AGEMA_signal_5101) );
  DFF_X1 new_AGEMA_reg_buffer_3217_s_current_state_reg ( .D(
        new_AGEMA_signal_5104), .CK(clk), .Q(new_AGEMA_signal_5105) );
  DFF_X1 new_AGEMA_reg_buffer_3221_s_current_state_reg ( .D(
        new_AGEMA_signal_5108), .CK(clk), .Q(new_AGEMA_signal_5109) );
  DFF_X1 new_AGEMA_reg_buffer_3225_s_current_state_reg ( .D(
        new_AGEMA_signal_5112), .CK(clk), .Q(new_AGEMA_signal_5113) );
  DFF_X1 new_AGEMA_reg_buffer_3229_s_current_state_reg ( .D(
        new_AGEMA_signal_5116), .CK(clk), .Q(new_AGEMA_signal_5117) );
  DFF_X1 new_AGEMA_reg_buffer_3233_s_current_state_reg ( .D(
        new_AGEMA_signal_5120), .CK(clk), .Q(new_AGEMA_signal_5121) );
  DFF_X1 new_AGEMA_reg_buffer_3237_s_current_state_reg ( .D(
        new_AGEMA_signal_5124), .CK(clk), .Q(new_AGEMA_signal_5125) );
  DFF_X1 new_AGEMA_reg_buffer_3241_s_current_state_reg ( .D(
        new_AGEMA_signal_5128), .CK(clk), .Q(new_AGEMA_signal_5129) );
  DFF_X1 new_AGEMA_reg_buffer_3245_s_current_state_reg ( .D(
        new_AGEMA_signal_5132), .CK(clk), .Q(new_AGEMA_signal_5133) );
  DFF_X1 new_AGEMA_reg_buffer_3249_s_current_state_reg ( .D(
        new_AGEMA_signal_5136), .CK(clk), .Q(new_AGEMA_signal_5137) );
  DFF_X1 new_AGEMA_reg_buffer_3253_s_current_state_reg ( .D(
        new_AGEMA_signal_5140), .CK(clk), .Q(new_AGEMA_signal_5141) );
  DFF_X1 new_AGEMA_reg_buffer_3257_s_current_state_reg ( .D(
        new_AGEMA_signal_5144), .CK(clk), .Q(new_AGEMA_signal_5145) );
  DFF_X1 new_AGEMA_reg_buffer_3261_s_current_state_reg ( .D(
        new_AGEMA_signal_5148), .CK(clk), .Q(new_AGEMA_signal_5149) );
  DFF_X1 new_AGEMA_reg_buffer_3265_s_current_state_reg ( .D(
        new_AGEMA_signal_5152), .CK(clk), .Q(new_AGEMA_signal_5153) );
  DFF_X1 new_AGEMA_reg_buffer_3269_s_current_state_reg ( .D(
        new_AGEMA_signal_5156), .CK(clk), .Q(new_AGEMA_signal_5157) );
  DFF_X1 new_AGEMA_reg_buffer_3273_s_current_state_reg ( .D(
        new_AGEMA_signal_5160), .CK(clk), .Q(new_AGEMA_signal_5161) );
  DFF_X1 new_AGEMA_reg_buffer_3277_s_current_state_reg ( .D(
        new_AGEMA_signal_5164), .CK(clk), .Q(new_AGEMA_signal_5165) );
  DFF_X1 new_AGEMA_reg_buffer_3281_s_current_state_reg ( .D(
        new_AGEMA_signal_5168), .CK(clk), .Q(new_AGEMA_signal_5169) );
  DFF_X1 new_AGEMA_reg_buffer_3285_s_current_state_reg ( .D(
        new_AGEMA_signal_5172), .CK(clk), .Q(new_AGEMA_signal_5173) );
  DFF_X1 new_AGEMA_reg_buffer_3289_s_current_state_reg ( .D(
        new_AGEMA_signal_5176), .CK(clk), .Q(new_AGEMA_signal_5177) );
  DFF_X1 new_AGEMA_reg_buffer_3293_s_current_state_reg ( .D(
        new_AGEMA_signal_5180), .CK(clk), .Q(new_AGEMA_signal_5181) );
  DFF_X1 new_AGEMA_reg_buffer_3297_s_current_state_reg ( .D(
        new_AGEMA_signal_5184), .CK(clk), .Q(new_AGEMA_signal_5185) );
  DFF_X1 new_AGEMA_reg_buffer_3301_s_current_state_reg ( .D(
        new_AGEMA_signal_5188), .CK(clk), .Q(new_AGEMA_signal_5189) );
  DFF_X1 new_AGEMA_reg_buffer_3305_s_current_state_reg ( .D(
        new_AGEMA_signal_5192), .CK(clk), .Q(new_AGEMA_signal_5193) );
  DFF_X1 new_AGEMA_reg_buffer_3309_s_current_state_reg ( .D(
        new_AGEMA_signal_5196), .CK(clk), .Q(new_AGEMA_signal_5197) );
  DFF_X1 new_AGEMA_reg_buffer_3313_s_current_state_reg ( .D(
        new_AGEMA_signal_5200), .CK(clk), .Q(new_AGEMA_signal_5201) );
  DFF_X1 new_AGEMA_reg_buffer_3317_s_current_state_reg ( .D(
        new_AGEMA_signal_5204), .CK(clk), .Q(new_AGEMA_signal_5205) );
  DFF_X1 new_AGEMA_reg_buffer_3321_s_current_state_reg ( .D(
        new_AGEMA_signal_5208), .CK(clk), .Q(new_AGEMA_signal_5209) );
  DFF_X1 new_AGEMA_reg_buffer_3325_s_current_state_reg ( .D(
        new_AGEMA_signal_5212), .CK(clk), .Q(new_AGEMA_signal_5213) );
  DFF_X1 new_AGEMA_reg_buffer_3329_s_current_state_reg ( .D(
        new_AGEMA_signal_5216), .CK(clk), .Q(new_AGEMA_signal_5217) );
  DFF_X1 new_AGEMA_reg_buffer_3333_s_current_state_reg ( .D(
        new_AGEMA_signal_5220), .CK(clk), .Q(new_AGEMA_signal_5221) );
  DFF_X1 new_AGEMA_reg_buffer_3337_s_current_state_reg ( .D(
        new_AGEMA_signal_5224), .CK(clk), .Q(new_AGEMA_signal_5225) );
  DFF_X1 new_AGEMA_reg_buffer_3341_s_current_state_reg ( .D(
        new_AGEMA_signal_5228), .CK(clk), .Q(new_AGEMA_signal_5229) );
  DFF_X1 new_AGEMA_reg_buffer_3345_s_current_state_reg ( .D(
        new_AGEMA_signal_5232), .CK(clk), .Q(new_AGEMA_signal_5233) );
  DFF_X1 new_AGEMA_reg_buffer_3349_s_current_state_reg ( .D(
        new_AGEMA_signal_5236), .CK(clk), .Q(new_AGEMA_signal_5237) );
  DFF_X1 new_AGEMA_reg_buffer_3353_s_current_state_reg ( .D(
        new_AGEMA_signal_5240), .CK(clk), .Q(new_AGEMA_signal_5241) );
  DFF_X1 new_AGEMA_reg_buffer_3357_s_current_state_reg ( .D(
        new_AGEMA_signal_5244), .CK(clk), .Q(new_AGEMA_signal_5245) );
  DFF_X1 new_AGEMA_reg_buffer_3361_s_current_state_reg ( .D(
        new_AGEMA_signal_5248), .CK(clk), .Q(new_AGEMA_signal_5249) );
  DFF_X1 new_AGEMA_reg_buffer_3365_s_current_state_reg ( .D(
        new_AGEMA_signal_5252), .CK(clk), .Q(new_AGEMA_signal_5253) );
  DFF_X1 new_AGEMA_reg_buffer_3369_s_current_state_reg ( .D(
        new_AGEMA_signal_5256), .CK(clk), .Q(new_AGEMA_signal_5257) );
  DFF_X1 new_AGEMA_reg_buffer_3373_s_current_state_reg ( .D(
        new_AGEMA_signal_5260), .CK(clk), .Q(new_AGEMA_signal_5261) );
  DFF_X1 new_AGEMA_reg_buffer_3377_s_current_state_reg ( .D(
        new_AGEMA_signal_5264), .CK(clk), .Q(new_AGEMA_signal_5265) );
  DFF_X1 new_AGEMA_reg_buffer_3381_s_current_state_reg ( .D(
        new_AGEMA_signal_5268), .CK(clk), .Q(new_AGEMA_signal_5269) );
  DFF_X1 new_AGEMA_reg_buffer_3385_s_current_state_reg ( .D(
        new_AGEMA_signal_5272), .CK(clk), .Q(new_AGEMA_signal_5273) );
  DFF_X1 new_AGEMA_reg_buffer_3389_s_current_state_reg ( .D(
        new_AGEMA_signal_5276), .CK(clk), .Q(new_AGEMA_signal_5277) );
  DFF_X1 new_AGEMA_reg_buffer_3393_s_current_state_reg ( .D(
        new_AGEMA_signal_5280), .CK(clk), .Q(new_AGEMA_signal_5281) );
  DFF_X1 new_AGEMA_reg_buffer_3397_s_current_state_reg ( .D(
        new_AGEMA_signal_5284), .CK(clk), .Q(new_AGEMA_signal_5285) );
  DFF_X1 new_AGEMA_reg_buffer_3401_s_current_state_reg ( .D(
        new_AGEMA_signal_5288), .CK(clk), .Q(new_AGEMA_signal_5289) );
  DFF_X1 new_AGEMA_reg_buffer_3405_s_current_state_reg ( .D(
        new_AGEMA_signal_5292), .CK(clk), .Q(new_AGEMA_signal_5293) );
  DFF_X1 new_AGEMA_reg_buffer_3409_s_current_state_reg ( .D(
        new_AGEMA_signal_5296), .CK(clk), .Q(new_AGEMA_signal_5297) );
  DFF_X1 new_AGEMA_reg_buffer_3413_s_current_state_reg ( .D(
        new_AGEMA_signal_5300), .CK(clk), .Q(new_AGEMA_signal_5301) );
  DFF_X1 new_AGEMA_reg_buffer_3417_s_current_state_reg ( .D(
        new_AGEMA_signal_5304), .CK(clk), .Q(new_AGEMA_signal_5305) );
  DFF_X1 new_AGEMA_reg_buffer_3421_s_current_state_reg ( .D(
        new_AGEMA_signal_5308), .CK(clk), .Q(new_AGEMA_signal_5309) );
  DFF_X1 new_AGEMA_reg_buffer_3425_s_current_state_reg ( .D(
        new_AGEMA_signal_5312), .CK(clk), .Q(new_AGEMA_signal_5313) );
  DFF_X1 new_AGEMA_reg_buffer_3429_s_current_state_reg ( .D(
        new_AGEMA_signal_5316), .CK(clk), .Q(new_AGEMA_signal_5317) );
  DFF_X1 new_AGEMA_reg_buffer_3433_s_current_state_reg ( .D(
        new_AGEMA_signal_5320), .CK(clk), .Q(new_AGEMA_signal_5321) );
  DFF_X1 new_AGEMA_reg_buffer_3437_s_current_state_reg ( .D(
        new_AGEMA_signal_5324), .CK(clk), .Q(new_AGEMA_signal_5325) );
  DFF_X1 new_AGEMA_reg_buffer_3441_s_current_state_reg ( .D(
        new_AGEMA_signal_5328), .CK(clk), .Q(new_AGEMA_signal_5329) );
  DFF_X1 new_AGEMA_reg_buffer_3445_s_current_state_reg ( .D(
        new_AGEMA_signal_5332), .CK(clk), .Q(new_AGEMA_signal_5333) );
  DFF_X1 new_AGEMA_reg_buffer_3449_s_current_state_reg ( .D(
        new_AGEMA_signal_5336), .CK(clk), .Q(new_AGEMA_signal_5337) );
  DFF_X1 new_AGEMA_reg_buffer_3453_s_current_state_reg ( .D(
        new_AGEMA_signal_5340), .CK(clk), .Q(new_AGEMA_signal_5341) );
  DFF_X1 new_AGEMA_reg_buffer_3457_s_current_state_reg ( .D(
        new_AGEMA_signal_5344), .CK(clk), .Q(new_AGEMA_signal_5345) );
  DFF_X1 new_AGEMA_reg_buffer_3461_s_current_state_reg ( .D(
        new_AGEMA_signal_5348), .CK(clk), .Q(new_AGEMA_signal_5349) );
  DFF_X1 new_AGEMA_reg_buffer_3465_s_current_state_reg ( .D(
        new_AGEMA_signal_5352), .CK(clk), .Q(new_AGEMA_signal_5353) );
  DFF_X1 new_AGEMA_reg_buffer_3469_s_current_state_reg ( .D(
        new_AGEMA_signal_5356), .CK(clk), .Q(new_AGEMA_signal_5357) );
  DFF_X1 new_AGEMA_reg_buffer_3473_s_current_state_reg ( .D(
        new_AGEMA_signal_5360), .CK(clk), .Q(new_AGEMA_signal_5361) );
  DFF_X1 new_AGEMA_reg_buffer_3477_s_current_state_reg ( .D(
        new_AGEMA_signal_5364), .CK(clk), .Q(new_AGEMA_signal_5365) );
  DFF_X1 new_AGEMA_reg_buffer_3481_s_current_state_reg ( .D(
        new_AGEMA_signal_5368), .CK(clk), .Q(new_AGEMA_signal_5369) );
  DFF_X1 new_AGEMA_reg_buffer_3485_s_current_state_reg ( .D(
        new_AGEMA_signal_5372), .CK(clk), .Q(new_AGEMA_signal_5373) );
  DFF_X1 new_AGEMA_reg_buffer_3489_s_current_state_reg ( .D(
        new_AGEMA_signal_5376), .CK(clk), .Q(new_AGEMA_signal_5377) );
  DFF_X1 new_AGEMA_reg_buffer_3493_s_current_state_reg ( .D(
        new_AGEMA_signal_5380), .CK(clk), .Q(new_AGEMA_signal_5381) );
  DFF_X1 new_AGEMA_reg_buffer_3497_s_current_state_reg ( .D(
        new_AGEMA_signal_5384), .CK(clk), .Q(new_AGEMA_signal_5385) );
  DFF_X1 new_AGEMA_reg_buffer_3501_s_current_state_reg ( .D(
        new_AGEMA_signal_5388), .CK(clk), .Q(new_AGEMA_signal_5389) );
  DFF_X1 new_AGEMA_reg_buffer_3505_s_current_state_reg ( .D(
        new_AGEMA_signal_5392), .CK(clk), .Q(new_AGEMA_signal_5393) );
  DFF_X1 new_AGEMA_reg_buffer_3509_s_current_state_reg ( .D(
        new_AGEMA_signal_5396), .CK(clk), .Q(new_AGEMA_signal_5397) );
  DFF_X1 new_AGEMA_reg_buffer_3513_s_current_state_reg ( .D(
        new_AGEMA_signal_5400), .CK(clk), .Q(new_AGEMA_signal_5401) );
  DFF_X1 new_AGEMA_reg_buffer_3517_s_current_state_reg ( .D(
        new_AGEMA_signal_5404), .CK(clk), .Q(new_AGEMA_signal_5405) );
  DFF_X1 new_AGEMA_reg_buffer_3521_s_current_state_reg ( .D(
        new_AGEMA_signal_5408), .CK(clk), .Q(new_AGEMA_signal_5409) );
  DFF_X1 new_AGEMA_reg_buffer_3525_s_current_state_reg ( .D(
        new_AGEMA_signal_5412), .CK(clk), .Q(new_AGEMA_signal_5413) );
  DFF_X1 new_AGEMA_reg_buffer_3529_s_current_state_reg ( .D(
        new_AGEMA_signal_5416), .CK(clk), .Q(new_AGEMA_signal_5417) );
  DFF_X1 new_AGEMA_reg_buffer_3533_s_current_state_reg ( .D(
        new_AGEMA_signal_5420), .CK(clk), .Q(new_AGEMA_signal_5421) );
  DFF_X1 new_AGEMA_reg_buffer_3537_s_current_state_reg ( .D(
        new_AGEMA_signal_5424), .CK(clk), .Q(new_AGEMA_signal_5425) );
  DFF_X1 new_AGEMA_reg_buffer_3541_s_current_state_reg ( .D(
        new_AGEMA_signal_5428), .CK(clk), .Q(new_AGEMA_signal_5429) );
  DFF_X1 new_AGEMA_reg_buffer_3545_s_current_state_reg ( .D(
        new_AGEMA_signal_5432), .CK(clk), .Q(new_AGEMA_signal_5433) );
  DFF_X1 new_AGEMA_reg_buffer_3549_s_current_state_reg ( .D(
        new_AGEMA_signal_5436), .CK(clk), .Q(new_AGEMA_signal_5437) );
  DFF_X1 new_AGEMA_reg_buffer_3553_s_current_state_reg ( .D(
        new_AGEMA_signal_5440), .CK(clk), .Q(new_AGEMA_signal_5441) );
  DFF_X1 new_AGEMA_reg_buffer_3557_s_current_state_reg ( .D(
        new_AGEMA_signal_5444), .CK(clk), .Q(new_AGEMA_signal_5445) );
  DFF_X1 new_AGEMA_reg_buffer_3561_s_current_state_reg ( .D(
        new_AGEMA_signal_5448), .CK(clk), .Q(new_AGEMA_signal_5449) );
  DFF_X1 new_AGEMA_reg_buffer_3565_s_current_state_reg ( .D(
        new_AGEMA_signal_5452), .CK(clk), .Q(new_AGEMA_signal_5453) );
  DFF_X1 new_AGEMA_reg_buffer_3569_s_current_state_reg ( .D(
        new_AGEMA_signal_5456), .CK(clk), .Q(new_AGEMA_signal_5457) );
  DFF_X1 new_AGEMA_reg_buffer_3573_s_current_state_reg ( .D(
        new_AGEMA_signal_5460), .CK(clk), .Q(new_AGEMA_signal_5461) );
  DFF_X1 new_AGEMA_reg_buffer_3577_s_current_state_reg ( .D(
        new_AGEMA_signal_5464), .CK(clk), .Q(new_AGEMA_signal_5465) );
  DFF_X1 new_AGEMA_reg_buffer_3581_s_current_state_reg ( .D(
        new_AGEMA_signal_5468), .CK(clk), .Q(new_AGEMA_signal_5469) );
  DFF_X1 new_AGEMA_reg_buffer_3585_s_current_state_reg ( .D(
        new_AGEMA_signal_5472), .CK(clk), .Q(new_AGEMA_signal_5473) );
  DFF_X1 new_AGEMA_reg_buffer_3589_s_current_state_reg ( .D(
        new_AGEMA_signal_5476), .CK(clk), .Q(new_AGEMA_signal_5477) );
  DFF_X1 new_AGEMA_reg_buffer_3593_s_current_state_reg ( .D(
        new_AGEMA_signal_5480), .CK(clk), .Q(new_AGEMA_signal_5481) );
  DFF_X1 new_AGEMA_reg_buffer_3597_s_current_state_reg ( .D(
        new_AGEMA_signal_5484), .CK(clk), .Q(new_AGEMA_signal_5485) );
  DFF_X1 new_AGEMA_reg_buffer_3601_s_current_state_reg ( .D(
        new_AGEMA_signal_5488), .CK(clk), .Q(new_AGEMA_signal_5489) );
  DFF_X1 new_AGEMA_reg_buffer_3605_s_current_state_reg ( .D(
        new_AGEMA_signal_5492), .CK(clk), .Q(new_AGEMA_signal_5493) );
  DFF_X1 new_AGEMA_reg_buffer_3609_s_current_state_reg ( .D(
        new_AGEMA_signal_5496), .CK(clk), .Q(new_AGEMA_signal_5497) );
  DFF_X1 new_AGEMA_reg_buffer_3613_s_current_state_reg ( .D(
        new_AGEMA_signal_5500), .CK(clk), .Q(new_AGEMA_signal_5501) );
  DFF_X1 new_AGEMA_reg_buffer_3617_s_current_state_reg ( .D(
        new_AGEMA_signal_5504), .CK(clk), .Q(new_AGEMA_signal_5505) );
  DFF_X1 new_AGEMA_reg_buffer_3621_s_current_state_reg ( .D(
        new_AGEMA_signal_5508), .CK(clk), .Q(new_AGEMA_signal_5509) );
  DFF_X1 new_AGEMA_reg_buffer_3625_s_current_state_reg ( .D(
        new_AGEMA_signal_5512), .CK(clk), .Q(new_AGEMA_signal_5513) );
  DFF_X1 new_AGEMA_reg_buffer_3629_s_current_state_reg ( .D(
        new_AGEMA_signal_5516), .CK(clk), .Q(new_AGEMA_signal_5517) );
  DFF_X1 new_AGEMA_reg_buffer_3633_s_current_state_reg ( .D(
        new_AGEMA_signal_5520), .CK(clk), .Q(new_AGEMA_signal_5521) );
  DFF_X1 new_AGEMA_reg_buffer_3637_s_current_state_reg ( .D(
        new_AGEMA_signal_5524), .CK(clk), .Q(new_AGEMA_signal_5525) );
  DFF_X1 new_AGEMA_reg_buffer_3641_s_current_state_reg ( .D(
        new_AGEMA_signal_5528), .CK(clk), .Q(new_AGEMA_signal_5529) );
  DFF_X1 new_AGEMA_reg_buffer_3645_s_current_state_reg ( .D(
        new_AGEMA_signal_5532), .CK(clk), .Q(new_AGEMA_signal_5533) );
  DFF_X1 new_AGEMA_reg_buffer_3649_s_current_state_reg ( .D(
        new_AGEMA_signal_5536), .CK(clk), .Q(new_AGEMA_signal_5537) );
  DFF_X1 new_AGEMA_reg_buffer_3653_s_current_state_reg ( .D(
        new_AGEMA_signal_5540), .CK(clk), .Q(new_AGEMA_signal_5541) );
  DFF_X1 new_AGEMA_reg_buffer_3657_s_current_state_reg ( .D(
        new_AGEMA_signal_5544), .CK(clk), .Q(new_AGEMA_signal_5545) );
  DFF_X1 new_AGEMA_reg_buffer_3661_s_current_state_reg ( .D(
        new_AGEMA_signal_5548), .CK(clk), .Q(new_AGEMA_signal_5549) );
  DFF_X1 new_AGEMA_reg_buffer_3665_s_current_state_reg ( .D(
        new_AGEMA_signal_5552), .CK(clk), .Q(new_AGEMA_signal_5553) );
  DFF_X1 new_AGEMA_reg_buffer_3669_s_current_state_reg ( .D(
        new_AGEMA_signal_5556), .CK(clk), .Q(new_AGEMA_signal_5557) );
  DFF_X1 new_AGEMA_reg_buffer_3673_s_current_state_reg ( .D(
        new_AGEMA_signal_5560), .CK(clk), .Q(new_AGEMA_signal_5561) );
  DFF_X1 new_AGEMA_reg_buffer_3677_s_current_state_reg ( .D(
        new_AGEMA_signal_5564), .CK(clk), .Q(new_AGEMA_signal_5565) );
  DFF_X1 new_AGEMA_reg_buffer_3681_s_current_state_reg ( .D(
        new_AGEMA_signal_5568), .CK(clk), .Q(new_AGEMA_signal_5569) );
  DFF_X1 new_AGEMA_reg_buffer_3685_s_current_state_reg ( .D(
        new_AGEMA_signal_5572), .CK(clk), .Q(new_AGEMA_signal_5573) );
  DFF_X1 new_AGEMA_reg_buffer_3689_s_current_state_reg ( .D(
        new_AGEMA_signal_5576), .CK(clk), .Q(new_AGEMA_signal_5577) );
  DFF_X1 new_AGEMA_reg_buffer_3693_s_current_state_reg ( .D(
        new_AGEMA_signal_5580), .CK(clk), .Q(new_AGEMA_signal_5581) );
  DFF_X1 new_AGEMA_reg_buffer_3697_s_current_state_reg ( .D(
        new_AGEMA_signal_5584), .CK(clk), .Q(new_AGEMA_signal_5585) );
  DFF_X1 new_AGEMA_reg_buffer_3701_s_current_state_reg ( .D(
        new_AGEMA_signal_5588), .CK(clk), .Q(new_AGEMA_signal_5589) );
  DFF_X1 new_AGEMA_reg_buffer_3705_s_current_state_reg ( .D(
        new_AGEMA_signal_5592), .CK(clk), .Q(new_AGEMA_signal_5593) );
  DFF_X1 new_AGEMA_reg_buffer_3709_s_current_state_reg ( .D(
        new_AGEMA_signal_5596), .CK(clk), .Q(new_AGEMA_signal_5597) );
  DFF_X1 new_AGEMA_reg_buffer_3713_s_current_state_reg ( .D(
        new_AGEMA_signal_5600), .CK(clk), .Q(new_AGEMA_signal_5601) );
  DFF_X1 new_AGEMA_reg_buffer_3717_s_current_state_reg ( .D(
        new_AGEMA_signal_5604), .CK(clk), .Q(new_AGEMA_signal_5605) );
  DFF_X1 new_AGEMA_reg_buffer_3721_s_current_state_reg ( .D(
        new_AGEMA_signal_5608), .CK(clk), .Q(new_AGEMA_signal_5609) );
  DFF_X1 new_AGEMA_reg_buffer_3725_s_current_state_reg ( .D(
        new_AGEMA_signal_5612), .CK(clk), .Q(new_AGEMA_signal_5613) );
  DFF_X1 new_AGEMA_reg_buffer_3729_s_current_state_reg ( .D(
        new_AGEMA_signal_5616), .CK(clk), .Q(new_AGEMA_signal_5617) );
  DFF_X1 new_AGEMA_reg_buffer_3733_s_current_state_reg ( .D(
        new_AGEMA_signal_5620), .CK(clk), .Q(new_AGEMA_signal_5621) );
  DFF_X1 new_AGEMA_reg_buffer_3737_s_current_state_reg ( .D(
        new_AGEMA_signal_5624), .CK(clk), .Q(new_AGEMA_signal_5625) );
  DFF_X1 new_AGEMA_reg_buffer_3741_s_current_state_reg ( .D(
        new_AGEMA_signal_5628), .CK(clk), .Q(new_AGEMA_signal_5629) );
  DFF_X1 new_AGEMA_reg_buffer_3745_s_current_state_reg ( .D(
        new_AGEMA_signal_5632), .CK(clk), .Q(new_AGEMA_signal_5633) );
  DFF_X1 new_AGEMA_reg_buffer_3749_s_current_state_reg ( .D(
        new_AGEMA_signal_5636), .CK(clk), .Q(new_AGEMA_signal_5637) );
  DFF_X1 new_AGEMA_reg_buffer_3753_s_current_state_reg ( .D(
        new_AGEMA_signal_5640), .CK(clk), .Q(new_AGEMA_signal_5641) );
  DFF_X1 new_AGEMA_reg_buffer_3757_s_current_state_reg ( .D(
        new_AGEMA_signal_5644), .CK(clk), .Q(new_AGEMA_signal_5645) );
  DFF_X1 new_AGEMA_reg_buffer_3761_s_current_state_reg ( .D(
        new_AGEMA_signal_5648), .CK(clk), .Q(new_AGEMA_signal_5649) );
  DFF_X1 new_AGEMA_reg_buffer_3765_s_current_state_reg ( .D(
        new_AGEMA_signal_5652), .CK(clk), .Q(new_AGEMA_signal_5653) );
  DFF_X1 new_AGEMA_reg_buffer_3769_s_current_state_reg ( .D(
        new_AGEMA_signal_5656), .CK(clk), .Q(new_AGEMA_signal_5657) );
  DFF_X1 new_AGEMA_reg_buffer_3773_s_current_state_reg ( .D(
        new_AGEMA_signal_5660), .CK(clk), .Q(new_AGEMA_signal_5661) );
  DFF_X1 new_AGEMA_reg_buffer_3777_s_current_state_reg ( .D(
        new_AGEMA_signal_5664), .CK(clk), .Q(new_AGEMA_signal_5665) );
  DFF_X1 new_AGEMA_reg_buffer_3781_s_current_state_reg ( .D(
        new_AGEMA_signal_5668), .CK(clk), .Q(new_AGEMA_signal_5669) );
  DFF_X1 new_AGEMA_reg_buffer_3785_s_current_state_reg ( .D(
        new_AGEMA_signal_5672), .CK(clk), .Q(new_AGEMA_signal_5673) );
  DFF_X1 new_AGEMA_reg_buffer_3789_s_current_state_reg ( .D(
        new_AGEMA_signal_5676), .CK(clk), .Q(new_AGEMA_signal_5677) );
  DFF_X1 new_AGEMA_reg_buffer_3793_s_current_state_reg ( .D(
        new_AGEMA_signal_5680), .CK(clk), .Q(new_AGEMA_signal_5681) );
  DFF_X1 new_AGEMA_reg_buffer_3797_s_current_state_reg ( .D(
        new_AGEMA_signal_5684), .CK(clk), .Q(new_AGEMA_signal_5685) );
  DFF_X1 new_AGEMA_reg_buffer_3801_s_current_state_reg ( .D(
        new_AGEMA_signal_5688), .CK(clk), .Q(new_AGEMA_signal_5689) );
  DFF_X1 new_AGEMA_reg_buffer_3805_s_current_state_reg ( .D(
        new_AGEMA_signal_5692), .CK(clk), .Q(new_AGEMA_signal_5693) );
  DFF_X1 new_AGEMA_reg_buffer_3809_s_current_state_reg ( .D(
        new_AGEMA_signal_5696), .CK(clk), .Q(new_AGEMA_signal_5697) );
  DFF_X1 new_AGEMA_reg_buffer_3813_s_current_state_reg ( .D(
        new_AGEMA_signal_5700), .CK(clk), .Q(new_AGEMA_signal_5701) );
  DFF_X1 new_AGEMA_reg_buffer_3817_s_current_state_reg ( .D(
        new_AGEMA_signal_5704), .CK(clk), .Q(new_AGEMA_signal_5705) );
  DFF_X1 new_AGEMA_reg_buffer_3821_s_current_state_reg ( .D(
        new_AGEMA_signal_5708), .CK(clk), .Q(new_AGEMA_signal_5709) );
  DFF_X1 new_AGEMA_reg_buffer_3825_s_current_state_reg ( .D(
        new_AGEMA_signal_5712), .CK(clk), .Q(new_AGEMA_signal_5713) );
  DFF_X1 new_AGEMA_reg_buffer_3829_s_current_state_reg ( .D(
        new_AGEMA_signal_5716), .CK(clk), .Q(new_AGEMA_signal_5717) );
  DFF_X1 new_AGEMA_reg_buffer_3833_s_current_state_reg ( .D(
        new_AGEMA_signal_5720), .CK(clk), .Q(new_AGEMA_signal_5721) );
  DFF_X1 new_AGEMA_reg_buffer_3837_s_current_state_reg ( .D(
        new_AGEMA_signal_5724), .CK(clk), .Q(new_AGEMA_signal_5725) );
  DFF_X1 new_AGEMA_reg_buffer_3841_s_current_state_reg ( .D(
        new_AGEMA_signal_5728), .CK(clk), .Q(new_AGEMA_signal_5729) );
  DFF_X1 new_AGEMA_reg_buffer_3845_s_current_state_reg ( .D(
        new_AGEMA_signal_5732), .CK(clk), .Q(new_AGEMA_signal_5733) );
  DFF_X1 new_AGEMA_reg_buffer_3849_s_current_state_reg ( .D(
        new_AGEMA_signal_5736), .CK(clk), .Q(new_AGEMA_signal_5737) );
  DFF_X1 new_AGEMA_reg_buffer_3853_s_current_state_reg ( .D(
        new_AGEMA_signal_5740), .CK(clk), .Q(new_AGEMA_signal_5741) );
  DFF_X1 new_AGEMA_reg_buffer_3857_s_current_state_reg ( .D(
        new_AGEMA_signal_5744), .CK(clk), .Q(new_AGEMA_signal_5745) );
  DFF_X1 new_AGEMA_reg_buffer_3861_s_current_state_reg ( .D(
        new_AGEMA_signal_5748), .CK(clk), .Q(new_AGEMA_signal_5749) );
  DFF_X1 new_AGEMA_reg_buffer_3865_s_current_state_reg ( .D(
        new_AGEMA_signal_5752), .CK(clk), .Q(new_AGEMA_signal_5753) );
  DFF_X1 new_AGEMA_reg_buffer_3869_s_current_state_reg ( .D(
        new_AGEMA_signal_5756), .CK(clk), .Q(new_AGEMA_signal_5757) );
  DFF_X1 new_AGEMA_reg_buffer_3873_s_current_state_reg ( .D(
        new_AGEMA_signal_5760), .CK(clk), .Q(new_AGEMA_signal_5761) );
  DFF_X1 new_AGEMA_reg_buffer_3877_s_current_state_reg ( .D(
        new_AGEMA_signal_5764), .CK(clk), .Q(new_AGEMA_signal_5765) );
  DFF_X1 new_AGEMA_reg_buffer_3881_s_current_state_reg ( .D(
        new_AGEMA_signal_5768), .CK(clk), .Q(new_AGEMA_signal_5769) );
  DFF_X1 new_AGEMA_reg_buffer_3885_s_current_state_reg ( .D(
        new_AGEMA_signal_5772), .CK(clk), .Q(new_AGEMA_signal_5773) );
  DFF_X1 new_AGEMA_reg_buffer_3889_s_current_state_reg ( .D(
        new_AGEMA_signal_5776), .CK(clk), .Q(new_AGEMA_signal_5777) );
  DFF_X1 new_AGEMA_reg_buffer_3893_s_current_state_reg ( .D(
        new_AGEMA_signal_5780), .CK(clk), .Q(new_AGEMA_signal_5781) );
  DFF_X1 new_AGEMA_reg_buffer_3897_s_current_state_reg ( .D(
        new_AGEMA_signal_5784), .CK(clk), .Q(new_AGEMA_signal_5785) );
  DFF_X1 new_AGEMA_reg_buffer_3901_s_current_state_reg ( .D(
        new_AGEMA_signal_5788), .CK(clk), .Q(new_AGEMA_signal_5789) );
  DFF_X1 new_AGEMA_reg_buffer_3905_s_current_state_reg ( .D(
        new_AGEMA_signal_5792), .CK(clk), .Q(new_AGEMA_signal_5793) );
  DFF_X1 new_AGEMA_reg_buffer_3909_s_current_state_reg ( .D(
        new_AGEMA_signal_5796), .CK(clk), .Q(new_AGEMA_signal_5797) );
  DFF_X1 new_AGEMA_reg_buffer_3913_s_current_state_reg ( .D(
        new_AGEMA_signal_5800), .CK(clk), .Q(new_AGEMA_signal_5801) );
  DFF_X1 new_AGEMA_reg_buffer_3917_s_current_state_reg ( .D(
        new_AGEMA_signal_5804), .CK(clk), .Q(new_AGEMA_signal_5805) );
  DFF_X1 new_AGEMA_reg_buffer_3921_s_current_state_reg ( .D(
        new_AGEMA_signal_5808), .CK(clk), .Q(new_AGEMA_signal_5809) );
  DFF_X1 new_AGEMA_reg_buffer_3925_s_current_state_reg ( .D(
        new_AGEMA_signal_5812), .CK(clk), .Q(new_AGEMA_signal_5813) );
  DFF_X1 new_AGEMA_reg_buffer_3929_s_current_state_reg ( .D(
        new_AGEMA_signal_5816), .CK(clk), .Q(new_AGEMA_signal_5817) );
  DFF_X1 new_AGEMA_reg_buffer_3933_s_current_state_reg ( .D(
        new_AGEMA_signal_5820), .CK(clk), .Q(new_AGEMA_signal_5821) );
  DFF_X1 new_AGEMA_reg_buffer_3937_s_current_state_reg ( .D(
        new_AGEMA_signal_5824), .CK(clk), .Q(new_AGEMA_signal_5825) );
  DFF_X1 new_AGEMA_reg_buffer_3941_s_current_state_reg ( .D(
        new_AGEMA_signal_5828), .CK(clk), .Q(new_AGEMA_signal_5829) );
  DFF_X1 new_AGEMA_reg_buffer_3945_s_current_state_reg ( .D(
        new_AGEMA_signal_5832), .CK(clk), .Q(new_AGEMA_signal_5833) );
  DFF_X1 new_AGEMA_reg_buffer_3949_s_current_state_reg ( .D(
        new_AGEMA_signal_5836), .CK(clk), .Q(new_AGEMA_signal_5837) );
  DFF_X1 new_AGEMA_reg_buffer_3953_s_current_state_reg ( .D(
        new_AGEMA_signal_5840), .CK(clk), .Q(new_AGEMA_signal_5841) );
  DFF_X1 new_AGEMA_reg_buffer_3957_s_current_state_reg ( .D(
        new_AGEMA_signal_5844), .CK(clk), .Q(new_AGEMA_signal_5845) );
  DFF_X1 new_AGEMA_reg_buffer_3961_s_current_state_reg ( .D(
        new_AGEMA_signal_5848), .CK(clk), .Q(new_AGEMA_signal_5849) );
  DFF_X1 new_AGEMA_reg_buffer_3965_s_current_state_reg ( .D(
        new_AGEMA_signal_5852), .CK(clk), .Q(new_AGEMA_signal_5853) );
  DFF_X1 new_AGEMA_reg_buffer_3969_s_current_state_reg ( .D(
        new_AGEMA_signal_5856), .CK(clk), .Q(new_AGEMA_signal_5857) );
  DFF_X1 new_AGEMA_reg_buffer_3973_s_current_state_reg ( .D(
        new_AGEMA_signal_5860), .CK(clk), .Q(new_AGEMA_signal_5861) );
  DFF_X1 new_AGEMA_reg_buffer_3977_s_current_state_reg ( .D(
        new_AGEMA_signal_5864), .CK(clk), .Q(new_AGEMA_signal_5865) );
  DFF_X1 new_AGEMA_reg_buffer_3981_s_current_state_reg ( .D(
        new_AGEMA_signal_5868), .CK(clk), .Q(new_AGEMA_signal_5869) );
  DFF_X1 new_AGEMA_reg_buffer_3985_s_current_state_reg ( .D(
        new_AGEMA_signal_5872), .CK(clk), .Q(new_AGEMA_signal_5873) );
  DFF_X1 new_AGEMA_reg_buffer_3989_s_current_state_reg ( .D(
        new_AGEMA_signal_5876), .CK(clk), .Q(new_AGEMA_signal_5877) );
  DFF_X1 new_AGEMA_reg_buffer_3993_s_current_state_reg ( .D(
        new_AGEMA_signal_5880), .CK(clk), .Q(new_AGEMA_signal_5881) );
  DFF_X1 new_AGEMA_reg_buffer_3997_s_current_state_reg ( .D(
        new_AGEMA_signal_5884), .CK(clk), .Q(new_AGEMA_signal_5885) );
  DFF_X1 new_AGEMA_reg_buffer_4001_s_current_state_reg ( .D(
        new_AGEMA_signal_5888), .CK(clk), .Q(new_AGEMA_signal_5889) );
  DFF_X1 new_AGEMA_reg_buffer_4005_s_current_state_reg ( .D(
        new_AGEMA_signal_5892), .CK(clk), .Q(new_AGEMA_signal_5893) );
  DFF_X1 new_AGEMA_reg_buffer_4009_s_current_state_reg ( .D(
        new_AGEMA_signal_5896), .CK(clk), .Q(new_AGEMA_signal_5897) );
  DFF_X1 new_AGEMA_reg_buffer_4013_s_current_state_reg ( .D(
        new_AGEMA_signal_5900), .CK(clk), .Q(new_AGEMA_signal_5901) );
  DFF_X1 new_AGEMA_reg_buffer_4017_s_current_state_reg ( .D(
        new_AGEMA_signal_5904), .CK(clk), .Q(new_AGEMA_signal_5905) );
  DFF_X1 new_AGEMA_reg_buffer_4021_s_current_state_reg ( .D(
        new_AGEMA_signal_5908), .CK(clk), .Q(new_AGEMA_signal_5909) );
  DFF_X1 new_AGEMA_reg_buffer_4025_s_current_state_reg ( .D(
        new_AGEMA_signal_5912), .CK(clk), .Q(new_AGEMA_signal_5913) );
  DFF_X1 new_AGEMA_reg_buffer_4029_s_current_state_reg ( .D(
        new_AGEMA_signal_5916), .CK(clk), .Q(new_AGEMA_signal_5917) );
  DFF_X1 new_AGEMA_reg_buffer_4033_s_current_state_reg ( .D(
        new_AGEMA_signal_5920), .CK(clk), .Q(new_AGEMA_signal_5921) );
  DFF_X1 new_AGEMA_reg_buffer_4037_s_current_state_reg ( .D(
        new_AGEMA_signal_5924), .CK(clk), .Q(new_AGEMA_signal_5925) );
  DFF_X1 new_AGEMA_reg_buffer_4041_s_current_state_reg ( .D(
        new_AGEMA_signal_5928), .CK(clk), .Q(new_AGEMA_signal_5929) );
  DFF_X1 new_AGEMA_reg_buffer_4045_s_current_state_reg ( .D(
        new_AGEMA_signal_5932), .CK(clk), .Q(new_AGEMA_signal_5933) );
  DFF_X1 new_AGEMA_reg_buffer_4049_s_current_state_reg ( .D(
        new_AGEMA_signal_5936), .CK(clk), .Q(new_AGEMA_signal_5937) );
  DFF_X1 new_AGEMA_reg_buffer_4053_s_current_state_reg ( .D(
        new_AGEMA_signal_5940), .CK(clk), .Q(new_AGEMA_signal_5941) );
  DFF_X1 new_AGEMA_reg_buffer_4057_s_current_state_reg ( .D(
        new_AGEMA_signal_5944), .CK(clk), .Q(new_AGEMA_signal_5945) );
  DFF_X1 new_AGEMA_reg_buffer_4061_s_current_state_reg ( .D(
        new_AGEMA_signal_5948), .CK(clk), .Q(new_AGEMA_signal_5949) );
  DFF_X1 new_AGEMA_reg_buffer_4065_s_current_state_reg ( .D(
        new_AGEMA_signal_5952), .CK(clk), .Q(new_AGEMA_signal_5953) );
  DFF_X1 new_AGEMA_reg_buffer_4069_s_current_state_reg ( .D(
        new_AGEMA_signal_5956), .CK(clk), .Q(new_AGEMA_signal_5957) );
  DFF_X1 new_AGEMA_reg_buffer_4073_s_current_state_reg ( .D(
        new_AGEMA_signal_5960), .CK(clk), .Q(new_AGEMA_signal_5961) );
  DFF_X1 new_AGEMA_reg_buffer_4077_s_current_state_reg ( .D(
        new_AGEMA_signal_5964), .CK(clk), .Q(new_AGEMA_signal_5965) );
  DFF_X1 new_AGEMA_reg_buffer_4081_s_current_state_reg ( .D(
        new_AGEMA_signal_5968), .CK(clk), .Q(new_AGEMA_signal_5969) );
  DFF_X1 new_AGEMA_reg_buffer_4085_s_current_state_reg ( .D(
        new_AGEMA_signal_5972), .CK(clk), .Q(new_AGEMA_signal_5973) );
  DFF_X1 new_AGEMA_reg_buffer_4089_s_current_state_reg ( .D(
        new_AGEMA_signal_5976), .CK(clk), .Q(new_AGEMA_signal_5977) );
  DFF_X1 new_AGEMA_reg_buffer_4093_s_current_state_reg ( .D(
        new_AGEMA_signal_5980), .CK(clk), .Q(new_AGEMA_signal_5981) );
  DFF_X1 new_AGEMA_reg_buffer_4097_s_current_state_reg ( .D(
        new_AGEMA_signal_5984), .CK(clk), .Q(new_AGEMA_signal_5985) );
  DFF_X1 new_AGEMA_reg_buffer_4101_s_current_state_reg ( .D(
        new_AGEMA_signal_5988), .CK(clk), .Q(new_AGEMA_signal_5989) );
  DFF_X1 new_AGEMA_reg_buffer_4105_s_current_state_reg ( .D(
        new_AGEMA_signal_5992), .CK(clk), .Q(new_AGEMA_signal_5993) );
  DFF_X1 new_AGEMA_reg_buffer_4109_s_current_state_reg ( .D(
        new_AGEMA_signal_5996), .CK(clk), .Q(new_AGEMA_signal_5997) );
  DFF_X1 new_AGEMA_reg_buffer_4113_s_current_state_reg ( .D(
        new_AGEMA_signal_6000), .CK(clk), .Q(new_AGEMA_signal_6001) );
  DFF_X1 new_AGEMA_reg_buffer_4117_s_current_state_reg ( .D(
        new_AGEMA_signal_6004), .CK(clk), .Q(new_AGEMA_signal_6005) );
  DFF_X1 new_AGEMA_reg_buffer_4121_s_current_state_reg ( .D(
        new_AGEMA_signal_6008), .CK(clk), .Q(new_AGEMA_signal_6009) );
  DFF_X1 new_AGEMA_reg_buffer_4125_s_current_state_reg ( .D(
        new_AGEMA_signal_6012), .CK(clk), .Q(new_AGEMA_signal_6013) );
  DFF_X1 new_AGEMA_reg_buffer_4129_s_current_state_reg ( .D(
        new_AGEMA_signal_6016), .CK(clk), .Q(new_AGEMA_signal_6017) );
  DFF_X1 new_AGEMA_reg_buffer_4133_s_current_state_reg ( .D(
        new_AGEMA_signal_6020), .CK(clk), .Q(new_AGEMA_signal_6021) );
  DFF_X1 new_AGEMA_reg_buffer_4137_s_current_state_reg ( .D(
        new_AGEMA_signal_6024), .CK(clk), .Q(new_AGEMA_signal_6025) );
  DFF_X1 new_AGEMA_reg_buffer_4141_s_current_state_reg ( .D(
        new_AGEMA_signal_6028), .CK(clk), .Q(new_AGEMA_signal_6029) );
  DFF_X1 new_AGEMA_reg_buffer_4145_s_current_state_reg ( .D(
        new_AGEMA_signal_6032), .CK(clk), .Q(new_AGEMA_signal_6033) );
  DFF_X1 new_AGEMA_reg_buffer_4149_s_current_state_reg ( .D(
        new_AGEMA_signal_6036), .CK(clk), .Q(new_AGEMA_signal_6037) );
  DFF_X1 new_AGEMA_reg_buffer_4153_s_current_state_reg ( .D(
        new_AGEMA_signal_6040), .CK(clk), .Q(new_AGEMA_signal_6041) );
  DFF_X1 new_AGEMA_reg_buffer_4157_s_current_state_reg ( .D(
        new_AGEMA_signal_6044), .CK(clk), .Q(new_AGEMA_signal_6045) );
  DFF_X1 new_AGEMA_reg_buffer_4161_s_current_state_reg ( .D(
        new_AGEMA_signal_6048), .CK(clk), .Q(new_AGEMA_signal_6049) );
  DFF_X1 new_AGEMA_reg_buffer_4165_s_current_state_reg ( .D(
        new_AGEMA_signal_6052), .CK(clk), .Q(new_AGEMA_signal_6053) );
  DFF_X1 new_AGEMA_reg_buffer_4169_s_current_state_reg ( .D(
        new_AGEMA_signal_6056), .CK(clk), .Q(new_AGEMA_signal_6057) );
  DFF_X1 new_AGEMA_reg_buffer_4173_s_current_state_reg ( .D(
        new_AGEMA_signal_6060), .CK(clk), .Q(new_AGEMA_signal_6061) );
  DFF_X1 new_AGEMA_reg_buffer_4177_s_current_state_reg ( .D(
        new_AGEMA_signal_6064), .CK(clk), .Q(new_AGEMA_signal_6065) );
  DFF_X1 new_AGEMA_reg_buffer_4181_s_current_state_reg ( .D(
        new_AGEMA_signal_6068), .CK(clk), .Q(new_AGEMA_signal_6069) );
  DFF_X1 new_AGEMA_reg_buffer_4185_s_current_state_reg ( .D(
        new_AGEMA_signal_6072), .CK(clk), .Q(new_AGEMA_signal_6073) );
  DFF_X1 new_AGEMA_reg_buffer_4189_s_current_state_reg ( .D(
        new_AGEMA_signal_6076), .CK(clk), .Q(new_AGEMA_signal_6077) );
  DFF_X1 new_AGEMA_reg_buffer_4193_s_current_state_reg ( .D(
        new_AGEMA_signal_6080), .CK(clk), .Q(new_AGEMA_signal_6081) );
  DFF_X1 new_AGEMA_reg_buffer_4197_s_current_state_reg ( .D(
        new_AGEMA_signal_6084), .CK(clk), .Q(new_AGEMA_signal_6085) );
  DFF_X1 new_AGEMA_reg_buffer_4201_s_current_state_reg ( .D(
        new_AGEMA_signal_6088), .CK(clk), .Q(new_AGEMA_signal_6089) );
  DFF_X1 new_AGEMA_reg_buffer_4205_s_current_state_reg ( .D(
        new_AGEMA_signal_6092), .CK(clk), .Q(new_AGEMA_signal_6093) );
  DFF_X1 new_AGEMA_reg_buffer_4209_s_current_state_reg ( .D(
        new_AGEMA_signal_6096), .CK(clk), .Q(new_AGEMA_signal_6097) );
  DFF_X1 new_AGEMA_reg_buffer_4213_s_current_state_reg ( .D(
        new_AGEMA_signal_6100), .CK(clk), .Q(new_AGEMA_signal_6101) );
  DFF_X1 new_AGEMA_reg_buffer_4217_s_current_state_reg ( .D(
        new_AGEMA_signal_6104), .CK(clk), .Q(new_AGEMA_signal_6105) );
  DFF_X1 new_AGEMA_reg_buffer_4221_s_current_state_reg ( .D(
        new_AGEMA_signal_6108), .CK(clk), .Q(new_AGEMA_signal_6109) );
  DFF_X1 new_AGEMA_reg_buffer_4225_s_current_state_reg ( .D(
        new_AGEMA_signal_6112), .CK(clk), .Q(new_AGEMA_signal_6113) );
  DFF_X1 new_AGEMA_reg_buffer_4229_s_current_state_reg ( .D(
        new_AGEMA_signal_6116), .CK(clk), .Q(new_AGEMA_signal_6117) );
  DFF_X1 new_AGEMA_reg_buffer_4233_s_current_state_reg ( .D(
        new_AGEMA_signal_6120), .CK(clk), .Q(new_AGEMA_signal_6121) );
  DFF_X1 new_AGEMA_reg_buffer_4237_s_current_state_reg ( .D(
        new_AGEMA_signal_6124), .CK(clk), .Q(new_AGEMA_signal_6125) );
  DFF_X1 new_AGEMA_reg_buffer_4241_s_current_state_reg ( .D(
        new_AGEMA_signal_6128), .CK(clk), .Q(new_AGEMA_signal_6129) );
  DFF_X1 new_AGEMA_reg_buffer_4245_s_current_state_reg ( .D(
        new_AGEMA_signal_6132), .CK(clk), .Q(new_AGEMA_signal_6133) );
  DFF_X1 new_AGEMA_reg_buffer_4249_s_current_state_reg ( .D(
        new_AGEMA_signal_6136), .CK(clk), .Q(new_AGEMA_signal_6137) );
  DFF_X1 new_AGEMA_reg_buffer_4253_s_current_state_reg ( .D(
        new_AGEMA_signal_6140), .CK(clk), .Q(new_AGEMA_signal_6141) );
  DFF_X1 new_AGEMA_reg_buffer_4257_s_current_state_reg ( .D(
        new_AGEMA_signal_6144), .CK(clk), .Q(new_AGEMA_signal_6145) );
  DFF_X1 new_AGEMA_reg_buffer_4261_s_current_state_reg ( .D(
        new_AGEMA_signal_6148), .CK(clk), .Q(new_AGEMA_signal_6149) );
  DFF_X1 new_AGEMA_reg_buffer_4265_s_current_state_reg ( .D(
        new_AGEMA_signal_6152), .CK(clk), .Q(new_AGEMA_signal_6153) );
  DFF_X1 new_AGEMA_reg_buffer_4269_s_current_state_reg ( .D(
        new_AGEMA_signal_6156), .CK(clk), .Q(new_AGEMA_signal_6157) );
  DFF_X1 new_AGEMA_reg_buffer_4273_s_current_state_reg ( .D(
        new_AGEMA_signal_6160), .CK(clk), .Q(new_AGEMA_signal_6161) );
  DFF_X1 new_AGEMA_reg_buffer_4277_s_current_state_reg ( .D(
        new_AGEMA_signal_6164), .CK(clk), .Q(new_AGEMA_signal_6165) );
  DFF_X1 new_AGEMA_reg_buffer_4281_s_current_state_reg ( .D(
        new_AGEMA_signal_6168), .CK(clk), .Q(new_AGEMA_signal_6169) );
  DFF_X1 new_AGEMA_reg_buffer_4285_s_current_state_reg ( .D(
        new_AGEMA_signal_6172), .CK(clk), .Q(new_AGEMA_signal_6173) );
  DFF_X1 new_AGEMA_reg_buffer_4289_s_current_state_reg ( .D(
        new_AGEMA_signal_6176), .CK(clk), .Q(new_AGEMA_signal_6177) );
  DFF_X1 new_AGEMA_reg_buffer_4293_s_current_state_reg ( .D(
        new_AGEMA_signal_6180), .CK(clk), .Q(new_AGEMA_signal_6181) );
  DFF_X1 new_AGEMA_reg_buffer_4297_s_current_state_reg ( .D(
        new_AGEMA_signal_6184), .CK(clk), .Q(new_AGEMA_signal_6185) );
  DFF_X1 new_AGEMA_reg_buffer_4301_s_current_state_reg ( .D(
        new_AGEMA_signal_6188), .CK(clk), .Q(new_AGEMA_signal_6189) );
  DFF_X1 new_AGEMA_reg_buffer_4305_s_current_state_reg ( .D(
        new_AGEMA_signal_6192), .CK(clk), .Q(new_AGEMA_signal_6193) );
  DFF_X1 new_AGEMA_reg_buffer_4309_s_current_state_reg ( .D(
        new_AGEMA_signal_6196), .CK(clk), .Q(new_AGEMA_signal_6197) );
  DFF_X1 new_AGEMA_reg_buffer_4313_s_current_state_reg ( .D(
        new_AGEMA_signal_6200), .CK(clk), .Q(new_AGEMA_signal_6201) );
  DFF_X1 new_AGEMA_reg_buffer_4317_s_current_state_reg ( .D(
        new_AGEMA_signal_6204), .CK(clk), .Q(new_AGEMA_signal_6205) );
  DFF_X1 new_AGEMA_reg_buffer_4321_s_current_state_reg ( .D(
        new_AGEMA_signal_6208), .CK(clk), .Q(new_AGEMA_signal_6209) );
  DFF_X1 new_AGEMA_reg_buffer_4325_s_current_state_reg ( .D(
        new_AGEMA_signal_6212), .CK(clk), .Q(new_AGEMA_signal_6213) );
  DFF_X1 new_AGEMA_reg_buffer_4329_s_current_state_reg ( .D(
        new_AGEMA_signal_6216), .CK(clk), .Q(new_AGEMA_signal_6217) );
  DFF_X1 new_AGEMA_reg_buffer_4333_s_current_state_reg ( .D(
        new_AGEMA_signal_6220), .CK(clk), .Q(new_AGEMA_signal_6221) );
  DFF_X1 new_AGEMA_reg_buffer_4337_s_current_state_reg ( .D(
        new_AGEMA_signal_6224), .CK(clk), .Q(new_AGEMA_signal_6225) );
  DFF_X1 new_AGEMA_reg_buffer_4341_s_current_state_reg ( .D(
        new_AGEMA_signal_6228), .CK(clk), .Q(new_AGEMA_signal_6229) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4277), .CK(clk), .Q(ciphertext_s0[120]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4281), .CK(clk), .Q(ciphertext_s1[120]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4285), .CK(clk), .Q(ciphertext_s0[121]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4289), .CK(clk), .Q(ciphertext_s1[121]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4293), .CK(clk), .Q(ciphertext_s0[122]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4297), .CK(clk), .Q(ciphertext_s1[122]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4301), .CK(clk), .Q(ciphertext_s0[123]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4305), .CK(clk), .Q(ciphertext_s1[123]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4309), .CK(clk), .Q(ciphertext_s0[124]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4313), .CK(clk), .Q(ciphertext_s1[124]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4317), .CK(clk), .Q(ciphertext_s0[125]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4321), .CK(clk), .Q(ciphertext_s1[125]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4325), .CK(clk), .Q(ciphertext_s0[126]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4329), .CK(clk), .Q(ciphertext_s1[126]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4333), .CK(clk), .Q(ciphertext_s0[127]) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4337), .CK(clk), .Q(ciphertext_s1[127]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4341), .CK(clk), .Q(ciphertext_s0[112]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4345), .CK(clk), .Q(ciphertext_s1[112]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4349), .CK(clk), .Q(ciphertext_s0[113]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4353), .CK(clk), .Q(ciphertext_s1[113]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4357), .CK(clk), .Q(ciphertext_s0[114]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4361), .CK(clk), .Q(ciphertext_s1[114]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4365), .CK(clk), .Q(ciphertext_s0[115]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4369), .CK(clk), .Q(ciphertext_s1[115]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4373), .CK(clk), .Q(ciphertext_s0[116]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4377), .CK(clk), .Q(ciphertext_s1[116]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4381), .CK(clk), .Q(ciphertext_s0[117]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4385), .CK(clk), .Q(ciphertext_s1[117]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4389), .CK(clk), .Q(ciphertext_s0[118]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4393), .CK(clk), .Q(ciphertext_s1[118]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4397), .CK(clk), .Q(ciphertext_s0[119]) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4401), .CK(clk), .Q(ciphertext_s1[119]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4405), .CK(clk), .Q(ciphertext_s0[104]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4409), .CK(clk), .Q(ciphertext_s1[104]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4413), .CK(clk), .Q(ciphertext_s0[105]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4417), .CK(clk), .Q(ciphertext_s1[105]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4421), .CK(clk), .Q(ciphertext_s0[106]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4425), .CK(clk), .Q(ciphertext_s1[106]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4429), .CK(clk), .Q(ciphertext_s0[107]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4433), .CK(clk), .Q(ciphertext_s1[107]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4437), .CK(clk), .Q(ciphertext_s0[108]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4441), .CK(clk), .Q(ciphertext_s1[108]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4445), .CK(clk), .Q(ciphertext_s0[109]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4449), .CK(clk), .Q(ciphertext_s1[109]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4453), .CK(clk), .Q(ciphertext_s0[110]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4457), .CK(clk), .Q(ciphertext_s1[110]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4461), .CK(clk), .Q(ciphertext_s0[111]) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4465), .CK(clk), .Q(ciphertext_s1[111]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4469), .CK(clk), .Q(ciphertext_s0[96]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4473), .CK(clk), .Q(ciphertext_s1[96]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4477), .CK(clk), .Q(ciphertext_s0[97]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4481), .CK(clk), .Q(ciphertext_s1[97]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4485), .CK(clk), .Q(ciphertext_s0[98]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4489), .CK(clk), .Q(ciphertext_s1[98]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4493), .CK(clk), .Q(ciphertext_s0[99]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4497), .CK(clk), .Q(ciphertext_s1[99]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4501), .CK(clk), .Q(ciphertext_s0[100]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4505), .CK(clk), .Q(ciphertext_s1[100]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4509), .CK(clk), .Q(ciphertext_s0[101]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4513), .CK(clk), .Q(ciphertext_s1[101]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4517), .CK(clk), .Q(ciphertext_s0[102]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4521), .CK(clk), .Q(ciphertext_s1[102]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4525), .CK(clk), .Q(ciphertext_s0[103]) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4529), .CK(clk), .Q(ciphertext_s1[103]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4533), .CK(clk), .Q(ciphertext_s0[88]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4537), .CK(clk), .Q(ciphertext_s1[88]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4541), .CK(clk), .Q(ciphertext_s0[89]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4545), .CK(clk), .Q(ciphertext_s1[89]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4549), .CK(clk), .Q(ciphertext_s0[90]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4553), .CK(clk), .Q(ciphertext_s1[90]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4557), .CK(clk), .Q(ciphertext_s0[91]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4561), .CK(clk), .Q(ciphertext_s1[91]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4565), .CK(clk), .Q(ciphertext_s0[92]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4569), .CK(clk), .Q(ciphertext_s1[92]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4573), .CK(clk), .Q(ciphertext_s0[93]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4577), .CK(clk), .Q(ciphertext_s1[93]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4581), .CK(clk), .Q(ciphertext_s0[94]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4585), .CK(clk), .Q(ciphertext_s1[94]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4589), .CK(clk), .Q(ciphertext_s0[95]) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4593), .CK(clk), .Q(ciphertext_s1[95]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4597), .CK(clk), .Q(ciphertext_s0[80]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4601), .CK(clk), .Q(ciphertext_s1[80]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4605), .CK(clk), .Q(ciphertext_s0[81]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4609), .CK(clk), .Q(ciphertext_s1[81]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4613), .CK(clk), .Q(ciphertext_s0[82]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4617), .CK(clk), .Q(ciphertext_s1[82]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4621), .CK(clk), .Q(ciphertext_s0[83]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4625), .CK(clk), .Q(ciphertext_s1[83]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4629), .CK(clk), .Q(ciphertext_s0[84]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4633), .CK(clk), .Q(ciphertext_s1[84]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4637), .CK(clk), .Q(ciphertext_s0[85]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4641), .CK(clk), .Q(ciphertext_s1[85]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4645), .CK(clk), .Q(ciphertext_s0[86]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4649), .CK(clk), .Q(ciphertext_s1[86]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4653), .CK(clk), .Q(ciphertext_s0[87]) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4657), .CK(clk), .Q(ciphertext_s1[87]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4661), .CK(clk), .Q(ciphertext_s0[72]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4665), .CK(clk), .Q(ciphertext_s1[72]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4669), .CK(clk), .Q(ciphertext_s0[73]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4673), .CK(clk), .Q(ciphertext_s1[73]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4677), .CK(clk), .Q(ciphertext_s0[74]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4681), .CK(clk), .Q(ciphertext_s1[74]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4685), .CK(clk), .Q(ciphertext_s0[75]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4689), .CK(clk), .Q(ciphertext_s1[75]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4693), .CK(clk), .Q(ciphertext_s0[76]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4697), .CK(clk), .Q(ciphertext_s1[76]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4701), .CK(clk), .Q(ciphertext_s0[77]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4705), .CK(clk), .Q(ciphertext_s1[77]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4709), .CK(clk), .Q(ciphertext_s0[78]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4713), .CK(clk), .Q(ciphertext_s1[78]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4717), .CK(clk), .Q(ciphertext_s0[79]) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4721), .CK(clk), .Q(ciphertext_s1[79]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4725), .CK(clk), .Q(ciphertext_s0[64]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4729), .CK(clk), .Q(ciphertext_s1[64]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4733), .CK(clk), .Q(ciphertext_s0[65]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4737), .CK(clk), .Q(ciphertext_s1[65]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4741), .CK(clk), .Q(ciphertext_s0[66]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4745), .CK(clk), .Q(ciphertext_s1[66]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4749), .CK(clk), .Q(ciphertext_s0[67]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4753), .CK(clk), .Q(ciphertext_s1[67]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4757), .CK(clk), .Q(ciphertext_s0[68]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4761), .CK(clk), .Q(ciphertext_s1[68]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4765), .CK(clk), .Q(ciphertext_s0[69]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4769), .CK(clk), .Q(ciphertext_s1[69]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4773), .CK(clk), .Q(ciphertext_s0[70]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4777), .CK(clk), .Q(ciphertext_s1[70]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4781), .CK(clk), .Q(ciphertext_s0[71]) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4785), .CK(clk), .Q(ciphertext_s1[71]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4789), .CK(clk), .Q(ciphertext_s0[56]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4793), .CK(clk), .Q(ciphertext_s1[56]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4797), .CK(clk), .Q(ciphertext_s0[57]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4801), .CK(clk), .Q(ciphertext_s1[57]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4805), .CK(clk), .Q(ciphertext_s0[58]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4809), .CK(clk), .Q(ciphertext_s1[58]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4813), .CK(clk), .Q(ciphertext_s0[59]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4817), .CK(clk), .Q(ciphertext_s1[59]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4821), .CK(clk), .Q(ciphertext_s0[60]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4825), .CK(clk), .Q(ciphertext_s1[60]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4829), .CK(clk), .Q(ciphertext_s0[61]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4833), .CK(clk), .Q(ciphertext_s1[61]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4837), .CK(clk), .Q(ciphertext_s0[62]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4841), .CK(clk), .Q(ciphertext_s1[62]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4845), .CK(clk), .Q(ciphertext_s0[63]) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4849), .CK(clk), .Q(ciphertext_s1[63]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4853), .CK(clk), .Q(ciphertext_s0[48]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4857), .CK(clk), .Q(ciphertext_s1[48]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4861), .CK(clk), .Q(ciphertext_s0[49]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4865), .CK(clk), .Q(ciphertext_s1[49]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4869), .CK(clk), .Q(ciphertext_s0[50]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4873), .CK(clk), .Q(ciphertext_s1[50]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4877), .CK(clk), .Q(ciphertext_s0[51]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4881), .CK(clk), .Q(ciphertext_s1[51]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4885), .CK(clk), .Q(ciphertext_s0[52]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4889), .CK(clk), .Q(ciphertext_s1[52]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4893), .CK(clk), .Q(ciphertext_s0[53]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4897), .CK(clk), .Q(ciphertext_s1[53]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4901), .CK(clk), .Q(ciphertext_s0[54]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4905), .CK(clk), .Q(ciphertext_s1[54]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4909), .CK(clk), .Q(ciphertext_s0[55]) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4913), .CK(clk), .Q(ciphertext_s1[55]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4917), .CK(clk), .Q(ciphertext_s0[40]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4921), .CK(clk), .Q(ciphertext_s1[40]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4925), .CK(clk), .Q(ciphertext_s0[41]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4929), .CK(clk), .Q(ciphertext_s1[41]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4933), .CK(clk), .Q(ciphertext_s0[42]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4937), .CK(clk), .Q(ciphertext_s1[42]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4941), .CK(clk), .Q(ciphertext_s0[43]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4945), .CK(clk), .Q(ciphertext_s1[43]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4949), .CK(clk), .Q(ciphertext_s0[44]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4953), .CK(clk), .Q(ciphertext_s1[44]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4957), .CK(clk), .Q(ciphertext_s0[45]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4961), .CK(clk), .Q(ciphertext_s1[45]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4965), .CK(clk), .Q(ciphertext_s0[46]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4969), .CK(clk), .Q(ciphertext_s1[46]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4973), .CK(clk), .Q(ciphertext_s0[47]) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4977), .CK(clk), .Q(ciphertext_s1[47]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4981), .CK(clk), .Q(ciphertext_s0[32]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4985), .CK(clk), .Q(ciphertext_s1[32]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4989), .CK(clk), .Q(ciphertext_s0[33]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_4993), .CK(clk), .Q(ciphertext_s1[33]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_4997), .CK(clk), .Q(ciphertext_s0[34]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5001), .CK(clk), .Q(ciphertext_s1[34]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5005), .CK(clk), .Q(ciphertext_s0[35]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5009), .CK(clk), .Q(ciphertext_s1[35]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5013), .CK(clk), .Q(ciphertext_s0[36]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5017), .CK(clk), .Q(ciphertext_s1[36]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5021), .CK(clk), .Q(ciphertext_s0[37]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5025), .CK(clk), .Q(ciphertext_s1[37]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5029), .CK(clk), .Q(ciphertext_s0[38]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5033), .CK(clk), .Q(ciphertext_s1[38]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5037), .CK(clk), .Q(ciphertext_s0[39]) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5041), .CK(clk), .Q(ciphertext_s1[39]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5045), .CK(clk), .Q(ciphertext_s0[24]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5049), .CK(clk), .Q(ciphertext_s1[24]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5053), .CK(clk), .Q(ciphertext_s0[25]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5057), .CK(clk), .Q(ciphertext_s1[25]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5061), .CK(clk), .Q(ciphertext_s0[26]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5065), .CK(clk), .Q(ciphertext_s1[26]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5069), .CK(clk), .Q(ciphertext_s0[27]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5073), .CK(clk), .Q(ciphertext_s1[27]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5077), .CK(clk), .Q(ciphertext_s0[28]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5081), .CK(clk), .Q(ciphertext_s1[28]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5085), .CK(clk), .Q(ciphertext_s0[29]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5089), .CK(clk), .Q(ciphertext_s1[29]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5093), .CK(clk), .Q(ciphertext_s0[30]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5097), .CK(clk), .Q(ciphertext_s1[30]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5101), .CK(clk), .Q(ciphertext_s0[31]) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5105), .CK(clk), .Q(ciphertext_s1[31]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5109), .CK(clk), .Q(ciphertext_s0[16]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5113), .CK(clk), .Q(ciphertext_s1[16]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5117), .CK(clk), .Q(ciphertext_s0[17]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5121), .CK(clk), .Q(ciphertext_s1[17]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5125), .CK(clk), .Q(ciphertext_s0[18]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5129), .CK(clk), .Q(ciphertext_s1[18]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5133), .CK(clk), .Q(ciphertext_s0[19]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5137), .CK(clk), .Q(ciphertext_s1[19]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5141), .CK(clk), .Q(ciphertext_s0[20]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5145), .CK(clk), .Q(ciphertext_s1[20]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5149), .CK(clk), .Q(ciphertext_s0[21]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5153), .CK(clk), .Q(ciphertext_s1[21]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5157), .CK(clk), .Q(ciphertext_s0[22]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5161), .CK(clk), .Q(ciphertext_s1[22]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5165), .CK(clk), .Q(ciphertext_s0[23]) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5169), .CK(clk), .Q(ciphertext_s1[23]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5173), .CK(clk), .Q(ciphertext_s0[8]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5177), .CK(clk), .Q(ciphertext_s1[8]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5181), .CK(clk), .Q(ciphertext_s0[9]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5185), .CK(clk), .Q(ciphertext_s1[9]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5189), .CK(clk), .Q(ciphertext_s0[10]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5193), .CK(clk), .Q(ciphertext_s1[10]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5197), .CK(clk), .Q(ciphertext_s0[11]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5201), .CK(clk), .Q(ciphertext_s1[11]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5205), .CK(clk), .Q(ciphertext_s0[12]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5209), .CK(clk), .Q(ciphertext_s1[12]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5213), .CK(clk), .Q(ciphertext_s0[13]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5217), .CK(clk), .Q(ciphertext_s1[13]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5221), .CK(clk), .Q(ciphertext_s0[14]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5225), .CK(clk), .Q(ciphertext_s1[14]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5229), .CK(clk), .Q(ciphertext_s0[15]) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5233), .CK(clk), .Q(ciphertext_s1[15]) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(stateArray_S33reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext_s0[0])
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3497), .CK(clk), .Q(ciphertext_s1[0]) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(stateArray_S33reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext_s0[1])
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3520), .CK(clk), .Q(ciphertext_s1[1]) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(stateArray_S33reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext_s0[2])
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3521), .CK(clk), .Q(ciphertext_s1[2]) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(stateArray_S33reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext_s0[3])
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3522), .CK(clk), .Q(ciphertext_s1[3]) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(stateArray_S33reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext_s0[4])
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3523), .CK(clk), .Q(ciphertext_s1[4]) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(stateArray_S33reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext_s0[5])
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3524), .CK(clk), .Q(ciphertext_s1[5]) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(stateArray_S33reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext_s0[6])
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3525), .CK(clk), .Q(ciphertext_s1[6]) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(stateArray_S33reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext_s0[7])
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3526), .CK(clk), .Q(ciphertext_s1[7]) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5237), .CK(clk), .Q(keyStateIn[0]) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5241), .CK(clk), .Q(new_AGEMA_signal_1983) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5245), .CK(clk), .Q(keyStateIn[1]) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5249), .CK(clk), .Q(new_AGEMA_signal_1986) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5253), .CK(clk), .Q(keyStateIn[2]) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5257), .CK(clk), .Q(new_AGEMA_signal_1989) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5261), .CK(clk), .Q(keyStateIn[3]) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5265), .CK(clk), .Q(new_AGEMA_signal_1992) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5269), .CK(clk), .Q(keyStateIn[4]) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5273), .CK(clk), .Q(new_AGEMA_signal_1995) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5277), .CK(clk), .Q(keyStateIn[5]) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5281), .CK(clk), .Q(new_AGEMA_signal_1998) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5285), .CK(clk), .Q(keyStateIn[6]) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5289), .CK(clk), .Q(new_AGEMA_signal_2001) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5293), .CK(clk), .Q(keyStateIn[7]) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5297), .CK(clk), .Q(new_AGEMA_signal_2004) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5301), .CK(clk), .Q(KeyArray_outS01ser_0_) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5305), .CK(clk), .Q(new_AGEMA_signal_2020) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5309), .CK(clk), .Q(KeyArray_outS01ser_1_) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5313), .CK(clk), .Q(new_AGEMA_signal_2018) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5317), .CK(clk), .Q(KeyArray_outS01ser_2_) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5321), .CK(clk), .Q(new_AGEMA_signal_2016) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5325), .CK(clk), .Q(KeyArray_outS01ser_3_) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5329), .CK(clk), .Q(new_AGEMA_signal_2014) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5333), .CK(clk), .Q(KeyArray_outS01ser_4_) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5337), .CK(clk), .Q(new_AGEMA_signal_2012) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5341), .CK(clk), .Q(KeyArray_outS01ser_5_) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5345), .CK(clk), .Q(new_AGEMA_signal_2010) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5349), .CK(clk), .Q(KeyArray_outS01ser_6_) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5353), .CK(clk), .Q(new_AGEMA_signal_2008) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5357), .CK(clk), .Q(KeyArray_outS01ser_7_) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5361), .CK(clk), .Q(new_AGEMA_signal_2006) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5365), .CK(clk), .Q(KeyArray_outS02ser[0]) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5369), .CK(clk), .Q(new_AGEMA_signal_2443) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5373), .CK(clk), .Q(KeyArray_outS02ser[1]) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5377), .CK(clk), .Q(new_AGEMA_signal_2446) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5381), .CK(clk), .Q(KeyArray_outS02ser[2]) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5385), .CK(clk), .Q(new_AGEMA_signal_2449) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5389), .CK(clk), .Q(KeyArray_outS02ser[3]) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5393), .CK(clk), .Q(new_AGEMA_signal_2452) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5397), .CK(clk), .Q(KeyArray_outS02ser[4]) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5401), .CK(clk), .Q(new_AGEMA_signal_2455) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5405), .CK(clk), .Q(KeyArray_outS02ser[5]) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5409), .CK(clk), .Q(new_AGEMA_signal_2458) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5413), .CK(clk), .Q(KeyArray_outS02ser[6]) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5417), .CK(clk), .Q(new_AGEMA_signal_2461) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5421), .CK(clk), .Q(KeyArray_outS02ser[7]) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5425), .CK(clk), .Q(new_AGEMA_signal_2464) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5429), .CK(clk), .Q(KeyArray_outS03ser[0]) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5433), .CK(clk), .Q(new_AGEMA_signal_2467) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5437), .CK(clk), .Q(KeyArray_outS03ser[1]) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5441), .CK(clk), .Q(new_AGEMA_signal_2470) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5445), .CK(clk), .Q(KeyArray_outS03ser[2]) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5449), .CK(clk), .Q(new_AGEMA_signal_2473) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5453), .CK(clk), .Q(KeyArray_outS03ser[3]) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5457), .CK(clk), .Q(new_AGEMA_signal_2476) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5461), .CK(clk), .Q(KeyArray_outS03ser[4]) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5465), .CK(clk), .Q(new_AGEMA_signal_2479) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5469), .CK(clk), .Q(KeyArray_outS03ser[5]) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5473), .CK(clk), .Q(new_AGEMA_signal_2482) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5477), .CK(clk), .Q(KeyArray_outS03ser[6]) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5481), .CK(clk), .Q(new_AGEMA_signal_2485) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5485), .CK(clk), .Q(KeyArray_outS03ser[7]) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5489), .CK(clk), .Q(new_AGEMA_signal_2488) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5493), .CK(clk), .Q(KeyArray_outS10ser[0]) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5497), .CK(clk), .Q(new_AGEMA_signal_2491) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5501), .CK(clk), .Q(KeyArray_outS10ser[1]) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5505), .CK(clk), .Q(new_AGEMA_signal_2494) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5509), .CK(clk), .Q(KeyArray_outS10ser[2]) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5513), .CK(clk), .Q(new_AGEMA_signal_2497) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5517), .CK(clk), .Q(KeyArray_outS10ser[3]) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5521), .CK(clk), .Q(new_AGEMA_signal_2500) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5525), .CK(clk), .Q(KeyArray_outS10ser[4]) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5529), .CK(clk), .Q(new_AGEMA_signal_2503) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5533), .CK(clk), .Q(KeyArray_outS10ser[5]) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5537), .CK(clk), .Q(new_AGEMA_signal_2506) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5541), .CK(clk), .Q(KeyArray_outS10ser[6]) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5545), .CK(clk), .Q(new_AGEMA_signal_2509) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5549), .CK(clk), .Q(KeyArray_outS10ser[7]) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5553), .CK(clk), .Q(new_AGEMA_signal_2512) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5557), .CK(clk), .Q(KeyArray_outS11ser[0]) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5561), .CK(clk), .Q(new_AGEMA_signal_2515) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5565), .CK(clk), .Q(KeyArray_outS11ser[1]) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5569), .CK(clk), .Q(new_AGEMA_signal_2518) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5573), .CK(clk), .Q(KeyArray_outS11ser[2]) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5577), .CK(clk), .Q(new_AGEMA_signal_2521) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5581), .CK(clk), .Q(KeyArray_outS11ser[3]) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5585), .CK(clk), .Q(new_AGEMA_signal_2524) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5589), .CK(clk), .Q(KeyArray_outS11ser[4]) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5593), .CK(clk), .Q(new_AGEMA_signal_2527) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5597), .CK(clk), .Q(KeyArray_outS11ser[5]) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5601), .CK(clk), .Q(new_AGEMA_signal_2530) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5605), .CK(clk), .Q(KeyArray_outS11ser[6]) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5609), .CK(clk), .Q(new_AGEMA_signal_2533) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5613), .CK(clk), .Q(KeyArray_outS11ser[7]) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5617), .CK(clk), .Q(new_AGEMA_signal_2536) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5621), .CK(clk), .Q(KeyArray_outS12ser[0]) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5625), .CK(clk), .Q(new_AGEMA_signal_2539) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5629), .CK(clk), .Q(KeyArray_outS12ser[1]) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5633), .CK(clk), .Q(new_AGEMA_signal_2542) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5637), .CK(clk), .Q(KeyArray_outS12ser[2]) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5641), .CK(clk), .Q(new_AGEMA_signal_2545) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5645), .CK(clk), .Q(KeyArray_outS12ser[3]) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5649), .CK(clk), .Q(new_AGEMA_signal_2548) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5653), .CK(clk), .Q(KeyArray_outS12ser[4]) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5657), .CK(clk), .Q(new_AGEMA_signal_2551) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5661), .CK(clk), .Q(KeyArray_outS12ser[5]) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5665), .CK(clk), .Q(new_AGEMA_signal_2554) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5669), .CK(clk), .Q(KeyArray_outS12ser[6]) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5673), .CK(clk), .Q(new_AGEMA_signal_2557) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5677), .CK(clk), .Q(KeyArray_outS12ser[7]) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5681), .CK(clk), .Q(new_AGEMA_signal_2560) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5685), .CK(clk), .Q(keySBIn[0]) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5689), .CK(clk), .Q(new_AGEMA_signal_2563) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5693), .CK(clk), .Q(keySBIn[1]) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5697), .CK(clk), .Q(new_AGEMA_signal_2566) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5701), .CK(clk), .Q(keySBIn[2]) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5705), .CK(clk), .Q(new_AGEMA_signal_2569) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5709), .CK(clk), .Q(keySBIn[3]) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5713), .CK(clk), .Q(new_AGEMA_signal_2572) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5717), .CK(clk), .Q(keySBIn[4]) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5721), .CK(clk), .Q(new_AGEMA_signal_2575) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5725), .CK(clk), .Q(keySBIn[5]) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5729), .CK(clk), .Q(new_AGEMA_signal_2578) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5733), .CK(clk), .Q(keySBIn[6]) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5737), .CK(clk), .Q(new_AGEMA_signal_2581) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5741), .CK(clk), .Q(keySBIn[7]) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5745), .CK(clk), .Q(new_AGEMA_signal_2584) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5749), .CK(clk), .Q(KeyArray_outS20ser[0]) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5753), .CK(clk), .Q(new_AGEMA_signal_2587) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5757), .CK(clk), .Q(KeyArray_outS20ser[1]) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5761), .CK(clk), .Q(new_AGEMA_signal_2590) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5765), .CK(clk), .Q(KeyArray_outS20ser[2]) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5769), .CK(clk), .Q(new_AGEMA_signal_2593) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5773), .CK(clk), .Q(KeyArray_outS20ser[3]) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5777), .CK(clk), .Q(new_AGEMA_signal_2596) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5781), .CK(clk), .Q(KeyArray_outS20ser[4]) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5785), .CK(clk), .Q(new_AGEMA_signal_2599) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5789), .CK(clk), .Q(KeyArray_outS20ser[5]) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5793), .CK(clk), .Q(new_AGEMA_signal_2602) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5797), .CK(clk), .Q(KeyArray_outS20ser[6]) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5801), .CK(clk), .Q(new_AGEMA_signal_2605) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5805), .CK(clk), .Q(KeyArray_outS20ser[7]) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5809), .CK(clk), .Q(new_AGEMA_signal_2608) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5813), .CK(clk), .Q(KeyArray_outS21ser[0]) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5817), .CK(clk), .Q(new_AGEMA_signal_2611) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5821), .CK(clk), .Q(KeyArray_outS21ser[1]) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5825), .CK(clk), .Q(new_AGEMA_signal_2614) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5829), .CK(clk), .Q(KeyArray_outS21ser[2]) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5833), .CK(clk), .Q(new_AGEMA_signal_2617) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5837), .CK(clk), .Q(KeyArray_outS21ser[3]) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5841), .CK(clk), .Q(new_AGEMA_signal_2620) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5845), .CK(clk), .Q(KeyArray_outS21ser[4]) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5849), .CK(clk), .Q(new_AGEMA_signal_2623) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5853), .CK(clk), .Q(KeyArray_outS21ser[5]) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5857), .CK(clk), .Q(new_AGEMA_signal_2626) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5861), .CK(clk), .Q(KeyArray_outS21ser[6]) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5865), .CK(clk), .Q(new_AGEMA_signal_2629) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5869), .CK(clk), .Q(KeyArray_outS21ser[7]) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5873), .CK(clk), .Q(new_AGEMA_signal_2632) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5877), .CK(clk), .Q(KeyArray_outS22ser[0]) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5881), .CK(clk), .Q(new_AGEMA_signal_2635) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5885), .CK(clk), .Q(KeyArray_outS22ser[1]) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5889), .CK(clk), .Q(new_AGEMA_signal_2638) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5893), .CK(clk), .Q(KeyArray_outS22ser[2]) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5897), .CK(clk), .Q(new_AGEMA_signal_2641) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5901), .CK(clk), .Q(KeyArray_outS22ser[3]) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5905), .CK(clk), .Q(new_AGEMA_signal_2644) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5909), .CK(clk), .Q(KeyArray_outS22ser[4]) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5913), .CK(clk), .Q(new_AGEMA_signal_2647) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5917), .CK(clk), .Q(KeyArray_outS22ser[5]) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5921), .CK(clk), .Q(new_AGEMA_signal_2650) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5925), .CK(clk), .Q(KeyArray_outS22ser[6]) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5929), .CK(clk), .Q(new_AGEMA_signal_2653) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5933), .CK(clk), .Q(KeyArray_outS22ser[7]) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5937), .CK(clk), .Q(new_AGEMA_signal_2656) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5941), .CK(clk), .Q(KeyArray_outS23ser[0]) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5945), .CK(clk), .Q(new_AGEMA_signal_2659) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5949), .CK(clk), .Q(KeyArray_outS23ser[1]) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5953), .CK(clk), .Q(new_AGEMA_signal_2662) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5957), .CK(clk), .Q(KeyArray_outS23ser[2]) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5961), .CK(clk), .Q(new_AGEMA_signal_2665) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5965), .CK(clk), .Q(KeyArray_outS23ser[3]) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5969), .CK(clk), .Q(new_AGEMA_signal_2668) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5973), .CK(clk), .Q(KeyArray_outS23ser[4]) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5977), .CK(clk), .Q(new_AGEMA_signal_2671) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5981), .CK(clk), .Q(KeyArray_outS23ser[5]) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5985), .CK(clk), .Q(new_AGEMA_signal_2674) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5989), .CK(clk), .Q(KeyArray_outS23ser[6]) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_5993), .CK(clk), .Q(new_AGEMA_signal_2677) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_5997), .CK(clk), .Q(KeyArray_outS23ser[7]) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6001), .CK(clk), .Q(new_AGEMA_signal_2680) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(KeyArray_S30reg_gff_1_SFF_0_n5), .CK(clk), .Q(KeyArray_outS30ser[0]) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3512), .CK(clk), .Q(new_AGEMA_signal_2683) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(KeyArray_S30reg_gff_1_SFF_1_n5), .CK(clk), .Q(KeyArray_outS30ser[1]) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3527), .CK(clk), .Q(new_AGEMA_signal_2686) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(KeyArray_S30reg_gff_1_SFF_2_n5), .CK(clk), .Q(KeyArray_outS30ser[2]) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3528), .CK(clk), .Q(new_AGEMA_signal_2689) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(KeyArray_S30reg_gff_1_SFF_3_n5), .CK(clk), .Q(KeyArray_outS30ser[3]) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3529), .CK(clk), .Q(new_AGEMA_signal_2692) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(KeyArray_S30reg_gff_1_SFF_4_n5), .CK(clk), .Q(KeyArray_outS30ser[4]) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3530), .CK(clk), .Q(new_AGEMA_signal_2695) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(KeyArray_S30reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS30ser[5]) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3531), .CK(clk), .Q(new_AGEMA_signal_2698) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(KeyArray_S30reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS30ser[6]) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3532), .CK(clk), .Q(new_AGEMA_signal_2701) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(KeyArray_S30reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS30ser[7]) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_3533), .CK(clk), .Q(new_AGEMA_signal_2704) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6005), .CK(clk), .Q(KeyArray_outS31ser[0]) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6009), .CK(clk), .Q(new_AGEMA_signal_2707) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6013), .CK(clk), .Q(KeyArray_outS31ser[1]) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6017), .CK(clk), .Q(new_AGEMA_signal_2710) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6021), .CK(clk), .Q(KeyArray_outS31ser[2]) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6025), .CK(clk), .Q(new_AGEMA_signal_2713) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6029), .CK(clk), .Q(KeyArray_outS31ser[3]) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6033), .CK(clk), .Q(new_AGEMA_signal_2716) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6037), .CK(clk), .Q(KeyArray_outS31ser[4]) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6041), .CK(clk), .Q(new_AGEMA_signal_2719) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6045), .CK(clk), .Q(KeyArray_outS31ser[5]) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6049), .CK(clk), .Q(new_AGEMA_signal_2722) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6053), .CK(clk), .Q(KeyArray_outS31ser[6]) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6057), .CK(clk), .Q(new_AGEMA_signal_2725) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6061), .CK(clk), .Q(KeyArray_outS31ser[7]) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6065), .CK(clk), .Q(new_AGEMA_signal_2728) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6069), .CK(clk), .Q(KeyArray_outS32ser[0]) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6073), .CK(clk), .Q(new_AGEMA_signal_2731) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6077), .CK(clk), .Q(KeyArray_outS32ser[1]) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6081), .CK(clk), .Q(new_AGEMA_signal_2734) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6085), .CK(clk), .Q(KeyArray_outS32ser[2]) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6089), .CK(clk), .Q(new_AGEMA_signal_2737) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6093), .CK(clk), .Q(KeyArray_outS32ser[3]) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6097), .CK(clk), .Q(new_AGEMA_signal_2740) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6101), .CK(clk), .Q(KeyArray_outS32ser[4]) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6105), .CK(clk), .Q(new_AGEMA_signal_2743) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6109), .CK(clk), .Q(KeyArray_outS32ser[5]) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6113), .CK(clk), .Q(new_AGEMA_signal_2746) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6117), .CK(clk), .Q(KeyArray_outS32ser[6]) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6121), .CK(clk), .Q(new_AGEMA_signal_2749) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6125), .CK(clk), .Q(KeyArray_outS32ser[7]) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6129), .CK(clk), .Q(new_AGEMA_signal_2752) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6133), .CK(clk), .Q(KeyArray_outS33ser[0]) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6137), .CK(clk), .Q(new_AGEMA_signal_2755) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6141), .CK(clk), .Q(KeyArray_outS33ser[1]) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6145), .CK(clk), .Q(new_AGEMA_signal_2758) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6149), .CK(clk), .Q(KeyArray_outS33ser[2]) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6153), .CK(clk), .Q(new_AGEMA_signal_2761) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6157), .CK(clk), .Q(KeyArray_outS33ser[3]) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6161), .CK(clk), .Q(new_AGEMA_signal_2764) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6165), .CK(clk), .Q(KeyArray_outS33ser[4]) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6169), .CK(clk), .Q(new_AGEMA_signal_2767) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6173), .CK(clk), .Q(KeyArray_outS33ser[5]) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6177), .CK(clk), .Q(new_AGEMA_signal_2770) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6181), .CK(clk), .Q(KeyArray_outS33ser[6]) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6185), .CK(clk), .Q(new_AGEMA_signal_2773) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg (
        .D(new_AGEMA_signal_6189), .CK(clk), .Q(KeyArray_outS33ser[7]) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg (
        .D(new_AGEMA_signal_6193), .CK(clk), .Q(new_AGEMA_signal_2776) );
endmodule

