
module circuit ( ClkxCI, XxDI, Zmul1xDI, Zmul2xDI, Zmul3xDI, Zinv1xDI, 
        Zinv2xDI, Zinv3xDI, QxDO );
  input [23:0] XxDI;
  input [11:0] Zmul1xDI;
  input [11:0] Zmul2xDI;
  input [11:0] Zmul3xDI;
  input [5:0] Zinv1xDI;
  input [5:0] Zinv2xDI;
  input [5:0] Zinv3xDI;
  output [23:0] QxDO;
  input ClkxCI;
  wire   mappedxD_2__7_, mappedxD_2__6_, mappedxD_2__5_, mappedxD_2__4_,
         mappedxD_2__3_, mappedxD_2__1_, mappedxD_2__0_, mappedxD_1__7_,
         mappedxD_1__6_, mappedxD_1__5_, mappedxD_1__4_, mappedxD_1__3_,
         mappedxD_1__1_, mappedxD_1__0_, mappedxD_0__7_, mappedxD_0__6_,
         mappedxD_0__5_, mappedxD_0__4_, mappedxD_0__3_, mappedxD_0__1_,
         mappedxD_0__0_, InvMappedxD_0__6_, InvMappedxD_0__5_,
         InvMappedxD_0__1_, InvMappedxD_0__0_, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, input_mapping_2_n23, input_mapping_2_n22,
         input_mapping_2_n21, input_mapping_2_n20, input_mapping_2_n19,
         input_mapping_2_n18, input_mapping_2_n17, output_mapping_2_n9,
         output_mapping_2_n8, output_mapping_2_n7, input_mapping_1_n23,
         input_mapping_1_n22, input_mapping_1_n21, input_mapping_1_n20,
         input_mapping_1_n19, input_mapping_1_n18, input_mapping_1_n17,
         output_mapping_1_n9, output_mapping_1_n8, output_mapping_1_n7,
         input_mapping_0_n23, input_mapping_0_n22, input_mapping_0_n21,
         input_mapping_0_n20, input_mapping_0_n19, input_mapping_0_n18,
         input_mapping_0_n17, output_mapping_0_n9, output_mapping_0_n8,
         output_mapping_0_n7, mul_y0y1_n12, mul_y0y1_n11, mul_y0y1_n10,
         mul_y0y1_n9, mul_y0y1_n8, mul_y0y1_n7, mul_y0y1_n6, mul_y0y1_n5,
         mul_y0y1_n4, mul_y0y1_n3, mul_y0y1_n2, mul_y0y1_n1, mul_y0y1_n48,
         mul_y0y1_n47, mul_y0y1_n46, mul_y0y1_n45, mul_y0y1_n44, mul_y0y1_n43,
         mul_y0y1_n42, mul_y0y1_n41, mul_y0y1_n40, mul_y0y1_n39, mul_y0y1_n38,
         mul_y0y1_n37, mul_y0y1_n36, mul_y0y1_n35, mul_y0y1_n34, mul_y0y1_n33,
         mul_y0y1_n32, mul_y0y1_n31, mul_y0y1_n30, mul_y0y1_n29, mul_y0y1_n28,
         mul_y0y1_n27, mul_y0y1_n26, mul_y0y1_n25, mul_y0y1_n24, mul_y0y1_n23,
         mul_y0y1_n22, mul_y0y1_n21, mul_y0y1_n20, mul_y0y1_n19, mul_y0y1_n18,
         mul_y0y1_n17, mul_y0y1_n16, mul_y0y1_n15, mul_y0y1_n14, mul_y0y1_n13,
         mul_y0y1_Xi_mul_Yj_1__0_, mul_y0y1_Xi_mul_Yj_1__1_,
         mul_y0y1_Xi_mul_Yj_1__2_, mul_y0y1_Xi_mul_Yj_1__3_,
         mul_y0y1_Xi_mul_Yj_2__0_, mul_y0y1_Xi_mul_Yj_2__1_,
         mul_y0y1_Xi_mul_Yj_2__2_, mul_y0y1_Xi_mul_Yj_2__3_,
         mul_y0y1_Xi_mul_Yj_3__0_, mul_y0y1_Xi_mul_Yj_3__1_,
         mul_y0y1_Xi_mul_Yj_3__2_, mul_y0y1_Xi_mul_Yj_3__3_,
         mul_y0y1_Xi_mul_Yj_5__0_, mul_y0y1_Xi_mul_Yj_5__1_,
         mul_y0y1_Xi_mul_Yj_5__2_, mul_y0y1_Xi_mul_Yj_5__3_,
         mul_y0y1_Xi_mul_Yj_6__0_, mul_y0y1_Xi_mul_Yj_6__1_,
         mul_y0y1_Xi_mul_Yj_6__2_, mul_y0y1_Xi_mul_Yj_6__3_,
         mul_y0y1_Xi_mul_Yj_7__0_, mul_y0y1_Xi_mul_Yj_7__1_,
         mul_y0y1_Xi_mul_Yj_7__2_, mul_y0y1_Xi_mul_Yj_7__3_,
         mul_y0y1_gf4_mul_2_2_n77, mul_y0y1_gf4_mul_2_2_n76,
         mul_y0y1_gf4_mul_2_2_n75, mul_y0y1_gf4_mul_2_2_n74,
         mul_y0y1_gf4_mul_2_2_n73, mul_y0y1_gf4_mul_2_2_n72,
         mul_y0y1_gf4_mul_2_2_n71, mul_y0y1_gf4_mul_2_2_n70,
         mul_y0y1_gf4_mul_2_2_n69, mul_y0y1_gf4_mul_2_2_n68,
         mul_y0y1_gf4_mul_2_2_n67, mul_y0y1_gf4_mul_2_2_n66,
         mul_y0y1_gf4_mul_2_2_n65, mul_y0y1_gf4_mul_2_2_n64,
         mul_y0y1_gf4_mul_2_2_n63, mul_y0y1_gf4_mul_2_2_n62,
         mul_y0y1_gf4_mul_2_2_n61, mul_y0y1_gf4_mul_2_2_n60,
         mul_y0y1_gf4_mul_2_2_n59, mul_y0y1_gf4_mul_2_2_n58,
         mul_y0y1_gf4_mul_2_2_n57, mul_y0y1_gf4_mul_2_2_n56,
         mul_y0y1_gf4_mul_2_2_n55, mul_y0y1_gf4_mul_2_2_n54,
         mul_y0y1_gf4_mul_2_2_n53, mul_y0y1_gf4_mul_2_1_n77,
         mul_y0y1_gf4_mul_2_1_n76, mul_y0y1_gf4_mul_2_1_n75,
         mul_y0y1_gf4_mul_2_1_n74, mul_y0y1_gf4_mul_2_1_n73,
         mul_y0y1_gf4_mul_2_1_n72, mul_y0y1_gf4_mul_2_1_n71,
         mul_y0y1_gf4_mul_2_1_n70, mul_y0y1_gf4_mul_2_1_n69,
         mul_y0y1_gf4_mul_2_1_n68, mul_y0y1_gf4_mul_2_1_n67,
         mul_y0y1_gf4_mul_2_1_n66, mul_y0y1_gf4_mul_2_1_n65,
         mul_y0y1_gf4_mul_2_1_n64, mul_y0y1_gf4_mul_2_1_n63,
         mul_y0y1_gf4_mul_2_1_n62, mul_y0y1_gf4_mul_2_1_n61,
         mul_y0y1_gf4_mul_2_1_n60, mul_y0y1_gf4_mul_2_1_n59,
         mul_y0y1_gf4_mul_2_1_n58, mul_y0y1_gf4_mul_2_1_n57,
         mul_y0y1_gf4_mul_2_1_n56, mul_y0y1_gf4_mul_2_1_n55,
         mul_y0y1_gf4_mul_2_1_n54, mul_y0y1_gf4_mul_2_1_n53,
         mul_y0y1_gf4_mul_2_0_n77, mul_y0y1_gf4_mul_2_0_n76,
         mul_y0y1_gf4_mul_2_0_n75, mul_y0y1_gf4_mul_2_0_n74,
         mul_y0y1_gf4_mul_2_0_n73, mul_y0y1_gf4_mul_2_0_n72,
         mul_y0y1_gf4_mul_2_0_n71, mul_y0y1_gf4_mul_2_0_n70,
         mul_y0y1_gf4_mul_2_0_n69, mul_y0y1_gf4_mul_2_0_n68,
         mul_y0y1_gf4_mul_2_0_n67, mul_y0y1_gf4_mul_2_0_n66,
         mul_y0y1_gf4_mul_2_0_n65, mul_y0y1_gf4_mul_2_0_n64,
         mul_y0y1_gf4_mul_2_0_n63, mul_y0y1_gf4_mul_2_0_n62,
         mul_y0y1_gf4_mul_2_0_n61, mul_y0y1_gf4_mul_2_0_n60,
         mul_y0y1_gf4_mul_2_0_n59, mul_y0y1_gf4_mul_2_0_n58,
         mul_y0y1_gf4_mul_2_0_n57, mul_y0y1_gf4_mul_2_0_n56,
         mul_y0y1_gf4_mul_2_0_n55, mul_y0y1_gf4_mul_2_0_n54,
         mul_y0y1_gf4_mul_2_0_n53, mul_y0y1_gf4_mul_1_2_n77,
         mul_y0y1_gf4_mul_1_2_n76, mul_y0y1_gf4_mul_1_2_n75,
         mul_y0y1_gf4_mul_1_2_n74, mul_y0y1_gf4_mul_1_2_n73,
         mul_y0y1_gf4_mul_1_2_n72, mul_y0y1_gf4_mul_1_2_n71,
         mul_y0y1_gf4_mul_1_2_n70, mul_y0y1_gf4_mul_1_2_n69,
         mul_y0y1_gf4_mul_1_2_n68, mul_y0y1_gf4_mul_1_2_n67,
         mul_y0y1_gf4_mul_1_2_n66, mul_y0y1_gf4_mul_1_2_n65,
         mul_y0y1_gf4_mul_1_2_n64, mul_y0y1_gf4_mul_1_2_n63,
         mul_y0y1_gf4_mul_1_2_n62, mul_y0y1_gf4_mul_1_2_n61,
         mul_y0y1_gf4_mul_1_2_n60, mul_y0y1_gf4_mul_1_2_n59,
         mul_y0y1_gf4_mul_1_2_n58, mul_y0y1_gf4_mul_1_2_n57,
         mul_y0y1_gf4_mul_1_2_n56, mul_y0y1_gf4_mul_1_2_n55,
         mul_y0y1_gf4_mul_1_2_n54, mul_y0y1_gf4_mul_1_2_n53,
         mul_y0y1_gf4_mul_1_1_n77, mul_y0y1_gf4_mul_1_1_n76,
         mul_y0y1_gf4_mul_1_1_n75, mul_y0y1_gf4_mul_1_1_n74,
         mul_y0y1_gf4_mul_1_1_n73, mul_y0y1_gf4_mul_1_1_n72,
         mul_y0y1_gf4_mul_1_1_n71, mul_y0y1_gf4_mul_1_1_n70,
         mul_y0y1_gf4_mul_1_1_n69, mul_y0y1_gf4_mul_1_1_n68,
         mul_y0y1_gf4_mul_1_1_n67, mul_y0y1_gf4_mul_1_1_n66,
         mul_y0y1_gf4_mul_1_1_n65, mul_y0y1_gf4_mul_1_1_n64,
         mul_y0y1_gf4_mul_1_1_n63, mul_y0y1_gf4_mul_1_1_n62,
         mul_y0y1_gf4_mul_1_1_n61, mul_y0y1_gf4_mul_1_1_n60,
         mul_y0y1_gf4_mul_1_1_n59, mul_y0y1_gf4_mul_1_1_n58,
         mul_y0y1_gf4_mul_1_1_n57, mul_y0y1_gf4_mul_1_1_n56,
         mul_y0y1_gf4_mul_1_1_n55, mul_y0y1_gf4_mul_1_1_n54,
         mul_y0y1_gf4_mul_1_1_n53, mul_y0y1_gf4_mul_1_0_n77,
         mul_y0y1_gf4_mul_1_0_n76, mul_y0y1_gf4_mul_1_0_n75,
         mul_y0y1_gf4_mul_1_0_n74, mul_y0y1_gf4_mul_1_0_n73,
         mul_y0y1_gf4_mul_1_0_n72, mul_y0y1_gf4_mul_1_0_n71,
         mul_y0y1_gf4_mul_1_0_n70, mul_y0y1_gf4_mul_1_0_n69,
         mul_y0y1_gf4_mul_1_0_n68, mul_y0y1_gf4_mul_1_0_n67,
         mul_y0y1_gf4_mul_1_0_n66, mul_y0y1_gf4_mul_1_0_n65,
         mul_y0y1_gf4_mul_1_0_n64, mul_y0y1_gf4_mul_1_0_n63,
         mul_y0y1_gf4_mul_1_0_n62, mul_y0y1_gf4_mul_1_0_n61,
         mul_y0y1_gf4_mul_1_0_n60, mul_y0y1_gf4_mul_1_0_n59,
         mul_y0y1_gf4_mul_1_0_n58, mul_y0y1_gf4_mul_1_0_n57,
         mul_y0y1_gf4_mul_1_0_n56, mul_y0y1_gf4_mul_1_0_n55,
         mul_y0y1_gf4_mul_1_0_n54, mul_y0y1_gf4_mul_1_0_n53,
         mul_y0y1_gf4_mul_0_2_n77, mul_y0y1_gf4_mul_0_2_n76,
         mul_y0y1_gf4_mul_0_2_n75, mul_y0y1_gf4_mul_0_2_n74,
         mul_y0y1_gf4_mul_0_2_n73, mul_y0y1_gf4_mul_0_2_n72,
         mul_y0y1_gf4_mul_0_2_n71, mul_y0y1_gf4_mul_0_2_n70,
         mul_y0y1_gf4_mul_0_2_n69, mul_y0y1_gf4_mul_0_2_n68,
         mul_y0y1_gf4_mul_0_2_n67, mul_y0y1_gf4_mul_0_2_n66,
         mul_y0y1_gf4_mul_0_2_n65, mul_y0y1_gf4_mul_0_2_n64,
         mul_y0y1_gf4_mul_0_2_n63, mul_y0y1_gf4_mul_0_2_n62,
         mul_y0y1_gf4_mul_0_2_n61, mul_y0y1_gf4_mul_0_2_n60,
         mul_y0y1_gf4_mul_0_2_n59, mul_y0y1_gf4_mul_0_2_n58,
         mul_y0y1_gf4_mul_0_2_n57, mul_y0y1_gf4_mul_0_2_n56,
         mul_y0y1_gf4_mul_0_2_n55, mul_y0y1_gf4_mul_0_2_n54,
         mul_y0y1_gf4_mul_0_2_n53, mul_y0y1_gf4_mul_0_1_n77,
         mul_y0y1_gf4_mul_0_1_n76, mul_y0y1_gf4_mul_0_1_n75,
         mul_y0y1_gf4_mul_0_1_n74, mul_y0y1_gf4_mul_0_1_n73,
         mul_y0y1_gf4_mul_0_1_n72, mul_y0y1_gf4_mul_0_1_n71,
         mul_y0y1_gf4_mul_0_1_n70, mul_y0y1_gf4_mul_0_1_n69,
         mul_y0y1_gf4_mul_0_1_n68, mul_y0y1_gf4_mul_0_1_n67,
         mul_y0y1_gf4_mul_0_1_n66, mul_y0y1_gf4_mul_0_1_n65,
         mul_y0y1_gf4_mul_0_1_n64, mul_y0y1_gf4_mul_0_1_n63,
         mul_y0y1_gf4_mul_0_1_n62, mul_y0y1_gf4_mul_0_1_n61,
         mul_y0y1_gf4_mul_0_1_n60, mul_y0y1_gf4_mul_0_1_n59,
         mul_y0y1_gf4_mul_0_1_n58, mul_y0y1_gf4_mul_0_1_n57,
         mul_y0y1_gf4_mul_0_1_n56, mul_y0y1_gf4_mul_0_1_n55,
         mul_y0y1_gf4_mul_0_1_n54, mul_y0y1_gf4_mul_0_1_n53,
         mul_y0y1_gf4_mul_0_0_n77, mul_y0y1_gf4_mul_0_0_n76,
         mul_y0y1_gf4_mul_0_0_n75, mul_y0y1_gf4_mul_0_0_n74,
         mul_y0y1_gf4_mul_0_0_n73, mul_y0y1_gf4_mul_0_0_n72,
         mul_y0y1_gf4_mul_0_0_n71, mul_y0y1_gf4_mul_0_0_n70,
         mul_y0y1_gf4_mul_0_0_n69, mul_y0y1_gf4_mul_0_0_n68,
         mul_y0y1_gf4_mul_0_0_n67, mul_y0y1_gf4_mul_0_0_n66,
         mul_y0y1_gf4_mul_0_0_n65, mul_y0y1_gf4_mul_0_0_n64,
         mul_y0y1_gf4_mul_0_0_n63, mul_y0y1_gf4_mul_0_0_n62,
         mul_y0y1_gf4_mul_0_0_n61, mul_y0y1_gf4_mul_0_0_n60,
         mul_y0y1_gf4_mul_0_0_n59, mul_y0y1_gf4_mul_0_0_n58,
         mul_y0y1_gf4_mul_0_0_n57, mul_y0y1_gf4_mul_0_0_n56,
         mul_y0y1_gf4_mul_0_0_n55, mul_y0y1_gf4_mul_0_0_n54,
         mul_y0y1_gf4_mul_0_0_n53, inverter_gf24_n3, inverter_gf24_n2,
         inverter_gf24_n1, inverter_gf24_n12, inverter_gf24_n11,
         inverter_gf24_n10, inverter_gf24_n9, inverter_gf24_n8,
         inverter_gf24_n7, inverter_gf24_n6, inverter_gf24_n5,
         inverter_gf24_n4, inverter_gf24_d_0__0_, inverter_gf24_d_1__0_,
         inverter_gf24_d_2__0_, inverter_gf24_ExDP_0__0_,
         inverter_gf24_ExDP_0__1_, inverter_gf24_ExDP_1__0_,
         inverter_gf24_ExDP_1__1_, inverter_gf24_ExDP_2__0_,
         inverter_gf24_ExDP_2__1_, inverter_gf24_a_mul_b_n6,
         inverter_gf24_a_mul_b_n5, inverter_gf24_a_mul_b_n4,
         inverter_gf24_a_mul_b_n3, inverter_gf24_a_mul_b_n2,
         inverter_gf24_a_mul_b_n1, inverter_gf24_a_mul_b_n24,
         inverter_gf24_a_mul_b_n23, inverter_gf24_a_mul_b_n22,
         inverter_gf24_a_mul_b_n21, inverter_gf24_a_mul_b_n20,
         inverter_gf24_a_mul_b_n19, inverter_gf24_a_mul_b_n18,
         inverter_gf24_a_mul_b_n17, inverter_gf24_a_mul_b_n16,
         inverter_gf24_a_mul_b_n15, inverter_gf24_a_mul_b_n14,
         inverter_gf24_a_mul_b_n13, inverter_gf24_a_mul_b_n12,
         inverter_gf24_a_mul_b_n11, inverter_gf24_a_mul_b_n10,
         inverter_gf24_a_mul_b_n9, inverter_gf24_a_mul_b_n8,
         inverter_gf24_a_mul_b_n7, inverter_gf24_a_mul_b_Xi_mul_Yj_1__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_1__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_2__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_2__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_3__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_3__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_5__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_5__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_6__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_6__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_7__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_7__1_,
         inverter_gf24_a_mul_b_gf2_mul_2_2_n15,
         inverter_gf24_a_mul_b_gf2_mul_2_2_n14,
         inverter_gf24_a_mul_b_gf2_mul_2_2_n13,
         inverter_gf24_a_mul_b_gf2_mul_2_2_n12,
         inverter_gf24_a_mul_b_gf2_mul_2_2_n11,
         inverter_gf24_a_mul_b_gf2_mul_2_1_n15,
         inverter_gf24_a_mul_b_gf2_mul_2_1_n14,
         inverter_gf24_a_mul_b_gf2_mul_2_1_n13,
         inverter_gf24_a_mul_b_gf2_mul_2_1_n12,
         inverter_gf24_a_mul_b_gf2_mul_2_1_n11,
         inverter_gf24_a_mul_b_gf2_mul_2_0_n15,
         inverter_gf24_a_mul_b_gf2_mul_2_0_n14,
         inverter_gf24_a_mul_b_gf2_mul_2_0_n13,
         inverter_gf24_a_mul_b_gf2_mul_2_0_n12,
         inverter_gf24_a_mul_b_gf2_mul_2_0_n11,
         inverter_gf24_a_mul_b_gf2_mul_1_2_n15,
         inverter_gf24_a_mul_b_gf2_mul_1_2_n14,
         inverter_gf24_a_mul_b_gf2_mul_1_2_n13,
         inverter_gf24_a_mul_b_gf2_mul_1_2_n12,
         inverter_gf24_a_mul_b_gf2_mul_1_2_n11,
         inverter_gf24_a_mul_b_gf2_mul_1_1_n15,
         inverter_gf24_a_mul_b_gf2_mul_1_1_n14,
         inverter_gf24_a_mul_b_gf2_mul_1_1_n13,
         inverter_gf24_a_mul_b_gf2_mul_1_1_n12,
         inverter_gf24_a_mul_b_gf2_mul_1_1_n11,
         inverter_gf24_a_mul_b_gf2_mul_1_0_n15,
         inverter_gf24_a_mul_b_gf2_mul_1_0_n14,
         inverter_gf24_a_mul_b_gf2_mul_1_0_n13,
         inverter_gf24_a_mul_b_gf2_mul_1_0_n12,
         inverter_gf24_a_mul_b_gf2_mul_1_0_n11,
         inverter_gf24_a_mul_b_gf2_mul_0_2_n15,
         inverter_gf24_a_mul_b_gf2_mul_0_2_n14,
         inverter_gf24_a_mul_b_gf2_mul_0_2_n13,
         inverter_gf24_a_mul_b_gf2_mul_0_2_n12,
         inverter_gf24_a_mul_b_gf2_mul_0_2_n11,
         inverter_gf24_a_mul_b_gf2_mul_0_1_n15,
         inverter_gf24_a_mul_b_gf2_mul_0_1_n14,
         inverter_gf24_a_mul_b_gf2_mul_0_1_n13,
         inverter_gf24_a_mul_b_gf2_mul_0_1_n12,
         inverter_gf24_a_mul_b_gf2_mul_0_1_n11,
         inverter_gf24_a_mul_b_gf2_mul_0_0_n15,
         inverter_gf24_a_mul_b_gf2_mul_0_0_n14,
         inverter_gf24_a_mul_b_gf2_mul_0_0_n13,
         inverter_gf24_a_mul_b_gf2_mul_0_0_n12,
         inverter_gf24_a_mul_b_gf2_mul_0_0_n11, inverter_gf24_a_mul_e_n39,
         inverter_gf24_a_mul_e_n38, inverter_gf24_a_mul_e_n37,
         inverter_gf24_a_mul_e_n36, inverter_gf24_a_mul_e_n35,
         inverter_gf24_a_mul_e_n34, inverter_gf24_a_mul_e_n27,
         inverter_gf24_a_mul_e_n26, inverter_gf24_a_mul_e_n25,
         inverter_gf24_a_mul_e_n42, inverter_gf24_a_mul_e_n41,
         inverter_gf24_a_mul_e_n40, inverter_gf24_a_mul_e_n24,
         inverter_gf24_a_mul_e_n23, inverter_gf24_a_mul_e_n22,
         inverter_gf24_a_mul_e_n21, inverter_gf24_a_mul_e_n20,
         inverter_gf24_a_mul_e_n19, inverter_gf24_a_mul_e_n18,
         inverter_gf24_a_mul_e_n17, inverter_gf24_a_mul_e_n16,
         inverter_gf24_a_mul_e_n15, inverter_gf24_a_mul_e_n14,
         inverter_gf24_a_mul_e_n13, inverter_gf24_a_mul_e_n12,
         inverter_gf24_a_mul_e_n11, inverter_gf24_a_mul_e_n10,
         inverter_gf24_a_mul_e_n9, inverter_gf24_a_mul_e_n8,
         inverter_gf24_a_mul_e_n7, inverter_gf24_a_mul_e_Xi_mul_Yj_1__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_1__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_2__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_2__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_3__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_3__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_5__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_5__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_6__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_6__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_7__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_7__1_,
         inverter_gf24_a_mul_e_gf2_mul_2_2_n15,
         inverter_gf24_a_mul_e_gf2_mul_2_2_n14,
         inverter_gf24_a_mul_e_gf2_mul_2_2_n13,
         inverter_gf24_a_mul_e_gf2_mul_2_2_n12,
         inverter_gf24_a_mul_e_gf2_mul_2_2_n11,
         inverter_gf24_a_mul_e_gf2_mul_2_1_n15,
         inverter_gf24_a_mul_e_gf2_mul_2_1_n14,
         inverter_gf24_a_mul_e_gf2_mul_2_1_n13,
         inverter_gf24_a_mul_e_gf2_mul_2_1_n12,
         inverter_gf24_a_mul_e_gf2_mul_2_1_n11,
         inverter_gf24_a_mul_e_gf2_mul_2_0_n15,
         inverter_gf24_a_mul_e_gf2_mul_2_0_n14,
         inverter_gf24_a_mul_e_gf2_mul_2_0_n13,
         inverter_gf24_a_mul_e_gf2_mul_2_0_n12,
         inverter_gf24_a_mul_e_gf2_mul_2_0_n11,
         inverter_gf24_a_mul_e_gf2_mul_1_2_n15,
         inverter_gf24_a_mul_e_gf2_mul_1_2_n14,
         inverter_gf24_a_mul_e_gf2_mul_1_2_n13,
         inverter_gf24_a_mul_e_gf2_mul_1_2_n12,
         inverter_gf24_a_mul_e_gf2_mul_1_2_n11,
         inverter_gf24_a_mul_e_gf2_mul_1_1_n15,
         inverter_gf24_a_mul_e_gf2_mul_1_1_n14,
         inverter_gf24_a_mul_e_gf2_mul_1_1_n13,
         inverter_gf24_a_mul_e_gf2_mul_1_1_n12,
         inverter_gf24_a_mul_e_gf2_mul_1_1_n11,
         inverter_gf24_a_mul_e_gf2_mul_1_0_n15,
         inverter_gf24_a_mul_e_gf2_mul_1_0_n14,
         inverter_gf24_a_mul_e_gf2_mul_1_0_n13,
         inverter_gf24_a_mul_e_gf2_mul_1_0_n12,
         inverter_gf24_a_mul_e_gf2_mul_1_0_n11,
         inverter_gf24_a_mul_e_gf2_mul_0_2_n15,
         inverter_gf24_a_mul_e_gf2_mul_0_2_n14,
         inverter_gf24_a_mul_e_gf2_mul_0_2_n13,
         inverter_gf24_a_mul_e_gf2_mul_0_2_n12,
         inverter_gf24_a_mul_e_gf2_mul_0_2_n11,
         inverter_gf24_a_mul_e_gf2_mul_0_1_n15,
         inverter_gf24_a_mul_e_gf2_mul_0_1_n14,
         inverter_gf24_a_mul_e_gf2_mul_0_1_n13,
         inverter_gf24_a_mul_e_gf2_mul_0_1_n12,
         inverter_gf24_a_mul_e_gf2_mul_0_1_n11,
         inverter_gf24_a_mul_e_gf2_mul_0_0_n15,
         inverter_gf24_a_mul_e_gf2_mul_0_0_n14,
         inverter_gf24_a_mul_e_gf2_mul_0_0_n13,
         inverter_gf24_a_mul_e_gf2_mul_0_0_n12,
         inverter_gf24_a_mul_e_gf2_mul_0_0_n11, inverter_gf24_b_mul_e_n39,
         inverter_gf24_b_mul_e_n38, inverter_gf24_b_mul_e_n37,
         inverter_gf24_b_mul_e_n36, inverter_gf24_b_mul_e_n35,
         inverter_gf24_b_mul_e_n34, inverter_gf24_b_mul_e_n27,
         inverter_gf24_b_mul_e_n26, inverter_gf24_b_mul_e_n25,
         inverter_gf24_b_mul_e_n42, inverter_gf24_b_mul_e_n41,
         inverter_gf24_b_mul_e_n40, inverter_gf24_b_mul_e_n24,
         inverter_gf24_b_mul_e_n23, inverter_gf24_b_mul_e_n22,
         inverter_gf24_b_mul_e_n21, inverter_gf24_b_mul_e_n20,
         inverter_gf24_b_mul_e_n19, inverter_gf24_b_mul_e_n18,
         inverter_gf24_b_mul_e_n17, inverter_gf24_b_mul_e_n16,
         inverter_gf24_b_mul_e_n15, inverter_gf24_b_mul_e_n14,
         inverter_gf24_b_mul_e_n13, inverter_gf24_b_mul_e_n12,
         inverter_gf24_b_mul_e_n11, inverter_gf24_b_mul_e_n10,
         inverter_gf24_b_mul_e_n9, inverter_gf24_b_mul_e_n8,
         inverter_gf24_b_mul_e_n7, inverter_gf24_b_mul_e_Xi_mul_Yj_1__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_1__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_2__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_2__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_3__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_3__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_5__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_5__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_6__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_6__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_7__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_7__1_,
         inverter_gf24_b_mul_e_gf2_mul_2_2_n15,
         inverter_gf24_b_mul_e_gf2_mul_2_2_n14,
         inverter_gf24_b_mul_e_gf2_mul_2_2_n13,
         inverter_gf24_b_mul_e_gf2_mul_2_2_n12,
         inverter_gf24_b_mul_e_gf2_mul_2_2_n11,
         inverter_gf24_b_mul_e_gf2_mul_2_1_n15,
         inverter_gf24_b_mul_e_gf2_mul_2_1_n14,
         inverter_gf24_b_mul_e_gf2_mul_2_1_n13,
         inverter_gf24_b_mul_e_gf2_mul_2_1_n12,
         inverter_gf24_b_mul_e_gf2_mul_2_1_n11,
         inverter_gf24_b_mul_e_gf2_mul_2_0_n15,
         inverter_gf24_b_mul_e_gf2_mul_2_0_n14,
         inverter_gf24_b_mul_e_gf2_mul_2_0_n13,
         inverter_gf24_b_mul_e_gf2_mul_2_0_n12,
         inverter_gf24_b_mul_e_gf2_mul_2_0_n11,
         inverter_gf24_b_mul_e_gf2_mul_1_2_n15,
         inverter_gf24_b_mul_e_gf2_mul_1_2_n14,
         inverter_gf24_b_mul_e_gf2_mul_1_2_n13,
         inverter_gf24_b_mul_e_gf2_mul_1_2_n12,
         inverter_gf24_b_mul_e_gf2_mul_1_2_n11,
         inverter_gf24_b_mul_e_gf2_mul_1_1_n15,
         inverter_gf24_b_mul_e_gf2_mul_1_1_n14,
         inverter_gf24_b_mul_e_gf2_mul_1_1_n13,
         inverter_gf24_b_mul_e_gf2_mul_1_1_n12,
         inverter_gf24_b_mul_e_gf2_mul_1_1_n11,
         inverter_gf24_b_mul_e_gf2_mul_1_0_n15,
         inverter_gf24_b_mul_e_gf2_mul_1_0_n14,
         inverter_gf24_b_mul_e_gf2_mul_1_0_n13,
         inverter_gf24_b_mul_e_gf2_mul_1_0_n12,
         inverter_gf24_b_mul_e_gf2_mul_1_0_n11,
         inverter_gf24_b_mul_e_gf2_mul_0_2_n15,
         inverter_gf24_b_mul_e_gf2_mul_0_2_n14,
         inverter_gf24_b_mul_e_gf2_mul_0_2_n13,
         inverter_gf24_b_mul_e_gf2_mul_0_2_n12,
         inverter_gf24_b_mul_e_gf2_mul_0_2_n11,
         inverter_gf24_b_mul_e_gf2_mul_0_1_n15,
         inverter_gf24_b_mul_e_gf2_mul_0_1_n14,
         inverter_gf24_b_mul_e_gf2_mul_0_1_n13,
         inverter_gf24_b_mul_e_gf2_mul_0_1_n12,
         inverter_gf24_b_mul_e_gf2_mul_0_1_n11,
         inverter_gf24_b_mul_e_gf2_mul_0_0_n15,
         inverter_gf24_b_mul_e_gf2_mul_0_0_n14,
         inverter_gf24_b_mul_e_gf2_mul_0_0_n13,
         inverter_gf24_b_mul_e_gf2_mul_0_0_n12,
         inverter_gf24_b_mul_e_gf2_mul_0_0_n11, mult_msb_n60, mult_msb_n59,
         mult_msb_n58, mult_msb_n57, mult_msb_n56, mult_msb_n55, mult_msb_n54,
         mult_msb_n53, mult_msb_n52, mult_msb_n51, mult_msb_n50, mult_msb_n49,
         mult_msb_n48, mult_msb_n47, mult_msb_n46, mult_msb_n45, mult_msb_n44,
         mult_msb_n43, mult_msb_n42, mult_msb_n41, mult_msb_n40, mult_msb_n39,
         mult_msb_n38, mult_msb_n37, mult_msb_n36, mult_msb_n35, mult_msb_n34,
         mult_msb_n33, mult_msb_n32, mult_msb_n31, mult_msb_n30, mult_msb_n29,
         mult_msb_n28, mult_msb_n27, mult_msb_n26, mult_msb_n25, mult_msb_n24,
         mult_msb_n23, mult_msb_n22, mult_msb_n21, mult_msb_n20, mult_msb_n19,
         mult_msb_n18, mult_msb_n17, mult_msb_n16, mult_msb_n15, mult_msb_n14,
         mult_msb_n13, mult_msb_Xi_mul_Yj_1__0_, mult_msb_Xi_mul_Yj_1__1_,
         mult_msb_Xi_mul_Yj_1__2_, mult_msb_Xi_mul_Yj_1__3_,
         mult_msb_Xi_mul_Yj_2__0_, mult_msb_Xi_mul_Yj_2__1_,
         mult_msb_Xi_mul_Yj_2__2_, mult_msb_Xi_mul_Yj_2__3_,
         mult_msb_Xi_mul_Yj_3__0_, mult_msb_Xi_mul_Yj_3__1_,
         mult_msb_Xi_mul_Yj_3__2_, mult_msb_Xi_mul_Yj_3__3_,
         mult_msb_Xi_mul_Yj_5__0_, mult_msb_Xi_mul_Yj_5__1_,
         mult_msb_Xi_mul_Yj_5__2_, mult_msb_Xi_mul_Yj_5__3_,
         mult_msb_Xi_mul_Yj_6__0_, mult_msb_Xi_mul_Yj_6__1_,
         mult_msb_Xi_mul_Yj_6__2_, mult_msb_Xi_mul_Yj_6__3_,
         mult_msb_Xi_mul_Yj_7__0_, mult_msb_Xi_mul_Yj_7__1_,
         mult_msb_Xi_mul_Yj_7__2_, mult_msb_Xi_mul_Yj_7__3_,
         mult_msb_gf4_mul_2_2_n77, mult_msb_gf4_mul_2_2_n76,
         mult_msb_gf4_mul_2_2_n75, mult_msb_gf4_mul_2_2_n74,
         mult_msb_gf4_mul_2_2_n73, mult_msb_gf4_mul_2_2_n72,
         mult_msb_gf4_mul_2_2_n71, mult_msb_gf4_mul_2_2_n70,
         mult_msb_gf4_mul_2_2_n69, mult_msb_gf4_mul_2_2_n68,
         mult_msb_gf4_mul_2_2_n67, mult_msb_gf4_mul_2_2_n66,
         mult_msb_gf4_mul_2_2_n65, mult_msb_gf4_mul_2_2_n64,
         mult_msb_gf4_mul_2_2_n63, mult_msb_gf4_mul_2_2_n62,
         mult_msb_gf4_mul_2_2_n61, mult_msb_gf4_mul_2_2_n60,
         mult_msb_gf4_mul_2_2_n59, mult_msb_gf4_mul_2_2_n58,
         mult_msb_gf4_mul_2_2_n57, mult_msb_gf4_mul_2_2_n56,
         mult_msb_gf4_mul_2_2_n55, mult_msb_gf4_mul_2_2_n54,
         mult_msb_gf4_mul_2_2_n53, mult_msb_gf4_mul_2_1_n77,
         mult_msb_gf4_mul_2_1_n76, mult_msb_gf4_mul_2_1_n75,
         mult_msb_gf4_mul_2_1_n74, mult_msb_gf4_mul_2_1_n73,
         mult_msb_gf4_mul_2_1_n72, mult_msb_gf4_mul_2_1_n71,
         mult_msb_gf4_mul_2_1_n70, mult_msb_gf4_mul_2_1_n69,
         mult_msb_gf4_mul_2_1_n68, mult_msb_gf4_mul_2_1_n67,
         mult_msb_gf4_mul_2_1_n66, mult_msb_gf4_mul_2_1_n65,
         mult_msb_gf4_mul_2_1_n64, mult_msb_gf4_mul_2_1_n63,
         mult_msb_gf4_mul_2_1_n62, mult_msb_gf4_mul_2_1_n61,
         mult_msb_gf4_mul_2_1_n60, mult_msb_gf4_mul_2_1_n59,
         mult_msb_gf4_mul_2_1_n58, mult_msb_gf4_mul_2_1_n57,
         mult_msb_gf4_mul_2_1_n56, mult_msb_gf4_mul_2_1_n55,
         mult_msb_gf4_mul_2_1_n54, mult_msb_gf4_mul_2_1_n53,
         mult_msb_gf4_mul_2_0_n77, mult_msb_gf4_mul_2_0_n76,
         mult_msb_gf4_mul_2_0_n75, mult_msb_gf4_mul_2_0_n74,
         mult_msb_gf4_mul_2_0_n73, mult_msb_gf4_mul_2_0_n72,
         mult_msb_gf4_mul_2_0_n71, mult_msb_gf4_mul_2_0_n70,
         mult_msb_gf4_mul_2_0_n69, mult_msb_gf4_mul_2_0_n68,
         mult_msb_gf4_mul_2_0_n67, mult_msb_gf4_mul_2_0_n66,
         mult_msb_gf4_mul_2_0_n65, mult_msb_gf4_mul_2_0_n64,
         mult_msb_gf4_mul_2_0_n63, mult_msb_gf4_mul_2_0_n62,
         mult_msb_gf4_mul_2_0_n61, mult_msb_gf4_mul_2_0_n60,
         mult_msb_gf4_mul_2_0_n59, mult_msb_gf4_mul_2_0_n58,
         mult_msb_gf4_mul_2_0_n57, mult_msb_gf4_mul_2_0_n56,
         mult_msb_gf4_mul_2_0_n55, mult_msb_gf4_mul_2_0_n54,
         mult_msb_gf4_mul_2_0_n53, mult_msb_gf4_mul_1_2_n77,
         mult_msb_gf4_mul_1_2_n76, mult_msb_gf4_mul_1_2_n75,
         mult_msb_gf4_mul_1_2_n74, mult_msb_gf4_mul_1_2_n73,
         mult_msb_gf4_mul_1_2_n72, mult_msb_gf4_mul_1_2_n71,
         mult_msb_gf4_mul_1_2_n70, mult_msb_gf4_mul_1_2_n69,
         mult_msb_gf4_mul_1_2_n68, mult_msb_gf4_mul_1_2_n67,
         mult_msb_gf4_mul_1_2_n66, mult_msb_gf4_mul_1_2_n65,
         mult_msb_gf4_mul_1_2_n64, mult_msb_gf4_mul_1_2_n63,
         mult_msb_gf4_mul_1_2_n62, mult_msb_gf4_mul_1_2_n61,
         mult_msb_gf4_mul_1_2_n60, mult_msb_gf4_mul_1_2_n59,
         mult_msb_gf4_mul_1_2_n58, mult_msb_gf4_mul_1_2_n57,
         mult_msb_gf4_mul_1_2_n56, mult_msb_gf4_mul_1_2_n55,
         mult_msb_gf4_mul_1_2_n54, mult_msb_gf4_mul_1_2_n53,
         mult_msb_gf4_mul_1_1_n77, mult_msb_gf4_mul_1_1_n76,
         mult_msb_gf4_mul_1_1_n75, mult_msb_gf4_mul_1_1_n74,
         mult_msb_gf4_mul_1_1_n73, mult_msb_gf4_mul_1_1_n72,
         mult_msb_gf4_mul_1_1_n71, mult_msb_gf4_mul_1_1_n70,
         mult_msb_gf4_mul_1_1_n69, mult_msb_gf4_mul_1_1_n68,
         mult_msb_gf4_mul_1_1_n67, mult_msb_gf4_mul_1_1_n66,
         mult_msb_gf4_mul_1_1_n65, mult_msb_gf4_mul_1_1_n64,
         mult_msb_gf4_mul_1_1_n63, mult_msb_gf4_mul_1_1_n62,
         mult_msb_gf4_mul_1_1_n61, mult_msb_gf4_mul_1_1_n60,
         mult_msb_gf4_mul_1_1_n59, mult_msb_gf4_mul_1_1_n58,
         mult_msb_gf4_mul_1_1_n57, mult_msb_gf4_mul_1_1_n56,
         mult_msb_gf4_mul_1_1_n55, mult_msb_gf4_mul_1_1_n54,
         mult_msb_gf4_mul_1_1_n53, mult_msb_gf4_mul_1_0_n77,
         mult_msb_gf4_mul_1_0_n76, mult_msb_gf4_mul_1_0_n75,
         mult_msb_gf4_mul_1_0_n74, mult_msb_gf4_mul_1_0_n73,
         mult_msb_gf4_mul_1_0_n72, mult_msb_gf4_mul_1_0_n71,
         mult_msb_gf4_mul_1_0_n70, mult_msb_gf4_mul_1_0_n69,
         mult_msb_gf4_mul_1_0_n68, mult_msb_gf4_mul_1_0_n67,
         mult_msb_gf4_mul_1_0_n66, mult_msb_gf4_mul_1_0_n65,
         mult_msb_gf4_mul_1_0_n64, mult_msb_gf4_mul_1_0_n63,
         mult_msb_gf4_mul_1_0_n62, mult_msb_gf4_mul_1_0_n61,
         mult_msb_gf4_mul_1_0_n60, mult_msb_gf4_mul_1_0_n59,
         mult_msb_gf4_mul_1_0_n58, mult_msb_gf4_mul_1_0_n57,
         mult_msb_gf4_mul_1_0_n56, mult_msb_gf4_mul_1_0_n55,
         mult_msb_gf4_mul_1_0_n54, mult_msb_gf4_mul_1_0_n53,
         mult_msb_gf4_mul_0_2_n77, mult_msb_gf4_mul_0_2_n76,
         mult_msb_gf4_mul_0_2_n75, mult_msb_gf4_mul_0_2_n74,
         mult_msb_gf4_mul_0_2_n73, mult_msb_gf4_mul_0_2_n72,
         mult_msb_gf4_mul_0_2_n71, mult_msb_gf4_mul_0_2_n70,
         mult_msb_gf4_mul_0_2_n69, mult_msb_gf4_mul_0_2_n68,
         mult_msb_gf4_mul_0_2_n67, mult_msb_gf4_mul_0_2_n66,
         mult_msb_gf4_mul_0_2_n65, mult_msb_gf4_mul_0_2_n64,
         mult_msb_gf4_mul_0_2_n63, mult_msb_gf4_mul_0_2_n62,
         mult_msb_gf4_mul_0_2_n61, mult_msb_gf4_mul_0_2_n60,
         mult_msb_gf4_mul_0_2_n59, mult_msb_gf4_mul_0_2_n58,
         mult_msb_gf4_mul_0_2_n57, mult_msb_gf4_mul_0_2_n56,
         mult_msb_gf4_mul_0_2_n55, mult_msb_gf4_mul_0_2_n54,
         mult_msb_gf4_mul_0_2_n53, mult_msb_gf4_mul_0_1_n77,
         mult_msb_gf4_mul_0_1_n76, mult_msb_gf4_mul_0_1_n75,
         mult_msb_gf4_mul_0_1_n74, mult_msb_gf4_mul_0_1_n73,
         mult_msb_gf4_mul_0_1_n72, mult_msb_gf4_mul_0_1_n71,
         mult_msb_gf4_mul_0_1_n70, mult_msb_gf4_mul_0_1_n69,
         mult_msb_gf4_mul_0_1_n68, mult_msb_gf4_mul_0_1_n67,
         mult_msb_gf4_mul_0_1_n66, mult_msb_gf4_mul_0_1_n65,
         mult_msb_gf4_mul_0_1_n64, mult_msb_gf4_mul_0_1_n63,
         mult_msb_gf4_mul_0_1_n62, mult_msb_gf4_mul_0_1_n61,
         mult_msb_gf4_mul_0_1_n60, mult_msb_gf4_mul_0_1_n59,
         mult_msb_gf4_mul_0_1_n58, mult_msb_gf4_mul_0_1_n57,
         mult_msb_gf4_mul_0_1_n56, mult_msb_gf4_mul_0_1_n55,
         mult_msb_gf4_mul_0_1_n54, mult_msb_gf4_mul_0_1_n53,
         mult_msb_gf4_mul_0_0_n77, mult_msb_gf4_mul_0_0_n76,
         mult_msb_gf4_mul_0_0_n75, mult_msb_gf4_mul_0_0_n74,
         mult_msb_gf4_mul_0_0_n73, mult_msb_gf4_mul_0_0_n72,
         mult_msb_gf4_mul_0_0_n71, mult_msb_gf4_mul_0_0_n70,
         mult_msb_gf4_mul_0_0_n69, mult_msb_gf4_mul_0_0_n68,
         mult_msb_gf4_mul_0_0_n67, mult_msb_gf4_mul_0_0_n66,
         mult_msb_gf4_mul_0_0_n65, mult_msb_gf4_mul_0_0_n64,
         mult_msb_gf4_mul_0_0_n63, mult_msb_gf4_mul_0_0_n62,
         mult_msb_gf4_mul_0_0_n61, mult_msb_gf4_mul_0_0_n60,
         mult_msb_gf4_mul_0_0_n59, mult_msb_gf4_mul_0_0_n58,
         mult_msb_gf4_mul_0_0_n57, mult_msb_gf4_mul_0_0_n56,
         mult_msb_gf4_mul_0_0_n55, mult_msb_gf4_mul_0_0_n54,
         mult_msb_gf4_mul_0_0_n53, mult_lsb_n96, mult_lsb_n95, mult_lsb_n94,
         mult_lsb_n93, mult_lsb_n92, mult_lsb_n91, mult_lsb_n90, mult_lsb_n89,
         mult_lsb_n88, mult_lsb_n87, mult_lsb_n86, mult_lsb_n85, mult_lsb_n84,
         mult_lsb_n83, mult_lsb_n82, mult_lsb_n81, mult_lsb_n80, mult_lsb_n79,
         mult_lsb_n78, mult_lsb_n77, mult_lsb_n76, mult_lsb_n75, mult_lsb_n74,
         mult_lsb_n73, mult_lsb_n72, mult_lsb_n71, mult_lsb_n70, mult_lsb_n69,
         mult_lsb_n68, mult_lsb_n67, mult_lsb_n66, mult_lsb_n65, mult_lsb_n64,
         mult_lsb_n63, mult_lsb_n62, mult_lsb_n61, mult_lsb_n60, mult_lsb_n59,
         mult_lsb_n58, mult_lsb_n57, mult_lsb_n56, mult_lsb_n55, mult_lsb_n54,
         mult_lsb_n53, mult_lsb_n52, mult_lsb_n51, mult_lsb_n50, mult_lsb_n49,
         mult_lsb_Xi_mul_Yj_1__0_, mult_lsb_Xi_mul_Yj_1__1_,
         mult_lsb_Xi_mul_Yj_1__2_, mult_lsb_Xi_mul_Yj_1__3_,
         mult_lsb_Xi_mul_Yj_2__0_, mult_lsb_Xi_mul_Yj_2__1_,
         mult_lsb_Xi_mul_Yj_2__2_, mult_lsb_Xi_mul_Yj_2__3_,
         mult_lsb_Xi_mul_Yj_3__0_, mult_lsb_Xi_mul_Yj_3__1_,
         mult_lsb_Xi_mul_Yj_3__2_, mult_lsb_Xi_mul_Yj_3__3_,
         mult_lsb_Xi_mul_Yj_5__0_, mult_lsb_Xi_mul_Yj_5__1_,
         mult_lsb_Xi_mul_Yj_5__2_, mult_lsb_Xi_mul_Yj_5__3_,
         mult_lsb_Xi_mul_Yj_6__0_, mult_lsb_Xi_mul_Yj_6__1_,
         mult_lsb_Xi_mul_Yj_6__2_, mult_lsb_Xi_mul_Yj_6__3_,
         mult_lsb_Xi_mul_Yj_7__0_, mult_lsb_Xi_mul_Yj_7__1_,
         mult_lsb_Xi_mul_Yj_7__2_, mult_lsb_Xi_mul_Yj_7__3_,
         mult_lsb_gf4_mul_2_2_n77, mult_lsb_gf4_mul_2_2_n76,
         mult_lsb_gf4_mul_2_2_n75, mult_lsb_gf4_mul_2_2_n74,
         mult_lsb_gf4_mul_2_2_n73, mult_lsb_gf4_mul_2_2_n72,
         mult_lsb_gf4_mul_2_2_n71, mult_lsb_gf4_mul_2_2_n70,
         mult_lsb_gf4_mul_2_2_n69, mult_lsb_gf4_mul_2_2_n68,
         mult_lsb_gf4_mul_2_2_n67, mult_lsb_gf4_mul_2_2_n66,
         mult_lsb_gf4_mul_2_2_n65, mult_lsb_gf4_mul_2_2_n64,
         mult_lsb_gf4_mul_2_2_n63, mult_lsb_gf4_mul_2_2_n62,
         mult_lsb_gf4_mul_2_2_n61, mult_lsb_gf4_mul_2_2_n60,
         mult_lsb_gf4_mul_2_2_n59, mult_lsb_gf4_mul_2_2_n58,
         mult_lsb_gf4_mul_2_2_n57, mult_lsb_gf4_mul_2_2_n56,
         mult_lsb_gf4_mul_2_2_n55, mult_lsb_gf4_mul_2_2_n54,
         mult_lsb_gf4_mul_2_2_n53, mult_lsb_gf4_mul_2_1_n77,
         mult_lsb_gf4_mul_2_1_n76, mult_lsb_gf4_mul_2_1_n75,
         mult_lsb_gf4_mul_2_1_n74, mult_lsb_gf4_mul_2_1_n73,
         mult_lsb_gf4_mul_2_1_n72, mult_lsb_gf4_mul_2_1_n71,
         mult_lsb_gf4_mul_2_1_n70, mult_lsb_gf4_mul_2_1_n69,
         mult_lsb_gf4_mul_2_1_n68, mult_lsb_gf4_mul_2_1_n67,
         mult_lsb_gf4_mul_2_1_n66, mult_lsb_gf4_mul_2_1_n65,
         mult_lsb_gf4_mul_2_1_n64, mult_lsb_gf4_mul_2_1_n63,
         mult_lsb_gf4_mul_2_1_n62, mult_lsb_gf4_mul_2_1_n61,
         mult_lsb_gf4_mul_2_1_n60, mult_lsb_gf4_mul_2_1_n59,
         mult_lsb_gf4_mul_2_1_n58, mult_lsb_gf4_mul_2_1_n57,
         mult_lsb_gf4_mul_2_1_n56, mult_lsb_gf4_mul_2_1_n55,
         mult_lsb_gf4_mul_2_1_n54, mult_lsb_gf4_mul_2_1_n53,
         mult_lsb_gf4_mul_2_0_n77, mult_lsb_gf4_mul_2_0_n76,
         mult_lsb_gf4_mul_2_0_n75, mult_lsb_gf4_mul_2_0_n74,
         mult_lsb_gf4_mul_2_0_n73, mult_lsb_gf4_mul_2_0_n72,
         mult_lsb_gf4_mul_2_0_n71, mult_lsb_gf4_mul_2_0_n70,
         mult_lsb_gf4_mul_2_0_n69, mult_lsb_gf4_mul_2_0_n68,
         mult_lsb_gf4_mul_2_0_n67, mult_lsb_gf4_mul_2_0_n66,
         mult_lsb_gf4_mul_2_0_n65, mult_lsb_gf4_mul_2_0_n64,
         mult_lsb_gf4_mul_2_0_n63, mult_lsb_gf4_mul_2_0_n62,
         mult_lsb_gf4_mul_2_0_n61, mult_lsb_gf4_mul_2_0_n60,
         mult_lsb_gf4_mul_2_0_n59, mult_lsb_gf4_mul_2_0_n58,
         mult_lsb_gf4_mul_2_0_n57, mult_lsb_gf4_mul_2_0_n56,
         mult_lsb_gf4_mul_2_0_n55, mult_lsb_gf4_mul_2_0_n54,
         mult_lsb_gf4_mul_2_0_n53, mult_lsb_gf4_mul_1_2_n77,
         mult_lsb_gf4_mul_1_2_n76, mult_lsb_gf4_mul_1_2_n75,
         mult_lsb_gf4_mul_1_2_n74, mult_lsb_gf4_mul_1_2_n73,
         mult_lsb_gf4_mul_1_2_n72, mult_lsb_gf4_mul_1_2_n71,
         mult_lsb_gf4_mul_1_2_n70, mult_lsb_gf4_mul_1_2_n69,
         mult_lsb_gf4_mul_1_2_n68, mult_lsb_gf4_mul_1_2_n67,
         mult_lsb_gf4_mul_1_2_n66, mult_lsb_gf4_mul_1_2_n65,
         mult_lsb_gf4_mul_1_2_n64, mult_lsb_gf4_mul_1_2_n63,
         mult_lsb_gf4_mul_1_2_n62, mult_lsb_gf4_mul_1_2_n61,
         mult_lsb_gf4_mul_1_2_n60, mult_lsb_gf4_mul_1_2_n59,
         mult_lsb_gf4_mul_1_2_n58, mult_lsb_gf4_mul_1_2_n57,
         mult_lsb_gf4_mul_1_2_n56, mult_lsb_gf4_mul_1_2_n55,
         mult_lsb_gf4_mul_1_2_n54, mult_lsb_gf4_mul_1_2_n53,
         mult_lsb_gf4_mul_1_1_n77, mult_lsb_gf4_mul_1_1_n76,
         mult_lsb_gf4_mul_1_1_n75, mult_lsb_gf4_mul_1_1_n74,
         mult_lsb_gf4_mul_1_1_n73, mult_lsb_gf4_mul_1_1_n72,
         mult_lsb_gf4_mul_1_1_n71, mult_lsb_gf4_mul_1_1_n70,
         mult_lsb_gf4_mul_1_1_n69, mult_lsb_gf4_mul_1_1_n68,
         mult_lsb_gf4_mul_1_1_n67, mult_lsb_gf4_mul_1_1_n66,
         mult_lsb_gf4_mul_1_1_n65, mult_lsb_gf4_mul_1_1_n64,
         mult_lsb_gf4_mul_1_1_n63, mult_lsb_gf4_mul_1_1_n62,
         mult_lsb_gf4_mul_1_1_n61, mult_lsb_gf4_mul_1_1_n60,
         mult_lsb_gf4_mul_1_1_n59, mult_lsb_gf4_mul_1_1_n58,
         mult_lsb_gf4_mul_1_1_n57, mult_lsb_gf4_mul_1_1_n56,
         mult_lsb_gf4_mul_1_1_n55, mult_lsb_gf4_mul_1_1_n54,
         mult_lsb_gf4_mul_1_1_n53, mult_lsb_gf4_mul_1_0_n77,
         mult_lsb_gf4_mul_1_0_n76, mult_lsb_gf4_mul_1_0_n75,
         mult_lsb_gf4_mul_1_0_n74, mult_lsb_gf4_mul_1_0_n73,
         mult_lsb_gf4_mul_1_0_n72, mult_lsb_gf4_mul_1_0_n71,
         mult_lsb_gf4_mul_1_0_n70, mult_lsb_gf4_mul_1_0_n69,
         mult_lsb_gf4_mul_1_0_n68, mult_lsb_gf4_mul_1_0_n67,
         mult_lsb_gf4_mul_1_0_n66, mult_lsb_gf4_mul_1_0_n65,
         mult_lsb_gf4_mul_1_0_n64, mult_lsb_gf4_mul_1_0_n63,
         mult_lsb_gf4_mul_1_0_n62, mult_lsb_gf4_mul_1_0_n61,
         mult_lsb_gf4_mul_1_0_n60, mult_lsb_gf4_mul_1_0_n59,
         mult_lsb_gf4_mul_1_0_n58, mult_lsb_gf4_mul_1_0_n57,
         mult_lsb_gf4_mul_1_0_n56, mult_lsb_gf4_mul_1_0_n55,
         mult_lsb_gf4_mul_1_0_n54, mult_lsb_gf4_mul_1_0_n53,
         mult_lsb_gf4_mul_0_2_n77, mult_lsb_gf4_mul_0_2_n76,
         mult_lsb_gf4_mul_0_2_n75, mult_lsb_gf4_mul_0_2_n74,
         mult_lsb_gf4_mul_0_2_n73, mult_lsb_gf4_mul_0_2_n72,
         mult_lsb_gf4_mul_0_2_n71, mult_lsb_gf4_mul_0_2_n70,
         mult_lsb_gf4_mul_0_2_n69, mult_lsb_gf4_mul_0_2_n68,
         mult_lsb_gf4_mul_0_2_n67, mult_lsb_gf4_mul_0_2_n66,
         mult_lsb_gf4_mul_0_2_n65, mult_lsb_gf4_mul_0_2_n64,
         mult_lsb_gf4_mul_0_2_n63, mult_lsb_gf4_mul_0_2_n62,
         mult_lsb_gf4_mul_0_2_n61, mult_lsb_gf4_mul_0_2_n60,
         mult_lsb_gf4_mul_0_2_n59, mult_lsb_gf4_mul_0_2_n58,
         mult_lsb_gf4_mul_0_2_n57, mult_lsb_gf4_mul_0_2_n56,
         mult_lsb_gf4_mul_0_2_n55, mult_lsb_gf4_mul_0_2_n54,
         mult_lsb_gf4_mul_0_2_n53, mult_lsb_gf4_mul_0_1_n77,
         mult_lsb_gf4_mul_0_1_n76, mult_lsb_gf4_mul_0_1_n75,
         mult_lsb_gf4_mul_0_1_n74, mult_lsb_gf4_mul_0_1_n73,
         mult_lsb_gf4_mul_0_1_n72, mult_lsb_gf4_mul_0_1_n71,
         mult_lsb_gf4_mul_0_1_n70, mult_lsb_gf4_mul_0_1_n69,
         mult_lsb_gf4_mul_0_1_n68, mult_lsb_gf4_mul_0_1_n67,
         mult_lsb_gf4_mul_0_1_n66, mult_lsb_gf4_mul_0_1_n65,
         mult_lsb_gf4_mul_0_1_n64, mult_lsb_gf4_mul_0_1_n63,
         mult_lsb_gf4_mul_0_1_n62, mult_lsb_gf4_mul_0_1_n61,
         mult_lsb_gf4_mul_0_1_n60, mult_lsb_gf4_mul_0_1_n59,
         mult_lsb_gf4_mul_0_1_n58, mult_lsb_gf4_mul_0_1_n57,
         mult_lsb_gf4_mul_0_1_n56, mult_lsb_gf4_mul_0_1_n55,
         mult_lsb_gf4_mul_0_1_n54, mult_lsb_gf4_mul_0_1_n53,
         mult_lsb_gf4_mul_0_0_n77, mult_lsb_gf4_mul_0_0_n76,
         mult_lsb_gf4_mul_0_0_n75, mult_lsb_gf4_mul_0_0_n74,
         mult_lsb_gf4_mul_0_0_n73, mult_lsb_gf4_mul_0_0_n72,
         mult_lsb_gf4_mul_0_0_n71, mult_lsb_gf4_mul_0_0_n70,
         mult_lsb_gf4_mul_0_0_n69, mult_lsb_gf4_mul_0_0_n68,
         mult_lsb_gf4_mul_0_0_n67, mult_lsb_gf4_mul_0_0_n66,
         mult_lsb_gf4_mul_0_0_n65, mult_lsb_gf4_mul_0_0_n64,
         mult_lsb_gf4_mul_0_0_n63, mult_lsb_gf4_mul_0_0_n62,
         mult_lsb_gf4_mul_0_0_n61, mult_lsb_gf4_mul_0_0_n60,
         mult_lsb_gf4_mul_0_0_n59, mult_lsb_gf4_mul_0_0_n58,
         mult_lsb_gf4_mul_0_0_n57, mult_lsb_gf4_mul_0_0_n56,
         mult_lsb_gf4_mul_0_0_n55, mult_lsb_gf4_mul_0_0_n54,
         mult_lsb_gf4_mul_0_0_n53;
  wire   [11:0] Y1xD;
  wire   [11:0] Y0xD;
  wire   [11:0] InverterInxDP;
  wire   [11:0] InverterInxD;
  wire   [11:0] Y0_0xDP;
  wire   [11:0] Y0_1xDP;
  wire   [11:0] Y0_2xDP;
  wire   [11:0] Y0_3xDP;
  wire   [11:0] Y0_4xDP;
  wire   [11:0] Y1_0xDP;
  wire   [11:0] Y1_1xDP;
  wire   [11:0] Y1_2xDP;
  wire   [11:0] Y1_3xDP;
  wire   [11:0] Y1_4xDP;
  wire   [11:0] Y0xorY12xD;
  wire   [8:0] Y0xorY1xD;
  wire   [11:0] Y0mulY1xD;
  wire   [23:0] InvUnmappedxD;
  wire   [11:0] InverterOutxD;
  wire   [35:0] mul_y0y1_FFxDN;
  wire   [5:0] inverter_gf24_AmulBxD;
  wire   [5:0] inverter_gf24_ExD;
  wire   [5:0] inverter_gf24_pipelinedBxDP;
  wire   [5:0] inverter_gf24_pipelinedAxDP;
  wire   [5:0] inverter_gf24_BxDP;
  wire   [5:0] inverter_gf24_AxDP;
  wire   [17:0] inverter_gf24_a_mul_b_FFxDN;
  wire   [17:0] inverter_gf24_a_mul_e_FFxDN;
  wire   [17:0] inverter_gf24_b_mul_e_FFxDN;
  wire   [35:0] mult_msb_FFxDN;
  wire   [35:0] mult_lsb_FFxDN;

  DFF_X1 mappedxDP_reg_2__7_ ( .D(mappedxD_2__7_), .CK(ClkxCI), .Q(Y1xD[11]), 
        .QN(n10) );
  DFF_X1 mappedxDP_reg_2__6_ ( .D(mappedxD_2__6_), .CK(ClkxCI), .Q(Y1xD[10]), 
        .QN(n12) );
  DFF_X1 mappedxDP_reg_2__5_ ( .D(mappedxD_2__5_), .CK(ClkxCI), .Q(Y1xD[9]), 
        .QN(n14) );
  DFF_X1 mappedxDP_reg_2__4_ ( .D(mappedxD_2__4_), .CK(ClkxCI), .Q(Y1xD[8]), 
        .QN(n16) );
  DFF_X1 mappedxDP_reg_2__3_ ( .D(mappedxD_2__3_), .CK(ClkxCI), .Q(Y0xD[11]), 
        .QN(n9) );
  DFF_X1 mappedxDP_reg_2__2_ ( .D(XxDI[16]), .CK(ClkxCI), .Q(Y0xD[10]), .QN(
        n11) );
  DFF_X1 mappedxDP_reg_2__1_ ( .D(mappedxD_2__1_), .CK(ClkxCI), .Q(Y0xD[9]), 
        .QN(n13) );
  DFF_X1 mappedxDP_reg_2__0_ ( .D(mappedxD_2__0_), .CK(ClkxCI), .Q(Y0xD[8]), 
        .QN(n15) );
  DFF_X1 mappedxDP_reg_1__7_ ( .D(mappedxD_1__7_), .CK(ClkxCI), .Q(Y1xD[7]), 
        .QN(n18) );
  DFF_X1 mappedxDP_reg_1__6_ ( .D(mappedxD_1__6_), .CK(ClkxCI), .Q(Y1xD[6]), 
        .QN(n20) );
  DFF_X1 mappedxDP_reg_1__5_ ( .D(mappedxD_1__5_), .CK(ClkxCI), .Q(Y1xD[5]), 
        .QN(n22) );
  DFF_X1 mappedxDP_reg_1__4_ ( .D(mappedxD_1__4_), .CK(ClkxCI), .Q(Y1xD[4]), 
        .QN(n24) );
  DFF_X1 mappedxDP_reg_1__3_ ( .D(mappedxD_1__3_), .CK(ClkxCI), .Q(Y0xD[7]), 
        .QN(n17) );
  DFF_X1 mappedxDP_reg_1__2_ ( .D(XxDI[8]), .CK(ClkxCI), .Q(Y0xD[6]), .QN(n19)
         );
  DFF_X1 mappedxDP_reg_1__1_ ( .D(mappedxD_1__1_), .CK(ClkxCI), .Q(Y0xD[5]), 
        .QN(n21) );
  DFF_X1 mappedxDP_reg_1__0_ ( .D(mappedxD_1__0_), .CK(ClkxCI), .Q(Y0xD[4]), 
        .QN(n23) );
  DFF_X1 mappedxDP_reg_0__7_ ( .D(mappedxD_0__7_), .CK(ClkxCI), .Q(Y1xD[3]), 
        .QN(n26) );
  DFF_X1 mappedxDP_reg_0__6_ ( .D(mappedxD_0__6_), .CK(ClkxCI), .Q(Y1xD[2]), 
        .QN(n28) );
  DFF_X1 mappedxDP_reg_0__5_ ( .D(mappedxD_0__5_), .CK(ClkxCI), .Q(Y1xD[1]), 
        .QN(n30) );
  DFF_X1 mappedxDP_reg_0__4_ ( .D(mappedxD_0__4_), .CK(ClkxCI), .Q(Y1xD[0]), 
        .QN(n32) );
  DFF_X1 mappedxDP_reg_0__3_ ( .D(mappedxD_0__3_), .CK(ClkxCI), .Q(Y0xD[3]), 
        .QN(n25) );
  DFF_X1 mappedxDP_reg_0__2_ ( .D(XxDI[0]), .CK(ClkxCI), .Q(Y0xD[2]), .QN(n27)
         );
  DFF_X1 mappedxDP_reg_0__1_ ( .D(mappedxD_0__1_), .CK(ClkxCI), .Q(Y0xD[1]), 
        .QN(n29) );
  DFF_X1 mappedxDP_reg_0__0_ ( .D(mappedxD_0__0_), .CK(ClkxCI), .Q(Y0xD[0]), 
        .QN(n31) );
  DFF_X1 Y0xorY12xDP_reg_2__3_ ( .D(Y0xorY12xD[11]), .CK(ClkxCI), .Q(), .QN(
        n33) );
  DFF_X1 InverterInxDP_reg_2__3_ ( .D(InverterInxD[11]), .CK(ClkxCI), .Q(
        InverterInxDP[11]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_2__2_ ( .D(Y0xorY12xD[10]), .CK(ClkxCI), .Q(), .QN(
        n34) );
  DFF_X1 InverterInxDP_reg_2__2_ ( .D(InverterInxD[10]), .CK(ClkxCI), .Q(
        InverterInxDP[10]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_2__1_ ( .D(Y0xorY12xD[9]), .CK(ClkxCI), .Q(), .QN(n35) );
  DFF_X1 InverterInxDP_reg_2__1_ ( .D(InverterInxD[9]), .CK(ClkxCI), .Q(
        InverterInxDP[9]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_2__0_ ( .D(Y0xorY12xD[8]), .CK(ClkxCI), .Q(), .QN(n36) );
  DFF_X1 InverterInxDP_reg_2__0_ ( .D(InverterInxD[8]), .CK(ClkxCI), .Q(
        InverterInxDP[8]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_1__3_ ( .D(Y0xorY12xD[7]), .CK(ClkxCI), .Q(), .QN(n37) );
  DFF_X1 InverterInxDP_reg_1__3_ ( .D(InverterInxD[7]), .CK(ClkxCI), .Q(
        InverterInxDP[7]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_1__2_ ( .D(Y0xorY12xD[6]), .CK(ClkxCI), .Q(), .QN(n38) );
  DFF_X1 InverterInxDP_reg_1__2_ ( .D(InverterInxD[6]), .CK(ClkxCI), .Q(
        InverterInxDP[6]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_1__1_ ( .D(Y0xorY12xD[5]), .CK(ClkxCI), .Q(), .QN(n39) );
  DFF_X1 InverterInxDP_reg_1__1_ ( .D(InverterInxD[5]), .CK(ClkxCI), .Q(
        InverterInxDP[5]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_1__0_ ( .D(Y0xorY12xD[4]), .CK(ClkxCI), .Q(), .QN(n40) );
  DFF_X1 InverterInxDP_reg_1__0_ ( .D(InverterInxD[4]), .CK(ClkxCI), .Q(
        InverterInxDP[4]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_0__3_ ( .D(Y0xorY12xD[3]), .CK(ClkxCI), .Q(), .QN(n41) );
  DFF_X1 InverterInxDP_reg_0__3_ ( .D(InverterInxD[3]), .CK(ClkxCI), .Q(
        InverterInxDP[3]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_0__2_ ( .D(Y0xorY12xD[2]), .CK(ClkxCI), .Q(), .QN(n42) );
  DFF_X1 InverterInxDP_reg_0__2_ ( .D(InverterInxD[2]), .CK(ClkxCI), .Q(
        InverterInxDP[2]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_0__1_ ( .D(Y0xorY12xD[1]), .CK(ClkxCI), .Q(), .QN(n43) );
  DFF_X1 InverterInxDP_reg_0__1_ ( .D(InverterInxD[1]), .CK(ClkxCI), .Q(
        InverterInxDP[1]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_0__0_ ( .D(Y0xorY12xD[0]), .CK(ClkxCI), .Q(), .QN(n44) );
  DFF_X1 InverterInxDP_reg_0__0_ ( .D(InverterInxD[0]), .CK(ClkxCI), .Q(
        InverterInxDP[0]), .QN() );
  DFF_X1 Y0_0xDP_reg_2__3_ ( .D(Y0xD[11]), .CK(ClkxCI), .Q(Y0_0xDP[11]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_2__2_ ( .D(Y0xD[10]), .CK(ClkxCI), .Q(Y0_0xDP[10]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_2__1_ ( .D(Y0xD[9]), .CK(ClkxCI), .Q(Y0_0xDP[9]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_2__0_ ( .D(Y0xD[8]), .CK(ClkxCI), .Q(Y0_0xDP[8]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_1__3_ ( .D(Y0xD[7]), .CK(ClkxCI), .Q(Y0_0xDP[7]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_1__2_ ( .D(Y0xD[6]), .CK(ClkxCI), .Q(Y0_0xDP[6]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_1__1_ ( .D(Y0xD[5]), .CK(ClkxCI), .Q(Y0_0xDP[5]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_1__0_ ( .D(Y0xD[4]), .CK(ClkxCI), .Q(Y0_0xDP[4]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_0__3_ ( .D(Y0xD[3]), .CK(ClkxCI), .Q(Y0_0xDP[3]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_0__2_ ( .D(Y0xD[2]), .CK(ClkxCI), .Q(Y0_0xDP[2]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_0__1_ ( .D(Y0xD[1]), .CK(ClkxCI), .Q(Y0_0xDP[1]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_0__0_ ( .D(Y0xD[0]), .CK(ClkxCI), .Q(Y0_0xDP[0]), .QN()
         );
  DFF_X1 Y0_1xDP_reg_2__3_ ( .D(Y0_0xDP[11]), .CK(ClkxCI), .Q(Y0_1xDP[11]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_2__2_ ( .D(Y0_0xDP[10]), .CK(ClkxCI), .Q(Y0_1xDP[10]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_2__1_ ( .D(Y0_0xDP[9]), .CK(ClkxCI), .Q(Y0_1xDP[9]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_2__0_ ( .D(Y0_0xDP[8]), .CK(ClkxCI), .Q(Y0_1xDP[8]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_1__3_ ( .D(Y0_0xDP[7]), .CK(ClkxCI), .Q(Y0_1xDP[7]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_1__2_ ( .D(Y0_0xDP[6]), .CK(ClkxCI), .Q(Y0_1xDP[6]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_1__1_ ( .D(Y0_0xDP[5]), .CK(ClkxCI), .Q(Y0_1xDP[5]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_1__0_ ( .D(Y0_0xDP[4]), .CK(ClkxCI), .Q(Y0_1xDP[4]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_0__3_ ( .D(Y0_0xDP[3]), .CK(ClkxCI), .Q(Y0_1xDP[3]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_0__2_ ( .D(Y0_0xDP[2]), .CK(ClkxCI), .Q(Y0_1xDP[2]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_0__1_ ( .D(Y0_0xDP[1]), .CK(ClkxCI), .Q(Y0_1xDP[1]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_0__0_ ( .D(Y0_0xDP[0]), .CK(ClkxCI), .Q(Y0_1xDP[0]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_2__3_ ( .D(Y0_1xDP[11]), .CK(ClkxCI), .Q(Y0_2xDP[11]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_2__2_ ( .D(Y0_1xDP[10]), .CK(ClkxCI), .Q(Y0_2xDP[10]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_2__1_ ( .D(Y0_1xDP[9]), .CK(ClkxCI), .Q(Y0_2xDP[9]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_2__0_ ( .D(Y0_1xDP[8]), .CK(ClkxCI), .Q(Y0_2xDP[8]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_1__3_ ( .D(Y0_1xDP[7]), .CK(ClkxCI), .Q(Y0_2xDP[7]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_1__2_ ( .D(Y0_1xDP[6]), .CK(ClkxCI), .Q(Y0_2xDP[6]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_1__1_ ( .D(Y0_1xDP[5]), .CK(ClkxCI), .Q(Y0_2xDP[5]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_1__0_ ( .D(Y0_1xDP[4]), .CK(ClkxCI), .Q(Y0_2xDP[4]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_0__3_ ( .D(Y0_1xDP[3]), .CK(ClkxCI), .Q(Y0_2xDP[3]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_0__2_ ( .D(Y0_1xDP[2]), .CK(ClkxCI), .Q(Y0_2xDP[2]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_0__1_ ( .D(Y0_1xDP[1]), .CK(ClkxCI), .Q(Y0_2xDP[1]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_0__0_ ( .D(Y0_1xDP[0]), .CK(ClkxCI), .Q(Y0_2xDP[0]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_2__3_ ( .D(Y0_2xDP[11]), .CK(ClkxCI), .Q(Y0_3xDP[11]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_2__2_ ( .D(Y0_2xDP[10]), .CK(ClkxCI), .Q(Y0_3xDP[10]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_2__1_ ( .D(Y0_2xDP[9]), .CK(ClkxCI), .Q(Y0_3xDP[9]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_2__0_ ( .D(Y0_2xDP[8]), .CK(ClkxCI), .Q(Y0_3xDP[8]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_1__3_ ( .D(Y0_2xDP[7]), .CK(ClkxCI), .Q(Y0_3xDP[7]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_1__2_ ( .D(Y0_2xDP[6]), .CK(ClkxCI), .Q(Y0_3xDP[6]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_1__1_ ( .D(Y0_2xDP[5]), .CK(ClkxCI), .Q(Y0_3xDP[5]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_1__0_ ( .D(Y0_2xDP[4]), .CK(ClkxCI), .Q(Y0_3xDP[4]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_0__3_ ( .D(Y0_2xDP[3]), .CK(ClkxCI), .Q(Y0_3xDP[3]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_0__2_ ( .D(Y0_2xDP[2]), .CK(ClkxCI), .Q(Y0_3xDP[2]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_0__1_ ( .D(Y0_2xDP[1]), .CK(ClkxCI), .Q(Y0_3xDP[1]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_0__0_ ( .D(Y0_2xDP[0]), .CK(ClkxCI), .Q(Y0_3xDP[0]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_2__3_ ( .D(Y0_3xDP[11]), .CK(ClkxCI), .Q(Y0_4xDP[11]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_2__2_ ( .D(Y0_3xDP[10]), .CK(ClkxCI), .Q(Y0_4xDP[10]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_2__1_ ( .D(Y0_3xDP[9]), .CK(ClkxCI), .Q(Y0_4xDP[9]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_2__0_ ( .D(Y0_3xDP[8]), .CK(ClkxCI), .Q(Y0_4xDP[8]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_1__3_ ( .D(Y0_3xDP[7]), .CK(ClkxCI), .Q(Y0_4xDP[7]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_1__2_ ( .D(Y0_3xDP[6]), .CK(ClkxCI), .Q(Y0_4xDP[6]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_1__1_ ( .D(Y0_3xDP[5]), .CK(ClkxCI), .Q(Y0_4xDP[5]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_1__0_ ( .D(Y0_3xDP[4]), .CK(ClkxCI), .Q(Y0_4xDP[4]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_0__3_ ( .D(Y0_3xDP[3]), .CK(ClkxCI), .Q(Y0_4xDP[3]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_0__2_ ( .D(Y0_3xDP[2]), .CK(ClkxCI), .Q(Y0_4xDP[2]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_0__1_ ( .D(Y0_3xDP[1]), .CK(ClkxCI), .Q(Y0_4xDP[1]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_0__0_ ( .D(Y0_3xDP[0]), .CK(ClkxCI), .Q(Y0_4xDP[0]), 
        .QN() );
  DFF_X1 Y1_0xDP_reg_2__3_ ( .D(Y1xD[11]), .CK(ClkxCI), .Q(Y1_0xDP[11]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_2__2_ ( .D(Y1xD[10]), .CK(ClkxCI), .Q(Y1_0xDP[10]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_2__1_ ( .D(Y1xD[9]), .CK(ClkxCI), .Q(Y1_0xDP[9]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_2__0_ ( .D(Y1xD[8]), .CK(ClkxCI), .Q(Y1_0xDP[8]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_1__3_ ( .D(Y1xD[7]), .CK(ClkxCI), .Q(Y1_0xDP[7]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_1__2_ ( .D(Y1xD[6]), .CK(ClkxCI), .Q(Y1_0xDP[6]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_1__1_ ( .D(Y1xD[5]), .CK(ClkxCI), .Q(Y1_0xDP[5]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_1__0_ ( .D(Y1xD[4]), .CK(ClkxCI), .Q(Y1_0xDP[4]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_0__3_ ( .D(Y1xD[3]), .CK(ClkxCI), .Q(Y1_0xDP[3]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_0__2_ ( .D(Y1xD[2]), .CK(ClkxCI), .Q(Y1_0xDP[2]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_0__1_ ( .D(Y1xD[1]), .CK(ClkxCI), .Q(Y1_0xDP[1]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_0__0_ ( .D(Y1xD[0]), .CK(ClkxCI), .Q(Y1_0xDP[0]), .QN()
         );
  DFF_X1 Y1_1xDP_reg_2__3_ ( .D(Y1_0xDP[11]), .CK(ClkxCI), .Q(Y1_1xDP[11]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_2__2_ ( .D(Y1_0xDP[10]), .CK(ClkxCI), .Q(Y1_1xDP[10]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_2__1_ ( .D(Y1_0xDP[9]), .CK(ClkxCI), .Q(Y1_1xDP[9]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_2__0_ ( .D(Y1_0xDP[8]), .CK(ClkxCI), .Q(Y1_1xDP[8]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_1__3_ ( .D(Y1_0xDP[7]), .CK(ClkxCI), .Q(Y1_1xDP[7]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_1__2_ ( .D(Y1_0xDP[6]), .CK(ClkxCI), .Q(Y1_1xDP[6]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_1__1_ ( .D(Y1_0xDP[5]), .CK(ClkxCI), .Q(Y1_1xDP[5]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_1__0_ ( .D(Y1_0xDP[4]), .CK(ClkxCI), .Q(Y1_1xDP[4]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_0__3_ ( .D(Y1_0xDP[3]), .CK(ClkxCI), .Q(Y1_1xDP[3]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_0__2_ ( .D(Y1_0xDP[2]), .CK(ClkxCI), .Q(Y1_1xDP[2]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_0__1_ ( .D(Y1_0xDP[1]), .CK(ClkxCI), .Q(Y1_1xDP[1]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_0__0_ ( .D(Y1_0xDP[0]), .CK(ClkxCI), .Q(Y1_1xDP[0]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_2__3_ ( .D(Y1_1xDP[11]), .CK(ClkxCI), .Q(Y1_2xDP[11]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_2__2_ ( .D(Y1_1xDP[10]), .CK(ClkxCI), .Q(Y1_2xDP[10]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_2__1_ ( .D(Y1_1xDP[9]), .CK(ClkxCI), .Q(Y1_2xDP[9]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_2__0_ ( .D(Y1_1xDP[8]), .CK(ClkxCI), .Q(Y1_2xDP[8]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_1__3_ ( .D(Y1_1xDP[7]), .CK(ClkxCI), .Q(Y1_2xDP[7]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_1__2_ ( .D(Y1_1xDP[6]), .CK(ClkxCI), .Q(Y1_2xDP[6]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_1__1_ ( .D(Y1_1xDP[5]), .CK(ClkxCI), .Q(Y1_2xDP[5]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_1__0_ ( .D(Y1_1xDP[4]), .CK(ClkxCI), .Q(Y1_2xDP[4]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_0__3_ ( .D(Y1_1xDP[3]), .CK(ClkxCI), .Q(Y1_2xDP[3]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_0__2_ ( .D(Y1_1xDP[2]), .CK(ClkxCI), .Q(Y1_2xDP[2]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_0__1_ ( .D(Y1_1xDP[1]), .CK(ClkxCI), .Q(Y1_2xDP[1]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_0__0_ ( .D(Y1_1xDP[0]), .CK(ClkxCI), .Q(Y1_2xDP[0]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_2__3_ ( .D(Y1_2xDP[11]), .CK(ClkxCI), .Q(Y1_3xDP[11]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_2__3_ ( .D(Y1_3xDP[11]), .CK(ClkxCI), .Q(Y1_4xDP[11]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_2__2_ ( .D(Y1_2xDP[10]), .CK(ClkxCI), .Q(Y1_3xDP[10]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_2__2_ ( .D(Y1_3xDP[10]), .CK(ClkxCI), .Q(Y1_4xDP[10]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_2__1_ ( .D(Y1_2xDP[9]), .CK(ClkxCI), .Q(Y1_3xDP[9]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_2__1_ ( .D(Y1_3xDP[9]), .CK(ClkxCI), .Q(Y1_4xDP[9]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_2__0_ ( .D(Y1_2xDP[8]), .CK(ClkxCI), .Q(Y1_3xDP[8]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_2__0_ ( .D(Y1_3xDP[8]), .CK(ClkxCI), .Q(Y1_4xDP[8]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_1__3_ ( .D(Y1_2xDP[7]), .CK(ClkxCI), .Q(Y1_3xDP[7]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_1__3_ ( .D(Y1_3xDP[7]), .CK(ClkxCI), .Q(Y1_4xDP[7]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_1__2_ ( .D(Y1_2xDP[6]), .CK(ClkxCI), .Q(Y1_3xDP[6]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_1__2_ ( .D(Y1_3xDP[6]), .CK(ClkxCI), .Q(Y1_4xDP[6]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_1__1_ ( .D(Y1_2xDP[5]), .CK(ClkxCI), .Q(Y1_3xDP[5]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_1__1_ ( .D(Y1_3xDP[5]), .CK(ClkxCI), .Q(Y1_4xDP[5]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_1__0_ ( .D(Y1_2xDP[4]), .CK(ClkxCI), .Q(Y1_3xDP[4]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_1__0_ ( .D(Y1_3xDP[4]), .CK(ClkxCI), .Q(Y1_4xDP[4]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_0__3_ ( .D(Y1_2xDP[3]), .CK(ClkxCI), .Q(Y1_3xDP[3]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_0__3_ ( .D(Y1_3xDP[3]), .CK(ClkxCI), .Q(Y1_4xDP[3]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_0__2_ ( .D(Y1_2xDP[2]), .CK(ClkxCI), .Q(Y1_3xDP[2]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_0__2_ ( .D(Y1_3xDP[2]), .CK(ClkxCI), .Q(Y1_4xDP[2]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_0__1_ ( .D(Y1_2xDP[1]), .CK(ClkxCI), .Q(Y1_3xDP[1]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_0__1_ ( .D(Y1_3xDP[1]), .CK(ClkxCI), .Q(Y1_4xDP[1]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_0__0_ ( .D(Y1_2xDP[0]), .CK(ClkxCI), .Q(Y1_3xDP[0]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_0__0_ ( .D(Y1_3xDP[0]), .CK(ClkxCI), .Q(Y1_4xDP[0]), 
        .QN() );
  XNOR2_X1 U60 ( .A(Y0mulY1xD[0]), .B(n44), .ZN(InverterInxD[0]) );
  XNOR2_X1 U61 ( .A(Y0mulY1xD[1]), .B(n43), .ZN(InverterInxD[1]) );
  XNOR2_X1 U62 ( .A(Y0mulY1xD[2]), .B(n42), .ZN(InverterInxD[2]) );
  XNOR2_X1 U63 ( .A(Y0mulY1xD[3]), .B(n41), .ZN(InverterInxD[3]) );
  XNOR2_X1 U64 ( .A(Y0mulY1xD[4]), .B(n40), .ZN(InverterInxD[4]) );
  XNOR2_X1 U65 ( .A(Y0mulY1xD[5]), .B(n39), .ZN(InverterInxD[5]) );
  XNOR2_X1 U66 ( .A(Y0mulY1xD[6]), .B(n38), .ZN(InverterInxD[6]) );
  XNOR2_X1 U67 ( .A(Y0mulY1xD[7]), .B(n37), .ZN(InverterInxD[7]) );
  XNOR2_X1 U68 ( .A(Y0mulY1xD[8]), .B(n36), .ZN(InverterInxD[8]) );
  XNOR2_X1 U69 ( .A(Y0mulY1xD[9]), .B(n35), .ZN(InverterInxD[9]) );
  XNOR2_X1 U70 ( .A(Y0mulY1xD[10]), .B(n34), .ZN(InverterInxD[10]) );
  XNOR2_X1 U71 ( .A(Y0mulY1xD[11]), .B(n33), .ZN(InverterInxD[11]) );
  XOR2_X1 U72 ( .A(n32), .B(n31), .Z(Y0xorY12xD[0]) );
  XOR2_X1 U73 ( .A(n30), .B(n29), .Z(Y0xorY1xD[0]) );
  XOR2_X1 U74 ( .A(n28), .B(n27), .Z(Y0xorY1xD[1]) );
  XOR2_X1 U75 ( .A(n26), .B(n25), .Z(Y0xorY1xD[2]) );
  XOR2_X1 U76 ( .A(n24), .B(n23), .Z(Y0xorY12xD[4]) );
  XOR2_X1 U77 ( .A(n22), .B(n21), .Z(Y0xorY1xD[3]) );
  XOR2_X1 U78 ( .A(n20), .B(n19), .Z(Y0xorY1xD[4]) );
  XOR2_X1 U79 ( .A(n18), .B(n17), .Z(Y0xorY1xD[5]) );
  XOR2_X1 U80 ( .A(n16), .B(n15), .Z(Y0xorY12xD[8]) );
  XOR2_X1 U81 ( .A(n14), .B(n13), .Z(Y0xorY1xD[6]) );
  XOR2_X1 U82 ( .A(n12), .B(n11), .Z(Y0xorY1xD[7]) );
  XOR2_X1 U83 ( .A(n10), .B(n9), .Z(Y0xorY1xD[8]) );
  INV_X1 U84 ( .A(InvMappedxD_0__6_), .ZN(QxDO[6]) );
  INV_X1 U85 ( .A(InvMappedxD_0__5_), .ZN(QxDO[5]) );
  INV_X1 U86 ( .A(InvMappedxD_0__1_), .ZN(QxDO[1]) );
  INV_X1 U87 ( .A(InvMappedxD_0__0_), .ZN(QxDO[0]) );
  XNOR2_X1 input_mapping_2_U14 ( .A(input_mapping_2_n23), .B(
        input_mapping_2_n22), .ZN(mappedxD_2__7_) );
  XOR2_X1 input_mapping_2_U13 ( .A(XxDI[20]), .B(mappedxD_2__1_), .Z(
        mappedxD_2__6_) );
  XNOR2_X1 input_mapping_2_U12 ( .A(input_mapping_2_n21), .B(
        input_mapping_2_n20), .ZN(mappedxD_2__5_) );
  XNOR2_X1 input_mapping_2_U11 ( .A(XxDI[16]), .B(input_mapping_2_n22), .ZN(
        mappedxD_2__4_) );
  XNOR2_X1 input_mapping_2_U10 ( .A(XxDI[23]), .B(input_mapping_2_n21), .ZN(
        input_mapping_2_n22) );
  XNOR2_X1 input_mapping_2_U9 ( .A(input_mapping_2_n19), .B(
        input_mapping_2_n18), .ZN(mappedxD_2__3_) );
  XNOR2_X1 input_mapping_2_U8 ( .A(input_mapping_2_n20), .B(XxDI[19]), .ZN(
        input_mapping_2_n18) );
  XNOR2_X1 input_mapping_2_U7 ( .A(XxDI[23]), .B(XxDI[20]), .ZN(
        input_mapping_2_n19) );
  XOR2_X1 input_mapping_2_U6 ( .A(XxDI[16]), .B(input_mapping_2_n21), .Z(
        mappedxD_2__1_) );
  XOR2_X1 input_mapping_2_U5 ( .A(XxDI[22]), .B(XxDI[21]), .Z(
        input_mapping_2_n21) );
  XNOR2_X1 input_mapping_2_U4 ( .A(input_mapping_2_n23), .B(
        input_mapping_2_n17), .ZN(mappedxD_2__0_) );
  XNOR2_X1 input_mapping_2_U3 ( .A(XxDI[22]), .B(XxDI[19]), .ZN(
        input_mapping_2_n17) );
  XNOR2_X1 input_mapping_2_U2 ( .A(XxDI[18]), .B(input_mapping_2_n20), .ZN(
        input_mapping_2_n23) );
  XNOR2_X1 input_mapping_2_U1 ( .A(XxDI[16]), .B(XxDI[17]), .ZN(
        input_mapping_2_n20) );
  XOR2_X1 square_scaler_gf24_2_U3 ( .A(Y0xorY12xD[8]), .B(Y0xorY1xD[7]), .Z(
        Y0xorY12xD[11]) );
  XOR2_X1 square_scaler_gf24_2_U2 ( .A(Y0xorY1xD[6]), .B(Y0xorY1xD[8]), .Z(
        Y0xorY12xD[10]) );
  XOR2_X1 square_scaler_gf24_2_U1 ( .A(Y0xorY12xD[8]), .B(Y0xorY1xD[6]), .Z(
        Y0xorY12xD[9]) );
  XOR2_X1 output_mapping_2_U11 ( .A(InvUnmappedxD[19]), .B(InvUnmappedxD[23]), 
        .Z(QxDO[22]) );
  XNOR2_X1 output_mapping_2_U10 ( .A(QxDO[20]), .B(output_mapping_2_n9), .ZN(
        QxDO[19]) );
  XOR2_X1 output_mapping_2_U9 ( .A(QxDO[23]), .B(InvUnmappedxD[23]), .Z(
        QxDO[20]) );
  XNOR2_X1 output_mapping_2_U8 ( .A(output_mapping_2_n8), .B(QxDO[21]), .ZN(
        QxDO[18]) );
  XNOR2_X1 output_mapping_2_U7 ( .A(QxDO[23]), .B(InvUnmappedxD[18]), .ZN(
        output_mapping_2_n8) );
  XOR2_X1 output_mapping_2_U6 ( .A(InvUnmappedxD[22]), .B(InvUnmappedxD[16]), 
        .Z(QxDO[21]) );
  XOR2_X1 output_mapping_2_U5 ( .A(InvUnmappedxD[19]), .B(InvUnmappedxD[21]), 
        .Z(QxDO[23]) );
  XNOR2_X1 output_mapping_2_U4 ( .A(output_mapping_2_n7), .B(InvUnmappedxD[17]), .ZN(QxDO[17]) );
  XNOR2_X1 output_mapping_2_U3 ( .A(InvUnmappedxD[21]), .B(InvUnmappedxD[20]), 
        .ZN(output_mapping_2_n7) );
  XNOR2_X1 output_mapping_2_U2 ( .A(InvUnmappedxD[17]), .B(output_mapping_2_n9), .ZN(QxDO[16]) );
  XNOR2_X1 output_mapping_2_U1 ( .A(InvUnmappedxD[22]), .B(InvUnmappedxD[20]), 
        .ZN(output_mapping_2_n9) );
  XNOR2_X1 input_mapping_1_U14 ( .A(input_mapping_1_n23), .B(
        input_mapping_1_n22), .ZN(mappedxD_1__7_) );
  XOR2_X1 input_mapping_1_U13 ( .A(XxDI[12]), .B(mappedxD_1__1_), .Z(
        mappedxD_1__6_) );
  XNOR2_X1 input_mapping_1_U12 ( .A(input_mapping_1_n21), .B(
        input_mapping_1_n20), .ZN(mappedxD_1__5_) );
  XNOR2_X1 input_mapping_1_U11 ( .A(XxDI[8]), .B(input_mapping_1_n22), .ZN(
        mappedxD_1__4_) );
  XNOR2_X1 input_mapping_1_U10 ( .A(XxDI[15]), .B(input_mapping_1_n21), .ZN(
        input_mapping_1_n22) );
  XNOR2_X1 input_mapping_1_U9 ( .A(input_mapping_1_n19), .B(
        input_mapping_1_n18), .ZN(mappedxD_1__3_) );
  XNOR2_X1 input_mapping_1_U8 ( .A(input_mapping_1_n20), .B(XxDI[11]), .ZN(
        input_mapping_1_n18) );
  XNOR2_X1 input_mapping_1_U7 ( .A(XxDI[15]), .B(XxDI[12]), .ZN(
        input_mapping_1_n19) );
  XOR2_X1 input_mapping_1_U6 ( .A(XxDI[8]), .B(input_mapping_1_n21), .Z(
        mappedxD_1__1_) );
  XOR2_X1 input_mapping_1_U5 ( .A(XxDI[14]), .B(XxDI[13]), .Z(
        input_mapping_1_n21) );
  XNOR2_X1 input_mapping_1_U4 ( .A(input_mapping_1_n23), .B(
        input_mapping_1_n17), .ZN(mappedxD_1__0_) );
  XNOR2_X1 input_mapping_1_U3 ( .A(XxDI[14]), .B(XxDI[11]), .ZN(
        input_mapping_1_n17) );
  XNOR2_X1 input_mapping_1_U2 ( .A(XxDI[10]), .B(input_mapping_1_n20), .ZN(
        input_mapping_1_n23) );
  XNOR2_X1 input_mapping_1_U1 ( .A(XxDI[8]), .B(XxDI[9]), .ZN(
        input_mapping_1_n20) );
  XOR2_X1 square_scaler_gf24_1_U3 ( .A(Y0xorY12xD[4]), .B(Y0xorY1xD[4]), .Z(
        Y0xorY12xD[7]) );
  XOR2_X1 square_scaler_gf24_1_U2 ( .A(Y0xorY1xD[3]), .B(Y0xorY1xD[5]), .Z(
        Y0xorY12xD[6]) );
  XOR2_X1 square_scaler_gf24_1_U1 ( .A(Y0xorY12xD[4]), .B(Y0xorY1xD[3]), .Z(
        Y0xorY12xD[5]) );
  XOR2_X1 output_mapping_1_U11 ( .A(InvUnmappedxD[11]), .B(InvUnmappedxD[15]), 
        .Z(QxDO[14]) );
  XNOR2_X1 output_mapping_1_U10 ( .A(QxDO[12]), .B(output_mapping_1_n9), .ZN(
        QxDO[11]) );
  XOR2_X1 output_mapping_1_U9 ( .A(QxDO[15]), .B(InvUnmappedxD[15]), .Z(
        QxDO[12]) );
  XNOR2_X1 output_mapping_1_U8 ( .A(output_mapping_1_n8), .B(QxDO[13]), .ZN(
        QxDO[10]) );
  XNOR2_X1 output_mapping_1_U7 ( .A(QxDO[15]), .B(InvUnmappedxD[10]), .ZN(
        output_mapping_1_n8) );
  XOR2_X1 output_mapping_1_U6 ( .A(InvUnmappedxD[14]), .B(InvUnmappedxD[8]), 
        .Z(QxDO[13]) );
  XOR2_X1 output_mapping_1_U5 ( .A(InvUnmappedxD[11]), .B(InvUnmappedxD[13]), 
        .Z(QxDO[15]) );
  XNOR2_X1 output_mapping_1_U4 ( .A(output_mapping_1_n7), .B(InvUnmappedxD[9]), 
        .ZN(QxDO[9]) );
  XNOR2_X1 output_mapping_1_U3 ( .A(InvUnmappedxD[13]), .B(InvUnmappedxD[12]), 
        .ZN(output_mapping_1_n7) );
  XNOR2_X1 output_mapping_1_U2 ( .A(InvUnmappedxD[9]), .B(output_mapping_1_n9), 
        .ZN(QxDO[8]) );
  XNOR2_X1 output_mapping_1_U1 ( .A(InvUnmappedxD[14]), .B(InvUnmappedxD[12]), 
        .ZN(output_mapping_1_n9) );
  XNOR2_X1 input_mapping_0_U14 ( .A(input_mapping_0_n23), .B(
        input_mapping_0_n22), .ZN(mappedxD_0__7_) );
  XOR2_X1 input_mapping_0_U13 ( .A(XxDI[4]), .B(mappedxD_0__1_), .Z(
        mappedxD_0__6_) );
  XNOR2_X1 input_mapping_0_U12 ( .A(input_mapping_0_n21), .B(
        input_mapping_0_n20), .ZN(mappedxD_0__5_) );
  XNOR2_X1 input_mapping_0_U11 ( .A(XxDI[0]), .B(input_mapping_0_n22), .ZN(
        mappedxD_0__4_) );
  XNOR2_X1 input_mapping_0_U10 ( .A(XxDI[7]), .B(input_mapping_0_n21), .ZN(
        input_mapping_0_n22) );
  XNOR2_X1 input_mapping_0_U9 ( .A(input_mapping_0_n19), .B(
        input_mapping_0_n18), .ZN(mappedxD_0__3_) );
  XNOR2_X1 input_mapping_0_U8 ( .A(input_mapping_0_n20), .B(XxDI[3]), .ZN(
        input_mapping_0_n18) );
  XNOR2_X1 input_mapping_0_U7 ( .A(XxDI[7]), .B(XxDI[4]), .ZN(
        input_mapping_0_n19) );
  XOR2_X1 input_mapping_0_U6 ( .A(XxDI[0]), .B(input_mapping_0_n21), .Z(
        mappedxD_0__1_) );
  XOR2_X1 input_mapping_0_U5 ( .A(XxDI[6]), .B(XxDI[5]), .Z(
        input_mapping_0_n21) );
  XNOR2_X1 input_mapping_0_U4 ( .A(input_mapping_0_n23), .B(
        input_mapping_0_n17), .ZN(mappedxD_0__0_) );
  XNOR2_X1 input_mapping_0_U3 ( .A(XxDI[6]), .B(XxDI[3]), .ZN(
        input_mapping_0_n17) );
  XNOR2_X1 input_mapping_0_U2 ( .A(XxDI[2]), .B(input_mapping_0_n20), .ZN(
        input_mapping_0_n23) );
  XNOR2_X1 input_mapping_0_U1 ( .A(XxDI[0]), .B(XxDI[1]), .ZN(
        input_mapping_0_n20) );
  XOR2_X1 square_scaler_gf24_0_U3 ( .A(Y0xorY12xD[0]), .B(Y0xorY1xD[1]), .Z(
        Y0xorY12xD[3]) );
  XOR2_X1 square_scaler_gf24_0_U2 ( .A(Y0xorY1xD[0]), .B(Y0xorY1xD[2]), .Z(
        Y0xorY12xD[2]) );
  XOR2_X1 square_scaler_gf24_0_U1 ( .A(Y0xorY12xD[0]), .B(Y0xorY1xD[0]), .Z(
        Y0xorY12xD[1]) );
  XOR2_X1 output_mapping_0_U11 ( .A(InvUnmappedxD[3]), .B(InvUnmappedxD[7]), 
        .Z(InvMappedxD_0__6_) );
  XNOR2_X1 output_mapping_0_U10 ( .A(QxDO[4]), .B(output_mapping_0_n9), .ZN(
        QxDO[3]) );
  XOR2_X1 output_mapping_0_U9 ( .A(QxDO[7]), .B(InvUnmappedxD[7]), .Z(QxDO[4])
         );
  XNOR2_X1 output_mapping_0_U8 ( .A(output_mapping_0_n8), .B(InvMappedxD_0__5_), .ZN(QxDO[2]) );
  XNOR2_X1 output_mapping_0_U7 ( .A(QxDO[7]), .B(InvUnmappedxD[2]), .ZN(
        output_mapping_0_n8) );
  XOR2_X1 output_mapping_0_U6 ( .A(InvUnmappedxD[6]), .B(InvUnmappedxD[0]), 
        .Z(InvMappedxD_0__5_) );
  XOR2_X1 output_mapping_0_U5 ( .A(InvUnmappedxD[3]), .B(InvUnmappedxD[5]), 
        .Z(QxDO[7]) );
  XNOR2_X1 output_mapping_0_U4 ( .A(output_mapping_0_n7), .B(InvUnmappedxD[1]), 
        .ZN(InvMappedxD_0__1_) );
  XNOR2_X1 output_mapping_0_U3 ( .A(InvUnmappedxD[5]), .B(InvUnmappedxD[4]), 
        .ZN(output_mapping_0_n7) );
  XNOR2_X1 output_mapping_0_U2 ( .A(InvUnmappedxD[1]), .B(output_mapping_0_n9), 
        .ZN(InvMappedxD_0__0_) );
  XNOR2_X1 output_mapping_0_U1 ( .A(InvUnmappedxD[6]), .B(InvUnmappedxD[4]), 
        .ZN(output_mapping_0_n9) );
  XNOR2_X1 mul_y0y1_U50 ( .A(mul_y0y1_n13), .B(mul_y0y1_n12), .ZN(
        Y0mulY1xD[11]) );
  XOR2_X1 mul_y0y1_U49 ( .A(mul_y0y1_n15), .B(mul_y0y1_n14), .Z(mul_y0y1_n12)
         );
  XNOR2_X1 mul_y0y1_U48 ( .A(mul_y0y1_n16), .B(mul_y0y1_n11), .ZN(
        Y0mulY1xD[10]) );
  XOR2_X1 mul_y0y1_U47 ( .A(mul_y0y1_n18), .B(mul_y0y1_n17), .Z(mul_y0y1_n11)
         );
  XNOR2_X1 mul_y0y1_U46 ( .A(mul_y0y1_n19), .B(mul_y0y1_n10), .ZN(Y0mulY1xD[9]) );
  XOR2_X1 mul_y0y1_U45 ( .A(mul_y0y1_n21), .B(mul_y0y1_n20), .Z(mul_y0y1_n10)
         );
  XNOR2_X1 mul_y0y1_U44 ( .A(mul_y0y1_n22), .B(mul_y0y1_n9), .ZN(Y0mulY1xD[8])
         );
  XOR2_X1 mul_y0y1_U43 ( .A(mul_y0y1_n24), .B(mul_y0y1_n23), .Z(mul_y0y1_n9)
         );
  XNOR2_X1 mul_y0y1_U42 ( .A(mul_y0y1_n25), .B(mul_y0y1_n8), .ZN(Y0mulY1xD[7])
         );
  XOR2_X1 mul_y0y1_U41 ( .A(mul_y0y1_n27), .B(mul_y0y1_n26), .Z(mul_y0y1_n8)
         );
  XNOR2_X1 mul_y0y1_U40 ( .A(mul_y0y1_n28), .B(mul_y0y1_n7), .ZN(Y0mulY1xD[6])
         );
  XOR2_X1 mul_y0y1_U39 ( .A(mul_y0y1_n30), .B(mul_y0y1_n29), .Z(mul_y0y1_n7)
         );
  XNOR2_X1 mul_y0y1_U38 ( .A(mul_y0y1_n31), .B(mul_y0y1_n6), .ZN(Y0mulY1xD[5])
         );
  XOR2_X1 mul_y0y1_U37 ( .A(mul_y0y1_n33), .B(mul_y0y1_n32), .Z(mul_y0y1_n6)
         );
  XNOR2_X1 mul_y0y1_U36 ( .A(mul_y0y1_n34), .B(mul_y0y1_n5), .ZN(Y0mulY1xD[4])
         );
  XOR2_X1 mul_y0y1_U35 ( .A(mul_y0y1_n36), .B(mul_y0y1_n35), .Z(mul_y0y1_n5)
         );
  XNOR2_X1 mul_y0y1_U34 ( .A(mul_y0y1_n37), .B(mul_y0y1_n4), .ZN(Y0mulY1xD[3])
         );
  XOR2_X1 mul_y0y1_U33 ( .A(mul_y0y1_n39), .B(mul_y0y1_n38), .Z(mul_y0y1_n4)
         );
  XNOR2_X1 mul_y0y1_U32 ( .A(mul_y0y1_n40), .B(mul_y0y1_n3), .ZN(Y0mulY1xD[2])
         );
  XOR2_X1 mul_y0y1_U31 ( .A(mul_y0y1_n42), .B(mul_y0y1_n41), .Z(mul_y0y1_n3)
         );
  XNOR2_X1 mul_y0y1_U30 ( .A(mul_y0y1_n43), .B(mul_y0y1_n2), .ZN(Y0mulY1xD[1])
         );
  XOR2_X1 mul_y0y1_U29 ( .A(mul_y0y1_n45), .B(mul_y0y1_n44), .Z(mul_y0y1_n2)
         );
  XNOR2_X1 mul_y0y1_U28 ( .A(mul_y0y1_n46), .B(mul_y0y1_n1), .ZN(Y0mulY1xD[0])
         );
  XOR2_X1 mul_y0y1_U27 ( .A(mul_y0y1_n48), .B(mul_y0y1_n47), .Z(mul_y0y1_n1)
         );
  XOR2_X1 mul_y0y1_U26 ( .A(Zmul1xDI[11]), .B(mul_y0y1_Xi_mul_Yj_7__3_), .Z(
        mul_y0y1_FFxDN[31]) );
  XOR2_X1 mul_y0y1_U25 ( .A(Zmul1xDI[10]), .B(mul_y0y1_Xi_mul_Yj_7__2_), .Z(
        mul_y0y1_FFxDN[30]) );
  XOR2_X1 mul_y0y1_U24 ( .A(Zmul1xDI[9]), .B(mul_y0y1_Xi_mul_Yj_7__1_), .Z(
        mul_y0y1_FFxDN[29]) );
  XOR2_X1 mul_y0y1_U23 ( .A(Zmul1xDI[8]), .B(mul_y0y1_Xi_mul_Yj_7__0_), .Z(
        mul_y0y1_FFxDN[28]) );
  XOR2_X1 mul_y0y1_U22 ( .A(Zmul1xDI[7]), .B(mul_y0y1_Xi_mul_Yj_6__3_), .Z(
        mul_y0y1_FFxDN[27]) );
  XOR2_X1 mul_y0y1_U21 ( .A(Zmul1xDI[6]), .B(mul_y0y1_Xi_mul_Yj_6__2_), .Z(
        mul_y0y1_FFxDN[26]) );
  XOR2_X1 mul_y0y1_U20 ( .A(Zmul1xDI[5]), .B(mul_y0y1_Xi_mul_Yj_6__1_), .Z(
        mul_y0y1_FFxDN[25]) );
  XOR2_X1 mul_y0y1_U19 ( .A(Zmul1xDI[4]), .B(mul_y0y1_Xi_mul_Yj_6__0_), .Z(
        mul_y0y1_FFxDN[24]) );
  XOR2_X1 mul_y0y1_U18 ( .A(Zmul1xDI[11]), .B(mul_y0y1_Xi_mul_Yj_5__3_), .Z(
        mul_y0y1_FFxDN[23]) );
  XOR2_X1 mul_y0y1_U17 ( .A(Zmul1xDI[10]), .B(mul_y0y1_Xi_mul_Yj_5__2_), .Z(
        mul_y0y1_FFxDN[22]) );
  XOR2_X1 mul_y0y1_U16 ( .A(Zmul1xDI[9]), .B(mul_y0y1_Xi_mul_Yj_5__1_), .Z(
        mul_y0y1_FFxDN[21]) );
  XOR2_X1 mul_y0y1_U15 ( .A(Zmul1xDI[8]), .B(mul_y0y1_Xi_mul_Yj_5__0_), .Z(
        mul_y0y1_FFxDN[20]) );
  XOR2_X1 mul_y0y1_U14 ( .A(Zmul1xDI[3]), .B(mul_y0y1_Xi_mul_Yj_3__3_), .Z(
        mul_y0y1_FFxDN[15]) );
  XOR2_X1 mul_y0y1_U13 ( .A(Zmul1xDI[2]), .B(mul_y0y1_Xi_mul_Yj_3__2_), .Z(
        mul_y0y1_FFxDN[14]) );
  XOR2_X1 mul_y0y1_U12 ( .A(Zmul1xDI[1]), .B(mul_y0y1_Xi_mul_Yj_3__1_), .Z(
        mul_y0y1_FFxDN[13]) );
  XOR2_X1 mul_y0y1_U11 ( .A(Zmul1xDI[0]), .B(mul_y0y1_Xi_mul_Yj_3__0_), .Z(
        mul_y0y1_FFxDN[12]) );
  XOR2_X1 mul_y0y1_U10 ( .A(Zmul1xDI[7]), .B(mul_y0y1_Xi_mul_Yj_2__3_), .Z(
        mul_y0y1_FFxDN[11]) );
  XOR2_X1 mul_y0y1_U9 ( .A(Zmul1xDI[6]), .B(mul_y0y1_Xi_mul_Yj_2__2_), .Z(
        mul_y0y1_FFxDN[10]) );
  XOR2_X1 mul_y0y1_U8 ( .A(Zmul1xDI[5]), .B(mul_y0y1_Xi_mul_Yj_2__1_), .Z(
        mul_y0y1_FFxDN[9]) );
  XOR2_X1 mul_y0y1_U7 ( .A(Zmul1xDI[4]), .B(mul_y0y1_Xi_mul_Yj_2__0_), .Z(
        mul_y0y1_FFxDN[8]) );
  XOR2_X1 mul_y0y1_U6 ( .A(Zmul1xDI[3]), .B(mul_y0y1_Xi_mul_Yj_1__3_), .Z(
        mul_y0y1_FFxDN[7]) );
  XOR2_X1 mul_y0y1_U5 ( .A(Zmul1xDI[2]), .B(mul_y0y1_Xi_mul_Yj_1__2_), .Z(
        mul_y0y1_FFxDN[6]) );
  XOR2_X1 mul_y0y1_U4 ( .A(Zmul1xDI[1]), .B(mul_y0y1_Xi_mul_Yj_1__1_), .Z(
        mul_y0y1_FFxDN[5]) );
  XOR2_X1 mul_y0y1_U3 ( .A(Zmul1xDI[0]), .B(mul_y0y1_Xi_mul_Yj_1__0_), .Z(
        mul_y0y1_FFxDN[4]) );
  DFF_X1 mul_y0y1_FFxDP_reg_1__1_ ( .D(mul_y0y1_FFxDN[5]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n44) );
  DFF_X1 mul_y0y1_FFxDP_reg_1__3_ ( .D(mul_y0y1_FFxDN[7]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n38) );
  DFF_X1 mul_y0y1_FFxDP_reg_2__1_ ( .D(mul_y0y1_FFxDN[9]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n45) );
  DFF_X1 mul_y0y1_FFxDP_reg_2__3_ ( .D(mul_y0y1_FFxDN[11]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n39) );
  DFF_X1 mul_y0y1_FFxDP_reg_3__1_ ( .D(mul_y0y1_FFxDN[13]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n31) );
  DFF_X1 mul_y0y1_FFxDP_reg_3__3_ ( .D(mul_y0y1_FFxDN[15]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n25) );
  DFF_X1 mul_y0y1_FFxDP_reg_5__1_ ( .D(mul_y0y1_FFxDN[21]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n33) );
  DFF_X1 mul_y0y1_FFxDP_reg_5__3_ ( .D(mul_y0y1_FFxDN[23]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n27) );
  DFF_X1 mul_y0y1_FFxDP_reg_6__1_ ( .D(mul_y0y1_FFxDN[25]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n19) );
  DFF_X1 mul_y0y1_FFxDP_reg_6__3_ ( .D(mul_y0y1_FFxDN[27]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n13) );
  DFF_X1 mul_y0y1_FFxDP_reg_7__1_ ( .D(mul_y0y1_FFxDN[29]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n20) );
  DFF_X1 mul_y0y1_FFxDP_reg_7__3_ ( .D(mul_y0y1_FFxDN[31]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n14) );
  DFF_X1 mul_y0y1_FFxDP_reg_1__0_ ( .D(mul_y0y1_FFxDN[4]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n47) );
  DFF_X1 mul_y0y1_FFxDP_reg_1__2_ ( .D(mul_y0y1_FFxDN[6]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n41) );
  DFF_X1 mul_y0y1_FFxDP_reg_2__0_ ( .D(mul_y0y1_FFxDN[8]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n48) );
  DFF_X1 mul_y0y1_FFxDP_reg_2__2_ ( .D(mul_y0y1_FFxDN[10]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n42) );
  DFF_X1 mul_y0y1_FFxDP_reg_3__0_ ( .D(mul_y0y1_FFxDN[12]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n34) );
  DFF_X1 mul_y0y1_FFxDP_reg_3__2_ ( .D(mul_y0y1_FFxDN[14]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n28) );
  DFF_X1 mul_y0y1_FFxDP_reg_5__0_ ( .D(mul_y0y1_FFxDN[20]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n36) );
  DFF_X1 mul_y0y1_FFxDP_reg_5__2_ ( .D(mul_y0y1_FFxDN[22]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n30) );
  DFF_X1 mul_y0y1_FFxDP_reg_6__0_ ( .D(mul_y0y1_FFxDN[24]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n22) );
  DFF_X1 mul_y0y1_FFxDP_reg_6__2_ ( .D(mul_y0y1_FFxDN[26]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n16) );
  DFF_X1 mul_y0y1_FFxDP_reg_7__0_ ( .D(mul_y0y1_FFxDN[28]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n23) );
  DFF_X1 mul_y0y1_FFxDP_reg_7__2_ ( .D(mul_y0y1_FFxDN[30]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n17) );
  DFF_X1 mul_y0y1_FFxDP_reg_0__3_ ( .D(mul_y0y1_FFxDN[3]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n37) );
  DFF_X1 mul_y0y1_FFxDP_reg_4__3_ ( .D(mul_y0y1_FFxDN[19]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n26) );
  DFF_X1 mul_y0y1_FFxDP_reg_8__3_ ( .D(mul_y0y1_FFxDN[35]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n15) );
  DFF_X1 mul_y0y1_FFxDP_reg_0__1_ ( .D(mul_y0y1_FFxDN[1]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n43) );
  DFF_X1 mul_y0y1_FFxDP_reg_4__1_ ( .D(mul_y0y1_FFxDN[17]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n32) );
  DFF_X1 mul_y0y1_FFxDP_reg_8__1_ ( .D(mul_y0y1_FFxDN[33]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n21) );
  DFF_X1 mul_y0y1_FFxDP_reg_0__2_ ( .D(mul_y0y1_FFxDN[2]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n40) );
  DFF_X1 mul_y0y1_FFxDP_reg_4__2_ ( .D(mul_y0y1_FFxDN[18]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n29) );
  DFF_X1 mul_y0y1_FFxDP_reg_8__2_ ( .D(mul_y0y1_FFxDN[34]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n18) );
  DFF_X1 mul_y0y1_FFxDP_reg_0__0_ ( .D(mul_y0y1_FFxDN[0]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n46) );
  DFF_X1 mul_y0y1_FFxDP_reg_4__0_ ( .D(mul_y0y1_FFxDN[16]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n35) );
  DFF_X1 mul_y0y1_FFxDP_reg_8__0_ ( .D(mul_y0y1_FFxDN[32]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n24) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U29 ( .A(mul_y0y1_gf4_mul_2_2_n77), .B(
        mul_y0y1_gf4_mul_2_2_n76), .ZN(mul_y0y1_FFxDN[35]) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U28 ( .A1(Y1xD[11]), .A2(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_2_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U27 ( .A(mul_y0y1_gf4_mul_2_2_n75), .B(
        mul_y0y1_gf4_mul_2_2_n74), .Z(mul_y0y1_gf4_mul_2_2_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U26 ( .A(mul_y0y1_gf4_mul_2_2_n73), .B(
        mul_y0y1_gf4_mul_2_2_n72), .ZN(mul_y0y1_FFxDN[34]) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U25 ( .A1(Y1xD[10]), .A2(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_2_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U24 ( .A(mul_y0y1_gf4_mul_2_2_n74), .B(
        mul_y0y1_gf4_mul_2_2_n71), .Z(mul_y0y1_gf4_mul_2_2_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_2_2_U23 ( .A1(mul_y0y1_gf4_mul_2_2_n70), .A2(
        mul_y0y1_gf4_mul_2_2_n69), .ZN(mul_y0y1_gf4_mul_2_2_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U22 ( .A(Y1xD[10]), .B(Y1xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_2_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U21 ( .A(Y0xD[10]), .B(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_2_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U20 ( .A(mul_y0y1_gf4_mul_2_2_n68), .B(
        mul_y0y1_gf4_mul_2_2_n67), .ZN(mul_y0y1_FFxDN[33]) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U19 ( .A1(Y1xD[9]), .A2(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_2_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U18 ( .A(mul_y0y1_gf4_mul_2_2_n75), .B(
        mul_y0y1_gf4_mul_2_2_n66), .Z(mul_y0y1_gf4_mul_2_2_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U17 ( .A(mul_y0y1_gf4_mul_2_2_n65), .B(
        mul_y0y1_gf4_mul_2_2_n64), .ZN(mul_y0y1_gf4_mul_2_2_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U16 ( .A1(mul_y0y1_gf4_mul_2_2_n63), .A2(
        mul_y0y1_gf4_mul_2_2_n62), .ZN(mul_y0y1_gf4_mul_2_2_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U15 ( .A(mul_y0y1_gf4_mul_2_2_n61), .B(
        mul_y0y1_gf4_mul_2_2_n60), .ZN(mul_y0y1_gf4_mul_2_2_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U14 ( .A(mul_y0y1_gf4_mul_2_2_n59), .B(
        mul_y0y1_gf4_mul_2_2_n58), .ZN(mul_y0y1_gf4_mul_2_2_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U13 ( .A(mul_y0y1_gf4_mul_2_2_n57), .B(
        mul_y0y1_gf4_mul_2_2_n56), .ZN(mul_y0y1_FFxDN[32]) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U12 ( .A1(Y1xD[8]), .A2(Y0xD[8]), .ZN(
        mul_y0y1_gf4_mul_2_2_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U11 ( .A(mul_y0y1_gf4_mul_2_2_n66), .B(
        mul_y0y1_gf4_mul_2_2_n71), .Z(mul_y0y1_gf4_mul_2_2_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U10 ( .A(mul_y0y1_gf4_mul_2_2_n55), .B(
        mul_y0y1_gf4_mul_2_2_n65), .ZN(mul_y0y1_gf4_mul_2_2_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_2_2_U9 ( .A1(mul_y0y1_gf4_mul_2_2_n61), .A2(
        mul_y0y1_gf4_mul_2_2_n59), .ZN(mul_y0y1_gf4_mul_2_2_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U8 ( .A(Y1xD[8]), .B(Y1xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_2_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U7 ( .A(Y0xD[8]), .B(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_2_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U6 ( .A1(mul_y0y1_gf4_mul_2_2_n58), .A2(
        mul_y0y1_gf4_mul_2_2_n60), .ZN(mul_y0y1_gf4_mul_2_2_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U5 ( .A(Y0xD[9]), .B(Y0xD[11]), .Z(
        mul_y0y1_gf4_mul_2_2_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U4 ( .A(Y1xD[9]), .B(Y1xD[11]), .Z(
        mul_y0y1_gf4_mul_2_2_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_2_2_U3 ( .A1(mul_y0y1_gf4_mul_2_2_n54), .A2(
        mul_y0y1_gf4_mul_2_2_n53), .ZN(mul_y0y1_gf4_mul_2_2_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U2 ( .A(Y1xD[8]), .B(Y1xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_2_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U1 ( .A(Y0xD[8]), .B(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_2_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U29 ( .A(mul_y0y1_gf4_mul_2_1_n77), .B(
        mul_y0y1_gf4_mul_2_1_n76), .ZN(mul_y0y1_Xi_mul_Yj_7__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U28 ( .A1(Y1xD[11]), .A2(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_2_1_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U27 ( .A(mul_y0y1_gf4_mul_2_1_n75), .B(
        mul_y0y1_gf4_mul_2_1_n74), .Z(mul_y0y1_gf4_mul_2_1_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U26 ( .A(mul_y0y1_gf4_mul_2_1_n73), .B(
        mul_y0y1_gf4_mul_2_1_n72), .ZN(mul_y0y1_Xi_mul_Yj_7__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U25 ( .A1(Y1xD[10]), .A2(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_2_1_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U24 ( .A(mul_y0y1_gf4_mul_2_1_n74), .B(
        mul_y0y1_gf4_mul_2_1_n71), .Z(mul_y0y1_gf4_mul_2_1_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_2_1_U23 ( .A1(mul_y0y1_gf4_mul_2_1_n70), .A2(
        mul_y0y1_gf4_mul_2_1_n69), .ZN(mul_y0y1_gf4_mul_2_1_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U22 ( .A(Y1xD[10]), .B(Y1xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_1_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U21 ( .A(Y0xD[6]), .B(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_2_1_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U20 ( .A(mul_y0y1_gf4_mul_2_1_n68), .B(
        mul_y0y1_gf4_mul_2_1_n67), .ZN(mul_y0y1_Xi_mul_Yj_7__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U19 ( .A1(Y1xD[9]), .A2(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_2_1_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U18 ( .A(mul_y0y1_gf4_mul_2_1_n75), .B(
        mul_y0y1_gf4_mul_2_1_n66), .Z(mul_y0y1_gf4_mul_2_1_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U17 ( .A(mul_y0y1_gf4_mul_2_1_n65), .B(
        mul_y0y1_gf4_mul_2_1_n64), .ZN(mul_y0y1_gf4_mul_2_1_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U16 ( .A1(mul_y0y1_gf4_mul_2_1_n63), .A2(
        mul_y0y1_gf4_mul_2_1_n62), .ZN(mul_y0y1_gf4_mul_2_1_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U15 ( .A(mul_y0y1_gf4_mul_2_1_n61), .B(
        mul_y0y1_gf4_mul_2_1_n60), .ZN(mul_y0y1_gf4_mul_2_1_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U14 ( .A(mul_y0y1_gf4_mul_2_1_n59), .B(
        mul_y0y1_gf4_mul_2_1_n58), .ZN(mul_y0y1_gf4_mul_2_1_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U13 ( .A(mul_y0y1_gf4_mul_2_1_n57), .B(
        mul_y0y1_gf4_mul_2_1_n56), .ZN(mul_y0y1_Xi_mul_Yj_7__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U12 ( .A1(Y1xD[8]), .A2(Y0xD[4]), .ZN(
        mul_y0y1_gf4_mul_2_1_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U11 ( .A(mul_y0y1_gf4_mul_2_1_n66), .B(
        mul_y0y1_gf4_mul_2_1_n71), .Z(mul_y0y1_gf4_mul_2_1_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U10 ( .A(mul_y0y1_gf4_mul_2_1_n55), .B(
        mul_y0y1_gf4_mul_2_1_n65), .ZN(mul_y0y1_gf4_mul_2_1_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_2_1_U9 ( .A1(mul_y0y1_gf4_mul_2_1_n61), .A2(
        mul_y0y1_gf4_mul_2_1_n59), .ZN(mul_y0y1_gf4_mul_2_1_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U8 ( .A(Y1xD[8]), .B(Y1xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_1_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U7 ( .A(Y0xD[4]), .B(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_2_1_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U6 ( .A1(mul_y0y1_gf4_mul_2_1_n58), .A2(
        mul_y0y1_gf4_mul_2_1_n60), .ZN(mul_y0y1_gf4_mul_2_1_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U5 ( .A(Y0xD[5]), .B(Y0xD[7]), .Z(
        mul_y0y1_gf4_mul_2_1_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U4 ( .A(Y1xD[9]), .B(Y1xD[11]), .Z(
        mul_y0y1_gf4_mul_2_1_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_2_1_U3 ( .A1(mul_y0y1_gf4_mul_2_1_n54), .A2(
        mul_y0y1_gf4_mul_2_1_n53), .ZN(mul_y0y1_gf4_mul_2_1_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U2 ( .A(Y1xD[8]), .B(Y1xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_1_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U1 ( .A(Y0xD[4]), .B(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_2_1_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U29 ( .A(mul_y0y1_gf4_mul_2_0_n77), .B(
        mul_y0y1_gf4_mul_2_0_n76), .ZN(mul_y0y1_Xi_mul_Yj_6__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U28 ( .A1(Y1xD[11]), .A2(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_2_0_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U27 ( .A(mul_y0y1_gf4_mul_2_0_n75), .B(
        mul_y0y1_gf4_mul_2_0_n74), .Z(mul_y0y1_gf4_mul_2_0_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U26 ( .A(mul_y0y1_gf4_mul_2_0_n73), .B(
        mul_y0y1_gf4_mul_2_0_n72), .ZN(mul_y0y1_Xi_mul_Yj_6__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U25 ( .A1(Y1xD[10]), .A2(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_2_0_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U24 ( .A(mul_y0y1_gf4_mul_2_0_n74), .B(
        mul_y0y1_gf4_mul_2_0_n71), .Z(mul_y0y1_gf4_mul_2_0_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_2_0_U23 ( .A1(mul_y0y1_gf4_mul_2_0_n70), .A2(
        mul_y0y1_gf4_mul_2_0_n69), .ZN(mul_y0y1_gf4_mul_2_0_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U22 ( .A(Y1xD[10]), .B(Y1xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_0_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U21 ( .A(Y0xD[2]), .B(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_2_0_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U20 ( .A(mul_y0y1_gf4_mul_2_0_n68), .B(
        mul_y0y1_gf4_mul_2_0_n67), .ZN(mul_y0y1_Xi_mul_Yj_6__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U19 ( .A1(Y1xD[9]), .A2(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_2_0_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U18 ( .A(mul_y0y1_gf4_mul_2_0_n75), .B(
        mul_y0y1_gf4_mul_2_0_n66), .Z(mul_y0y1_gf4_mul_2_0_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U17 ( .A(mul_y0y1_gf4_mul_2_0_n65), .B(
        mul_y0y1_gf4_mul_2_0_n64), .ZN(mul_y0y1_gf4_mul_2_0_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U16 ( .A1(mul_y0y1_gf4_mul_2_0_n63), .A2(
        mul_y0y1_gf4_mul_2_0_n62), .ZN(mul_y0y1_gf4_mul_2_0_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U15 ( .A(mul_y0y1_gf4_mul_2_0_n61), .B(
        mul_y0y1_gf4_mul_2_0_n60), .ZN(mul_y0y1_gf4_mul_2_0_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U14 ( .A(mul_y0y1_gf4_mul_2_0_n59), .B(
        mul_y0y1_gf4_mul_2_0_n58), .ZN(mul_y0y1_gf4_mul_2_0_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U13 ( .A(mul_y0y1_gf4_mul_2_0_n57), .B(
        mul_y0y1_gf4_mul_2_0_n56), .ZN(mul_y0y1_Xi_mul_Yj_6__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U12 ( .A1(Y1xD[8]), .A2(Y0xD[0]), .ZN(
        mul_y0y1_gf4_mul_2_0_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U11 ( .A(mul_y0y1_gf4_mul_2_0_n66), .B(
        mul_y0y1_gf4_mul_2_0_n71), .Z(mul_y0y1_gf4_mul_2_0_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U10 ( .A(mul_y0y1_gf4_mul_2_0_n55), .B(
        mul_y0y1_gf4_mul_2_0_n65), .ZN(mul_y0y1_gf4_mul_2_0_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_2_0_U9 ( .A1(mul_y0y1_gf4_mul_2_0_n61), .A2(
        mul_y0y1_gf4_mul_2_0_n59), .ZN(mul_y0y1_gf4_mul_2_0_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U8 ( .A(Y1xD[8]), .B(Y1xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_0_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U7 ( .A(Y0xD[0]), .B(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_2_0_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U6 ( .A1(mul_y0y1_gf4_mul_2_0_n58), .A2(
        mul_y0y1_gf4_mul_2_0_n60), .ZN(mul_y0y1_gf4_mul_2_0_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U5 ( .A(Y0xD[1]), .B(Y0xD[3]), .Z(
        mul_y0y1_gf4_mul_2_0_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U4 ( .A(Y1xD[9]), .B(Y1xD[11]), .Z(
        mul_y0y1_gf4_mul_2_0_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_2_0_U3 ( .A1(mul_y0y1_gf4_mul_2_0_n54), .A2(
        mul_y0y1_gf4_mul_2_0_n53), .ZN(mul_y0y1_gf4_mul_2_0_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U2 ( .A(Y1xD[8]), .B(Y1xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_0_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U1 ( .A(Y0xD[0]), .B(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_2_0_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U29 ( .A(mul_y0y1_gf4_mul_1_2_n77), .B(
        mul_y0y1_gf4_mul_1_2_n76), .ZN(mul_y0y1_Xi_mul_Yj_5__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U28 ( .A1(Y1xD[7]), .A2(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_1_2_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U27 ( .A(mul_y0y1_gf4_mul_1_2_n75), .B(
        mul_y0y1_gf4_mul_1_2_n74), .Z(mul_y0y1_gf4_mul_1_2_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U26 ( .A(mul_y0y1_gf4_mul_1_2_n73), .B(
        mul_y0y1_gf4_mul_1_2_n72), .ZN(mul_y0y1_Xi_mul_Yj_5__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U25 ( .A1(Y1xD[6]), .A2(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_1_2_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U24 ( .A(mul_y0y1_gf4_mul_1_2_n74), .B(
        mul_y0y1_gf4_mul_1_2_n71), .Z(mul_y0y1_gf4_mul_1_2_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_1_2_U23 ( .A1(mul_y0y1_gf4_mul_1_2_n70), .A2(
        mul_y0y1_gf4_mul_1_2_n69), .ZN(mul_y0y1_gf4_mul_1_2_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U22 ( .A(Y1xD[6]), .B(Y1xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_2_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U21 ( .A(Y0xD[10]), .B(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_1_2_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U20 ( .A(mul_y0y1_gf4_mul_1_2_n68), .B(
        mul_y0y1_gf4_mul_1_2_n67), .ZN(mul_y0y1_Xi_mul_Yj_5__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U19 ( .A1(Y1xD[5]), .A2(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_1_2_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U18 ( .A(mul_y0y1_gf4_mul_1_2_n75), .B(
        mul_y0y1_gf4_mul_1_2_n66), .Z(mul_y0y1_gf4_mul_1_2_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U17 ( .A(mul_y0y1_gf4_mul_1_2_n65), .B(
        mul_y0y1_gf4_mul_1_2_n64), .ZN(mul_y0y1_gf4_mul_1_2_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U16 ( .A1(mul_y0y1_gf4_mul_1_2_n63), .A2(
        mul_y0y1_gf4_mul_1_2_n62), .ZN(mul_y0y1_gf4_mul_1_2_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U15 ( .A(mul_y0y1_gf4_mul_1_2_n61), .B(
        mul_y0y1_gf4_mul_1_2_n60), .ZN(mul_y0y1_gf4_mul_1_2_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U14 ( .A(mul_y0y1_gf4_mul_1_2_n59), .B(
        mul_y0y1_gf4_mul_1_2_n58), .ZN(mul_y0y1_gf4_mul_1_2_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U13 ( .A(mul_y0y1_gf4_mul_1_2_n57), .B(
        mul_y0y1_gf4_mul_1_2_n56), .ZN(mul_y0y1_Xi_mul_Yj_5__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U12 ( .A1(Y1xD[4]), .A2(Y0xD[8]), .ZN(
        mul_y0y1_gf4_mul_1_2_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U11 ( .A(mul_y0y1_gf4_mul_1_2_n66), .B(
        mul_y0y1_gf4_mul_1_2_n71), .Z(mul_y0y1_gf4_mul_1_2_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U10 ( .A(mul_y0y1_gf4_mul_1_2_n55), .B(
        mul_y0y1_gf4_mul_1_2_n65), .ZN(mul_y0y1_gf4_mul_1_2_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_1_2_U9 ( .A1(mul_y0y1_gf4_mul_1_2_n61), .A2(
        mul_y0y1_gf4_mul_1_2_n59), .ZN(mul_y0y1_gf4_mul_1_2_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U8 ( .A(Y1xD[4]), .B(Y1xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_2_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U7 ( .A(Y0xD[8]), .B(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_1_2_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U6 ( .A1(mul_y0y1_gf4_mul_1_2_n58), .A2(
        mul_y0y1_gf4_mul_1_2_n60), .ZN(mul_y0y1_gf4_mul_1_2_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U5 ( .A(Y0xD[9]), .B(Y0xD[11]), .Z(
        mul_y0y1_gf4_mul_1_2_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U4 ( .A(Y1xD[5]), .B(Y1xD[7]), .Z(
        mul_y0y1_gf4_mul_1_2_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_1_2_U3 ( .A1(mul_y0y1_gf4_mul_1_2_n54), .A2(
        mul_y0y1_gf4_mul_1_2_n53), .ZN(mul_y0y1_gf4_mul_1_2_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U2 ( .A(Y1xD[4]), .B(Y1xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_2_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U1 ( .A(Y0xD[8]), .B(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_1_2_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U29 ( .A(mul_y0y1_gf4_mul_1_1_n77), .B(
        mul_y0y1_gf4_mul_1_1_n76), .ZN(mul_y0y1_FFxDN[19]) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U28 ( .A1(Y1xD[7]), .A2(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_1_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U27 ( .A(mul_y0y1_gf4_mul_1_1_n75), .B(
        mul_y0y1_gf4_mul_1_1_n74), .Z(mul_y0y1_gf4_mul_1_1_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U26 ( .A(mul_y0y1_gf4_mul_1_1_n73), .B(
        mul_y0y1_gf4_mul_1_1_n72), .ZN(mul_y0y1_FFxDN[18]) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U25 ( .A1(Y1xD[6]), .A2(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_1_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U24 ( .A(mul_y0y1_gf4_mul_1_1_n74), .B(
        mul_y0y1_gf4_mul_1_1_n71), .Z(mul_y0y1_gf4_mul_1_1_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_1_1_U23 ( .A1(mul_y0y1_gf4_mul_1_1_n70), .A2(
        mul_y0y1_gf4_mul_1_1_n69), .ZN(mul_y0y1_gf4_mul_1_1_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U22 ( .A(Y1xD[6]), .B(Y1xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_1_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U21 ( .A(Y0xD[6]), .B(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_1_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U20 ( .A(mul_y0y1_gf4_mul_1_1_n68), .B(
        mul_y0y1_gf4_mul_1_1_n67), .ZN(mul_y0y1_FFxDN[17]) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U19 ( .A1(Y1xD[5]), .A2(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_1_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U18 ( .A(mul_y0y1_gf4_mul_1_1_n75), .B(
        mul_y0y1_gf4_mul_1_1_n66), .Z(mul_y0y1_gf4_mul_1_1_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U17 ( .A(mul_y0y1_gf4_mul_1_1_n65), .B(
        mul_y0y1_gf4_mul_1_1_n64), .ZN(mul_y0y1_gf4_mul_1_1_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U16 ( .A1(mul_y0y1_gf4_mul_1_1_n63), .A2(
        mul_y0y1_gf4_mul_1_1_n62), .ZN(mul_y0y1_gf4_mul_1_1_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U15 ( .A(mul_y0y1_gf4_mul_1_1_n61), .B(
        mul_y0y1_gf4_mul_1_1_n60), .ZN(mul_y0y1_gf4_mul_1_1_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U14 ( .A(mul_y0y1_gf4_mul_1_1_n59), .B(
        mul_y0y1_gf4_mul_1_1_n58), .ZN(mul_y0y1_gf4_mul_1_1_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U13 ( .A(mul_y0y1_gf4_mul_1_1_n57), .B(
        mul_y0y1_gf4_mul_1_1_n56), .ZN(mul_y0y1_FFxDN[16]) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U12 ( .A1(Y1xD[4]), .A2(Y0xD[4]), .ZN(
        mul_y0y1_gf4_mul_1_1_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U11 ( .A(mul_y0y1_gf4_mul_1_1_n66), .B(
        mul_y0y1_gf4_mul_1_1_n71), .Z(mul_y0y1_gf4_mul_1_1_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U10 ( .A(mul_y0y1_gf4_mul_1_1_n55), .B(
        mul_y0y1_gf4_mul_1_1_n65), .ZN(mul_y0y1_gf4_mul_1_1_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_1_1_U9 ( .A1(mul_y0y1_gf4_mul_1_1_n61), .A2(
        mul_y0y1_gf4_mul_1_1_n59), .ZN(mul_y0y1_gf4_mul_1_1_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U8 ( .A(Y1xD[4]), .B(Y1xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_1_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U7 ( .A(Y0xD[4]), .B(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_1_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U6 ( .A1(mul_y0y1_gf4_mul_1_1_n58), .A2(
        mul_y0y1_gf4_mul_1_1_n60), .ZN(mul_y0y1_gf4_mul_1_1_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U5 ( .A(Y0xD[5]), .B(Y0xD[7]), .Z(
        mul_y0y1_gf4_mul_1_1_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U4 ( .A(Y1xD[5]), .B(Y1xD[7]), .Z(
        mul_y0y1_gf4_mul_1_1_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_1_1_U3 ( .A1(mul_y0y1_gf4_mul_1_1_n54), .A2(
        mul_y0y1_gf4_mul_1_1_n53), .ZN(mul_y0y1_gf4_mul_1_1_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U2 ( .A(Y1xD[4]), .B(Y1xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_1_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U1 ( .A(Y0xD[4]), .B(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_1_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U29 ( .A(mul_y0y1_gf4_mul_1_0_n77), .B(
        mul_y0y1_gf4_mul_1_0_n76), .ZN(mul_y0y1_Xi_mul_Yj_3__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U28 ( .A1(Y1xD[7]), .A2(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_1_0_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U27 ( .A(mul_y0y1_gf4_mul_1_0_n75), .B(
        mul_y0y1_gf4_mul_1_0_n74), .Z(mul_y0y1_gf4_mul_1_0_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U26 ( .A(mul_y0y1_gf4_mul_1_0_n73), .B(
        mul_y0y1_gf4_mul_1_0_n72), .ZN(mul_y0y1_Xi_mul_Yj_3__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U25 ( .A1(Y1xD[6]), .A2(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_1_0_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U24 ( .A(mul_y0y1_gf4_mul_1_0_n74), .B(
        mul_y0y1_gf4_mul_1_0_n71), .Z(mul_y0y1_gf4_mul_1_0_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_1_0_U23 ( .A1(mul_y0y1_gf4_mul_1_0_n70), .A2(
        mul_y0y1_gf4_mul_1_0_n69), .ZN(mul_y0y1_gf4_mul_1_0_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U22 ( .A(Y1xD[6]), .B(Y1xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_0_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U21 ( .A(Y0xD[2]), .B(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_1_0_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U20 ( .A(mul_y0y1_gf4_mul_1_0_n68), .B(
        mul_y0y1_gf4_mul_1_0_n67), .ZN(mul_y0y1_Xi_mul_Yj_3__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U19 ( .A1(Y1xD[5]), .A2(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_1_0_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U18 ( .A(mul_y0y1_gf4_mul_1_0_n75), .B(
        mul_y0y1_gf4_mul_1_0_n66), .Z(mul_y0y1_gf4_mul_1_0_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U17 ( .A(mul_y0y1_gf4_mul_1_0_n65), .B(
        mul_y0y1_gf4_mul_1_0_n64), .ZN(mul_y0y1_gf4_mul_1_0_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U16 ( .A1(mul_y0y1_gf4_mul_1_0_n63), .A2(
        mul_y0y1_gf4_mul_1_0_n62), .ZN(mul_y0y1_gf4_mul_1_0_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U15 ( .A(mul_y0y1_gf4_mul_1_0_n61), .B(
        mul_y0y1_gf4_mul_1_0_n60), .ZN(mul_y0y1_gf4_mul_1_0_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U14 ( .A(mul_y0y1_gf4_mul_1_0_n59), .B(
        mul_y0y1_gf4_mul_1_0_n58), .ZN(mul_y0y1_gf4_mul_1_0_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U13 ( .A(mul_y0y1_gf4_mul_1_0_n57), .B(
        mul_y0y1_gf4_mul_1_0_n56), .ZN(mul_y0y1_Xi_mul_Yj_3__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U12 ( .A1(Y1xD[4]), .A2(Y0xD[0]), .ZN(
        mul_y0y1_gf4_mul_1_0_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U11 ( .A(mul_y0y1_gf4_mul_1_0_n66), .B(
        mul_y0y1_gf4_mul_1_0_n71), .Z(mul_y0y1_gf4_mul_1_0_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U10 ( .A(mul_y0y1_gf4_mul_1_0_n55), .B(
        mul_y0y1_gf4_mul_1_0_n65), .ZN(mul_y0y1_gf4_mul_1_0_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_1_0_U9 ( .A1(mul_y0y1_gf4_mul_1_0_n61), .A2(
        mul_y0y1_gf4_mul_1_0_n59), .ZN(mul_y0y1_gf4_mul_1_0_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U8 ( .A(Y1xD[4]), .B(Y1xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_0_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U7 ( .A(Y0xD[0]), .B(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_1_0_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U6 ( .A1(mul_y0y1_gf4_mul_1_0_n58), .A2(
        mul_y0y1_gf4_mul_1_0_n60), .ZN(mul_y0y1_gf4_mul_1_0_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U5 ( .A(Y0xD[1]), .B(Y0xD[3]), .Z(
        mul_y0y1_gf4_mul_1_0_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U4 ( .A(Y1xD[5]), .B(Y1xD[7]), .Z(
        mul_y0y1_gf4_mul_1_0_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_1_0_U3 ( .A1(mul_y0y1_gf4_mul_1_0_n54), .A2(
        mul_y0y1_gf4_mul_1_0_n53), .ZN(mul_y0y1_gf4_mul_1_0_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U2 ( .A(Y1xD[4]), .B(Y1xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_0_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U1 ( .A(Y0xD[0]), .B(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_1_0_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U29 ( .A(mul_y0y1_gf4_mul_0_2_n77), .B(
        mul_y0y1_gf4_mul_0_2_n76), .ZN(mul_y0y1_Xi_mul_Yj_2__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U28 ( .A1(Y1xD[3]), .A2(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_0_2_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U27 ( .A(mul_y0y1_gf4_mul_0_2_n75), .B(
        mul_y0y1_gf4_mul_0_2_n74), .Z(mul_y0y1_gf4_mul_0_2_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U26 ( .A(mul_y0y1_gf4_mul_0_2_n73), .B(
        mul_y0y1_gf4_mul_0_2_n72), .ZN(mul_y0y1_Xi_mul_Yj_2__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U25 ( .A1(Y1xD[2]), .A2(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_0_2_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U24 ( .A(mul_y0y1_gf4_mul_0_2_n74), .B(
        mul_y0y1_gf4_mul_0_2_n71), .Z(mul_y0y1_gf4_mul_0_2_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_0_2_U23 ( .A1(mul_y0y1_gf4_mul_0_2_n70), .A2(
        mul_y0y1_gf4_mul_0_2_n69), .ZN(mul_y0y1_gf4_mul_0_2_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U22 ( .A(Y1xD[2]), .B(Y1xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_2_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U21 ( .A(Y0xD[10]), .B(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_0_2_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U20 ( .A(mul_y0y1_gf4_mul_0_2_n68), .B(
        mul_y0y1_gf4_mul_0_2_n67), .ZN(mul_y0y1_Xi_mul_Yj_2__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U19 ( .A1(Y1xD[1]), .A2(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_0_2_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U18 ( .A(mul_y0y1_gf4_mul_0_2_n75), .B(
        mul_y0y1_gf4_mul_0_2_n66), .Z(mul_y0y1_gf4_mul_0_2_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U17 ( .A(mul_y0y1_gf4_mul_0_2_n65), .B(
        mul_y0y1_gf4_mul_0_2_n64), .ZN(mul_y0y1_gf4_mul_0_2_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U16 ( .A1(mul_y0y1_gf4_mul_0_2_n63), .A2(
        mul_y0y1_gf4_mul_0_2_n62), .ZN(mul_y0y1_gf4_mul_0_2_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U15 ( .A(mul_y0y1_gf4_mul_0_2_n61), .B(
        mul_y0y1_gf4_mul_0_2_n60), .ZN(mul_y0y1_gf4_mul_0_2_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U14 ( .A(mul_y0y1_gf4_mul_0_2_n59), .B(
        mul_y0y1_gf4_mul_0_2_n58), .ZN(mul_y0y1_gf4_mul_0_2_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U13 ( .A(mul_y0y1_gf4_mul_0_2_n57), .B(
        mul_y0y1_gf4_mul_0_2_n56), .ZN(mul_y0y1_Xi_mul_Yj_2__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U12 ( .A1(Y1xD[0]), .A2(Y0xD[8]), .ZN(
        mul_y0y1_gf4_mul_0_2_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U11 ( .A(mul_y0y1_gf4_mul_0_2_n66), .B(
        mul_y0y1_gf4_mul_0_2_n71), .Z(mul_y0y1_gf4_mul_0_2_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U10 ( .A(mul_y0y1_gf4_mul_0_2_n55), .B(
        mul_y0y1_gf4_mul_0_2_n65), .ZN(mul_y0y1_gf4_mul_0_2_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_0_2_U9 ( .A1(mul_y0y1_gf4_mul_0_2_n61), .A2(
        mul_y0y1_gf4_mul_0_2_n59), .ZN(mul_y0y1_gf4_mul_0_2_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U8 ( .A(Y1xD[0]), .B(Y1xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_2_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U7 ( .A(Y0xD[8]), .B(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_0_2_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U6 ( .A1(mul_y0y1_gf4_mul_0_2_n58), .A2(
        mul_y0y1_gf4_mul_0_2_n60), .ZN(mul_y0y1_gf4_mul_0_2_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U5 ( .A(Y0xD[9]), .B(Y0xD[11]), .Z(
        mul_y0y1_gf4_mul_0_2_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U4 ( .A(Y1xD[1]), .B(Y1xD[3]), .Z(
        mul_y0y1_gf4_mul_0_2_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_0_2_U3 ( .A1(mul_y0y1_gf4_mul_0_2_n54), .A2(
        mul_y0y1_gf4_mul_0_2_n53), .ZN(mul_y0y1_gf4_mul_0_2_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U2 ( .A(Y1xD[0]), .B(Y1xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_2_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U1 ( .A(Y0xD[8]), .B(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_0_2_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U29 ( .A(mul_y0y1_gf4_mul_0_1_n77), .B(
        mul_y0y1_gf4_mul_0_1_n76), .ZN(mul_y0y1_Xi_mul_Yj_1__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U28 ( .A1(Y1xD[3]), .A2(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_0_1_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U27 ( .A(mul_y0y1_gf4_mul_0_1_n75), .B(
        mul_y0y1_gf4_mul_0_1_n74), .Z(mul_y0y1_gf4_mul_0_1_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U26 ( .A(mul_y0y1_gf4_mul_0_1_n73), .B(
        mul_y0y1_gf4_mul_0_1_n72), .ZN(mul_y0y1_Xi_mul_Yj_1__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U25 ( .A1(Y1xD[2]), .A2(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_0_1_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U24 ( .A(mul_y0y1_gf4_mul_0_1_n74), .B(
        mul_y0y1_gf4_mul_0_1_n71), .Z(mul_y0y1_gf4_mul_0_1_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_0_1_U23 ( .A1(mul_y0y1_gf4_mul_0_1_n70), .A2(
        mul_y0y1_gf4_mul_0_1_n69), .ZN(mul_y0y1_gf4_mul_0_1_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U22 ( .A(Y1xD[2]), .B(Y1xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_1_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U21 ( .A(Y0xD[6]), .B(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_0_1_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U20 ( .A(mul_y0y1_gf4_mul_0_1_n68), .B(
        mul_y0y1_gf4_mul_0_1_n67), .ZN(mul_y0y1_Xi_mul_Yj_1__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U19 ( .A1(Y1xD[1]), .A2(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_0_1_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U18 ( .A(mul_y0y1_gf4_mul_0_1_n75), .B(
        mul_y0y1_gf4_mul_0_1_n66), .Z(mul_y0y1_gf4_mul_0_1_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U17 ( .A(mul_y0y1_gf4_mul_0_1_n65), .B(
        mul_y0y1_gf4_mul_0_1_n64), .ZN(mul_y0y1_gf4_mul_0_1_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U16 ( .A1(mul_y0y1_gf4_mul_0_1_n63), .A2(
        mul_y0y1_gf4_mul_0_1_n62), .ZN(mul_y0y1_gf4_mul_0_1_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U15 ( .A(mul_y0y1_gf4_mul_0_1_n61), .B(
        mul_y0y1_gf4_mul_0_1_n60), .ZN(mul_y0y1_gf4_mul_0_1_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U14 ( .A(mul_y0y1_gf4_mul_0_1_n59), .B(
        mul_y0y1_gf4_mul_0_1_n58), .ZN(mul_y0y1_gf4_mul_0_1_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U13 ( .A(mul_y0y1_gf4_mul_0_1_n57), .B(
        mul_y0y1_gf4_mul_0_1_n56), .ZN(mul_y0y1_Xi_mul_Yj_1__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U12 ( .A1(Y1xD[0]), .A2(Y0xD[4]), .ZN(
        mul_y0y1_gf4_mul_0_1_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U11 ( .A(mul_y0y1_gf4_mul_0_1_n66), .B(
        mul_y0y1_gf4_mul_0_1_n71), .Z(mul_y0y1_gf4_mul_0_1_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U10 ( .A(mul_y0y1_gf4_mul_0_1_n55), .B(
        mul_y0y1_gf4_mul_0_1_n65), .ZN(mul_y0y1_gf4_mul_0_1_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_0_1_U9 ( .A1(mul_y0y1_gf4_mul_0_1_n61), .A2(
        mul_y0y1_gf4_mul_0_1_n59), .ZN(mul_y0y1_gf4_mul_0_1_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U8 ( .A(Y1xD[0]), .B(Y1xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_1_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U7 ( .A(Y0xD[4]), .B(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_0_1_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U6 ( .A1(mul_y0y1_gf4_mul_0_1_n58), .A2(
        mul_y0y1_gf4_mul_0_1_n60), .ZN(mul_y0y1_gf4_mul_0_1_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U5 ( .A(Y0xD[5]), .B(Y0xD[7]), .Z(
        mul_y0y1_gf4_mul_0_1_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U4 ( .A(Y1xD[1]), .B(Y1xD[3]), .Z(
        mul_y0y1_gf4_mul_0_1_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_0_1_U3 ( .A1(mul_y0y1_gf4_mul_0_1_n54), .A2(
        mul_y0y1_gf4_mul_0_1_n53), .ZN(mul_y0y1_gf4_mul_0_1_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U2 ( .A(Y1xD[0]), .B(Y1xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_1_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U1 ( .A(Y0xD[4]), .B(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_0_1_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U29 ( .A(mul_y0y1_gf4_mul_0_0_n77), .B(
        mul_y0y1_gf4_mul_0_0_n76), .ZN(mul_y0y1_FFxDN[3]) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U28 ( .A1(Y1xD[3]), .A2(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_0_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U27 ( .A(mul_y0y1_gf4_mul_0_0_n75), .B(
        mul_y0y1_gf4_mul_0_0_n74), .Z(mul_y0y1_gf4_mul_0_0_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U26 ( .A(mul_y0y1_gf4_mul_0_0_n73), .B(
        mul_y0y1_gf4_mul_0_0_n72), .ZN(mul_y0y1_FFxDN[2]) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U25 ( .A1(Y1xD[2]), .A2(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_0_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U24 ( .A(mul_y0y1_gf4_mul_0_0_n74), .B(
        mul_y0y1_gf4_mul_0_0_n71), .Z(mul_y0y1_gf4_mul_0_0_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_0_0_U23 ( .A1(mul_y0y1_gf4_mul_0_0_n70), .A2(
        mul_y0y1_gf4_mul_0_0_n69), .ZN(mul_y0y1_gf4_mul_0_0_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U22 ( .A(Y1xD[2]), .B(Y1xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_0_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U21 ( .A(Y0xD[2]), .B(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_0_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U20 ( .A(mul_y0y1_gf4_mul_0_0_n68), .B(
        mul_y0y1_gf4_mul_0_0_n67), .ZN(mul_y0y1_FFxDN[1]) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U19 ( .A1(Y1xD[1]), .A2(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_0_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U18 ( .A(mul_y0y1_gf4_mul_0_0_n75), .B(
        mul_y0y1_gf4_mul_0_0_n66), .Z(mul_y0y1_gf4_mul_0_0_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U17 ( .A(mul_y0y1_gf4_mul_0_0_n65), .B(
        mul_y0y1_gf4_mul_0_0_n64), .ZN(mul_y0y1_gf4_mul_0_0_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U16 ( .A1(mul_y0y1_gf4_mul_0_0_n63), .A2(
        mul_y0y1_gf4_mul_0_0_n62), .ZN(mul_y0y1_gf4_mul_0_0_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U15 ( .A(mul_y0y1_gf4_mul_0_0_n61), .B(
        mul_y0y1_gf4_mul_0_0_n60), .ZN(mul_y0y1_gf4_mul_0_0_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U14 ( .A(mul_y0y1_gf4_mul_0_0_n59), .B(
        mul_y0y1_gf4_mul_0_0_n58), .ZN(mul_y0y1_gf4_mul_0_0_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U13 ( .A(mul_y0y1_gf4_mul_0_0_n57), .B(
        mul_y0y1_gf4_mul_0_0_n56), .ZN(mul_y0y1_FFxDN[0]) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U12 ( .A1(Y1xD[0]), .A2(Y0xD[0]), .ZN(
        mul_y0y1_gf4_mul_0_0_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U11 ( .A(mul_y0y1_gf4_mul_0_0_n66), .B(
        mul_y0y1_gf4_mul_0_0_n71), .Z(mul_y0y1_gf4_mul_0_0_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U10 ( .A(mul_y0y1_gf4_mul_0_0_n55), .B(
        mul_y0y1_gf4_mul_0_0_n65), .ZN(mul_y0y1_gf4_mul_0_0_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_0_0_U9 ( .A1(mul_y0y1_gf4_mul_0_0_n61), .A2(
        mul_y0y1_gf4_mul_0_0_n59), .ZN(mul_y0y1_gf4_mul_0_0_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U8 ( .A(Y1xD[0]), .B(Y1xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_0_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U7 ( .A(Y0xD[0]), .B(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_0_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U6 ( .A1(mul_y0y1_gf4_mul_0_0_n58), .A2(
        mul_y0y1_gf4_mul_0_0_n60), .ZN(mul_y0y1_gf4_mul_0_0_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U5 ( .A(Y0xD[1]), .B(Y0xD[3]), .Z(
        mul_y0y1_gf4_mul_0_0_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U4 ( .A(Y1xD[1]), .B(Y1xD[3]), .Z(
        mul_y0y1_gf4_mul_0_0_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_0_0_U3 ( .A1(mul_y0y1_gf4_mul_0_0_n54), .A2(
        mul_y0y1_gf4_mul_0_0_n53), .ZN(mul_y0y1_gf4_mul_0_0_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U2 ( .A(Y1xD[0]), .B(Y1xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_0_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U1 ( .A(Y0xD[0]), .B(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_0_n54) );
  XNOR2_X1 inverter_gf24_U18 ( .A(inverter_gf24_n3), .B(InverterInxDP[10]), 
        .ZN(inverter_gf24_n10) );
  XNOR2_X1 inverter_gf24_U17 ( .A(inverter_gf24_d_2__0_), .B(InverterInxDP[8]), 
        .ZN(inverter_gf24_n3) );
  XNOR2_X1 inverter_gf24_U16 ( .A(inverter_gf24_n2), .B(InverterInxDP[6]), 
        .ZN(inverter_gf24_n11) );
  XNOR2_X1 inverter_gf24_U15 ( .A(inverter_gf24_d_1__0_), .B(InverterInxDP[4]), 
        .ZN(inverter_gf24_n2) );
  XNOR2_X1 inverter_gf24_U14 ( .A(inverter_gf24_n1), .B(InverterInxDP[2]), 
        .ZN(inverter_gf24_n12) );
  XNOR2_X1 inverter_gf24_U13 ( .A(inverter_gf24_d_0__0_), .B(InverterInxDP[0]), 
        .ZN(inverter_gf24_n1) );
  XOR2_X1 inverter_gf24_U12 ( .A(InverterInxDP[9]), .B(InverterInxDP[11]), .Z(
        inverter_gf24_d_2__0_) );
  XOR2_X1 inverter_gf24_U11 ( .A(InverterInxDP[5]), .B(InverterInxDP[7]), .Z(
        inverter_gf24_d_1__0_) );
  XOR2_X1 inverter_gf24_U10 ( .A(InverterInxDP[1]), .B(InverterInxDP[3]), .Z(
        inverter_gf24_d_0__0_) );
  XNOR2_X1 inverter_gf24_U9 ( .A(inverter_gf24_AmulBxD[4]), .B(
        inverter_gf24_n4), .ZN(inverter_gf24_ExD[5]) );
  XNOR2_X1 inverter_gf24_U8 ( .A(inverter_gf24_AmulBxD[5]), .B(
        inverter_gf24_n5), .ZN(inverter_gf24_ExD[4]) );
  XNOR2_X1 inverter_gf24_U7 ( .A(inverter_gf24_AmulBxD[2]), .B(
        inverter_gf24_n6), .ZN(inverter_gf24_ExD[3]) );
  XNOR2_X1 inverter_gf24_U6 ( .A(inverter_gf24_AmulBxD[3]), .B(
        inverter_gf24_n7), .ZN(inverter_gf24_ExD[2]) );
  XNOR2_X1 inverter_gf24_U5 ( .A(inverter_gf24_AmulBxD[0]), .B(
        inverter_gf24_n8), .ZN(inverter_gf24_ExD[1]) );
  XNOR2_X1 inverter_gf24_U4 ( .A(inverter_gf24_AmulBxD[1]), .B(
        inverter_gf24_n9), .ZN(inverter_gf24_ExD[0]) );
  DFF_X1 inverter_gf24_CxDP_reg_0__0_ ( .D(inverter_gf24_n12), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n8) );
  DFF_X1 inverter_gf24_CxDP_reg_1__0_ ( .D(inverter_gf24_n11), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n6) );
  DFF_X1 inverter_gf24_CxDP_reg_2__0_ ( .D(inverter_gf24_n10), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n4) );
  DFF_X1 inverter_gf24_CxDP_reg_0__1_ ( .D(inverter_gf24_d_0__0_), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n9) );
  DFF_X1 inverter_gf24_CxDP_reg_1__1_ ( .D(inverter_gf24_d_1__0_), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n7) );
  DFF_X1 inverter_gf24_CxDP_reg_2__1_ ( .D(inverter_gf24_d_2__0_), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n5) );
  DFF_X1 inverter_gf24_ExDP_reg_0__0_ ( .D(inverter_gf24_ExD[0]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_0__0_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_0__1_ ( .D(inverter_gf24_ExD[1]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_0__1_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_1__0_ ( .D(inverter_gf24_ExD[2]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_1__0_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_1__1_ ( .D(inverter_gf24_ExD[3]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_1__1_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_2__0_ ( .D(inverter_gf24_ExD[4]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_2__0_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_2__1_ ( .D(inverter_gf24_ExD[5]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_2__1_), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_0__0_ ( .D(InverterInxDP[0]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[0]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_1__0_ ( .D(InverterInxDP[4]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[2]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_2__0_ ( .D(InverterInxDP[8]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[4]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_0__0_ ( .D(InverterInxDP[2]), .CK(ClkxCI), .Q(
        inverter_gf24_AxDP[0]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_1__0_ ( .D(InverterInxDP[6]), .CK(ClkxCI), .Q(
        inverter_gf24_AxDP[2]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_2__0_ ( .D(InverterInxDP[10]), .CK(ClkxCI), 
        .Q(inverter_gf24_AxDP[4]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_0__1_ ( .D(InverterInxDP[3]), .CK(ClkxCI), .Q(
        inverter_gf24_AxDP[1]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_1__1_ ( .D(InverterInxDP[7]), .CK(ClkxCI), .Q(
        inverter_gf24_AxDP[3]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_2__1_ ( .D(InverterInxDP[11]), .CK(ClkxCI), 
        .Q(inverter_gf24_AxDP[5]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_0__1_ ( .D(InverterInxDP[1]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[1]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_1__1_ ( .D(InverterInxDP[5]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[3]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_2__1_ ( .D(InverterInxDP[9]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[5]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_0__0_ ( .D(inverter_gf24_AxDP[0]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[0]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_0__1_ ( .D(inverter_gf24_AxDP[1]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[1]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_1__0_ ( .D(inverter_gf24_AxDP[2]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[2]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_1__1_ ( .D(inverter_gf24_AxDP[3]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[3]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_2__0_ ( .D(inverter_gf24_AxDP[4]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[4]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_2__1_ ( .D(inverter_gf24_AxDP[5]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[5]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_0__0_ ( .D(inverter_gf24_BxDP[0]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[0]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_0__1_ ( .D(inverter_gf24_BxDP[1]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[1]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_1__0_ ( .D(inverter_gf24_BxDP[2]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[2]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_1__1_ ( .D(inverter_gf24_BxDP[3]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[3]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_2__0_ ( .D(inverter_gf24_BxDP[4]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[4]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_2__1_ ( .D(inverter_gf24_BxDP[5]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[5]), .QN() );
  XNOR2_X1 inverter_gf24_a_mul_b_U26 ( .A(inverter_gf24_a_mul_b_n7), .B(
        inverter_gf24_a_mul_b_n6), .ZN(inverter_gf24_AmulBxD[5]) );
  XOR2_X1 inverter_gf24_a_mul_b_U25 ( .A(inverter_gf24_a_mul_b_n9), .B(
        inverter_gf24_a_mul_b_n8), .Z(inverter_gf24_a_mul_b_n6) );
  XNOR2_X1 inverter_gf24_a_mul_b_U24 ( .A(inverter_gf24_a_mul_b_n10), .B(
        inverter_gf24_a_mul_b_n5), .ZN(inverter_gf24_AmulBxD[4]) );
  XOR2_X1 inverter_gf24_a_mul_b_U23 ( .A(inverter_gf24_a_mul_b_n12), .B(
        inverter_gf24_a_mul_b_n11), .Z(inverter_gf24_a_mul_b_n5) );
  XNOR2_X1 inverter_gf24_a_mul_b_U22 ( .A(inverter_gf24_a_mul_b_n13), .B(
        inverter_gf24_a_mul_b_n4), .ZN(inverter_gf24_AmulBxD[3]) );
  XOR2_X1 inverter_gf24_a_mul_b_U21 ( .A(inverter_gf24_a_mul_b_n15), .B(
        inverter_gf24_a_mul_b_n14), .Z(inverter_gf24_a_mul_b_n4) );
  XNOR2_X1 inverter_gf24_a_mul_b_U20 ( .A(inverter_gf24_a_mul_b_n16), .B(
        inverter_gf24_a_mul_b_n3), .ZN(inverter_gf24_AmulBxD[2]) );
  XOR2_X1 inverter_gf24_a_mul_b_U19 ( .A(inverter_gf24_a_mul_b_n18), .B(
        inverter_gf24_a_mul_b_n17), .Z(inverter_gf24_a_mul_b_n3) );
  XNOR2_X1 inverter_gf24_a_mul_b_U18 ( .A(inverter_gf24_a_mul_b_n19), .B(
        inverter_gf24_a_mul_b_n2), .ZN(inverter_gf24_AmulBxD[1]) );
  XOR2_X1 inverter_gf24_a_mul_b_U17 ( .A(inverter_gf24_a_mul_b_n21), .B(
        inverter_gf24_a_mul_b_n20), .Z(inverter_gf24_a_mul_b_n2) );
  XNOR2_X1 inverter_gf24_a_mul_b_U16 ( .A(inverter_gf24_a_mul_b_n22), .B(
        inverter_gf24_a_mul_b_n1), .ZN(inverter_gf24_AmulBxD[0]) );
  XOR2_X1 inverter_gf24_a_mul_b_U15 ( .A(inverter_gf24_a_mul_b_n24), .B(
        inverter_gf24_a_mul_b_n23), .Z(inverter_gf24_a_mul_b_n1) );
  XOR2_X1 inverter_gf24_a_mul_b_U14 ( .A(Zinv1xDI[5]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_7__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[15]) );
  XOR2_X1 inverter_gf24_a_mul_b_U13 ( .A(Zinv1xDI[4]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_7__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[14]) );
  XOR2_X1 inverter_gf24_a_mul_b_U12 ( .A(Zinv1xDI[3]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_6__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[13]) );
  XOR2_X1 inverter_gf24_a_mul_b_U11 ( .A(Zinv1xDI[2]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_6__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[12]) );
  XOR2_X1 inverter_gf24_a_mul_b_U10 ( .A(Zinv1xDI[5]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_5__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[11]) );
  XOR2_X1 inverter_gf24_a_mul_b_U9 ( .A(Zinv1xDI[4]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_5__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[10]) );
  XOR2_X1 inverter_gf24_a_mul_b_U8 ( .A(Zinv1xDI[1]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_3__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[7]) );
  XOR2_X1 inverter_gf24_a_mul_b_U7 ( .A(Zinv1xDI[0]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_3__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[6]) );
  XOR2_X1 inverter_gf24_a_mul_b_U6 ( .A(Zinv1xDI[3]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_2__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[5]) );
  XOR2_X1 inverter_gf24_a_mul_b_U5 ( .A(Zinv1xDI[2]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_2__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[4]) );
  XOR2_X1 inverter_gf24_a_mul_b_U4 ( .A(Zinv1xDI[1]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_1__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[3]) );
  XOR2_X1 inverter_gf24_a_mul_b_U3 ( .A(Zinv1xDI[0]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_1__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[2]) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_1__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[2]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n23) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_1__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[3]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n20) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_2__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[4]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n24) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_2__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[5]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n21) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_3__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[6]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n16) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_3__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[7]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n13) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_5__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[10]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n18) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_5__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[11]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n15) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_6__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[12]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n10) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_6__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[13]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n7) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_7__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[14]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n11) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_7__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[15]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n8) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_0__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[0]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n22) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_0__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[1]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n19) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_4__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[8]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n17) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_4__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[9]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n14) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_8__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[16]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n12) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_8__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[17]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n9) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[17]) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U6 ( .A1(InverterInxDP[11]), .A2(
        InverterInxDP[9]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[16]) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U3 ( .A(InverterInxDP[11]), .B(
        InverterInxDP[10]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U2 ( .A(InverterInxDP[9]), .B(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U1 ( .A1(InverterInxDP[10]), .A2(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_7__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U6 ( .A1(InverterInxDP[11]), .A2(
        InverterInxDP[5]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_7__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U3 ( .A(InverterInxDP[11]), .B(
        InverterInxDP[10]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U2 ( .A(InverterInxDP[5]), .B(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U1 ( .A1(InverterInxDP[10]), .A2(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_6__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U6 ( .A1(InverterInxDP[11]), .A2(
        InverterInxDP[1]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_6__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U3 ( .A(InverterInxDP[11]), .B(
        InverterInxDP[10]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U2 ( .A(InverterInxDP[1]), .B(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U1 ( .A1(InverterInxDP[10]), .A2(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_5__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U6 ( .A1(InverterInxDP[7]), .A2(
        InverterInxDP[9]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_5__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U3 ( .A(InverterInxDP[7]), .B(
        InverterInxDP[6]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U2 ( .A(InverterInxDP[9]), .B(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U1 ( .A1(InverterInxDP[6]), .A2(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[9]) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U6 ( .A1(InverterInxDP[7]), .A2(
        InverterInxDP[5]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[8]) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U3 ( .A(InverterInxDP[7]), .B(
        InverterInxDP[6]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U2 ( .A(InverterInxDP[5]), .B(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U1 ( .A1(InverterInxDP[6]), .A2(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_3__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U6 ( .A1(InverterInxDP[7]), .A2(
        InverterInxDP[1]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_3__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U3 ( .A(InverterInxDP[7]), .B(
        InverterInxDP[6]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U2 ( .A(InverterInxDP[1]), .B(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U1 ( .A1(InverterInxDP[6]), .A2(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_2__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U6 ( .A1(InverterInxDP[3]), .A2(
        InverterInxDP[9]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_2__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U3 ( .A(InverterInxDP[3]), .B(
        InverterInxDP[2]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U2 ( .A(InverterInxDP[9]), .B(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U1 ( .A1(InverterInxDP[2]), .A2(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_1__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U6 ( .A1(InverterInxDP[3]), .A2(
        InverterInxDP[5]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_1__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U3 ( .A(InverterInxDP[3]), .B(
        InverterInxDP[2]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U2 ( .A(InverterInxDP[5]), .B(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U1 ( .A1(InverterInxDP[2]), .A2(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[1]) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U6 ( .A1(InverterInxDP[3]), .A2(
        InverterInxDP[1]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[0]) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U3 ( .A(InverterInxDP[3]), .B(
        InverterInxDP[2]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U2 ( .A(InverterInxDP[1]), .B(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U1 ( .A1(InverterInxDP[2]), .A2(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_0_n13) );
  XOR2_X1 inverter_gf24_a_mul_e_U32 ( .A(inverter_gf24_a_mul_e_n22), .B(
        inverter_gf24_a_mul_e_n8), .Z(inverter_gf24_a_mul_e_n39) );
  XOR2_X1 inverter_gf24_a_mul_e_U31 ( .A(inverter_gf24_a_mul_e_n19), .B(
        inverter_gf24_a_mul_e_n10), .Z(inverter_gf24_a_mul_e_n38) );
  XOR2_X1 inverter_gf24_a_mul_e_U30 ( .A(inverter_gf24_a_mul_e_n23), .B(
        inverter_gf24_a_mul_e_n12), .Z(inverter_gf24_a_mul_e_n37) );
  XOR2_X1 inverter_gf24_a_mul_e_U29 ( .A(inverter_gf24_a_mul_e_n20), .B(
        inverter_gf24_a_mul_e_n14), .Z(inverter_gf24_a_mul_e_n36) );
  XOR2_X1 inverter_gf24_a_mul_e_U28 ( .A(inverter_gf24_a_mul_e_n24), .B(
        inverter_gf24_a_mul_e_n16), .Z(inverter_gf24_a_mul_e_n35) );
  XOR2_X1 inverter_gf24_a_mul_e_U27 ( .A(inverter_gf24_a_mul_e_n21), .B(
        inverter_gf24_a_mul_e_n18), .Z(inverter_gf24_a_mul_e_n34) );
  XOR2_X1 inverter_gf24_a_mul_e_U26 ( .A(Zinv2xDI[5]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_7__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[15]) );
  XOR2_X1 inverter_gf24_a_mul_e_U25 ( .A(Zinv2xDI[4]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_7__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[14]) );
  XOR2_X1 inverter_gf24_a_mul_e_U24 ( .A(Zinv2xDI[3]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_6__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[13]) );
  XOR2_X1 inverter_gf24_a_mul_e_U23 ( .A(Zinv2xDI[2]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_6__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[12]) );
  XOR2_X1 inverter_gf24_a_mul_e_U22 ( .A(Zinv2xDI[5]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_5__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[11]) );
  XOR2_X1 inverter_gf24_a_mul_e_U21 ( .A(Zinv2xDI[4]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_5__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[10]) );
  XOR2_X1 inverter_gf24_a_mul_e_U20 ( .A(Zinv2xDI[1]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_3__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[7]) );
  XOR2_X1 inverter_gf24_a_mul_e_U19 ( .A(Zinv2xDI[0]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_3__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[6]) );
  XOR2_X1 inverter_gf24_a_mul_e_U18 ( .A(Zinv2xDI[3]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_2__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[5]) );
  XOR2_X1 inverter_gf24_a_mul_e_U17 ( .A(Zinv2xDI[2]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_2__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[4]) );
  XOR2_X1 inverter_gf24_a_mul_e_U16 ( .A(Zinv2xDI[1]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_1__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[3]) );
  XOR2_X1 inverter_gf24_a_mul_e_U15 ( .A(Zinv2xDI[0]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_1__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[2]) );
  INV_X1 inverter_gf24_a_mul_e_U14 ( .A(inverter_gf24_a_mul_e_n42), .ZN(
        InverterOutxD[0]) );
  XOR2_X1 inverter_gf24_a_mul_e_U13 ( .A(inverter_gf24_a_mul_e_n17), .B(
        inverter_gf24_a_mul_e_n34), .Z(inverter_gf24_a_mul_e_n42) );
  INV_X1 inverter_gf24_a_mul_e_U12 ( .A(inverter_gf24_a_mul_e_n41), .ZN(
        InverterOutxD[4]) );
  XOR2_X1 inverter_gf24_a_mul_e_U11 ( .A(inverter_gf24_a_mul_e_n13), .B(
        inverter_gf24_a_mul_e_n36), .Z(inverter_gf24_a_mul_e_n41) );
  INV_X1 inverter_gf24_a_mul_e_U10 ( .A(inverter_gf24_a_mul_e_n40), .ZN(
        InverterOutxD[8]) );
  XOR2_X1 inverter_gf24_a_mul_e_U9 ( .A(inverter_gf24_a_mul_e_n9), .B(
        inverter_gf24_a_mul_e_n38), .Z(inverter_gf24_a_mul_e_n40) );
  INV_X1 inverter_gf24_a_mul_e_U8 ( .A(inverter_gf24_a_mul_e_n27), .ZN(
        InverterOutxD[9]) );
  INV_X1 inverter_gf24_a_mul_e_U7 ( .A(inverter_gf24_a_mul_e_n26), .ZN(
        InverterOutxD[1]) );
  INV_X1 inverter_gf24_a_mul_e_U6 ( .A(inverter_gf24_a_mul_e_n25), .ZN(
        InverterOutxD[5]) );
  XOR2_X1 inverter_gf24_a_mul_e_U5 ( .A(inverter_gf24_a_mul_e_n7), .B(
        inverter_gf24_a_mul_e_n39), .Z(inverter_gf24_a_mul_e_n27) );
  XOR2_X1 inverter_gf24_a_mul_e_U4 ( .A(inverter_gf24_a_mul_e_n15), .B(
        inverter_gf24_a_mul_e_n35), .Z(inverter_gf24_a_mul_e_n26) );
  XOR2_X1 inverter_gf24_a_mul_e_U3 ( .A(inverter_gf24_a_mul_e_n11), .B(
        inverter_gf24_a_mul_e_n37), .Z(inverter_gf24_a_mul_e_n25) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_1__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[2]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n17) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_1__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[3]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n15) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_2__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[4]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n18) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_2__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[5]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n16) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_3__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[6]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n20) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_3__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[7]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n23) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_5__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[10]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n14) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_5__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[11]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n12) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_6__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[12]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n19) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_6__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[13]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n22) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_7__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[14]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n9) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_7__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[15]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n7) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_0__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[0]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n21) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_4__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[8]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n13) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_8__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[16]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n10) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_0__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[1]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n24) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_4__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[9]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n11) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_8__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[17]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n8) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[17]) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[5]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[16]) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U3 ( .A(
        inverter_gf24_pipelinedAxDP[5]), .B(inverter_gf24_pipelinedAxDP[4]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_2_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[4]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_7__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[5]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_7__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U3 ( .A(
        inverter_gf24_pipelinedAxDP[5]), .B(inverter_gf24_pipelinedAxDP[4]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_2_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[4]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_6__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[5]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_6__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U3 ( .A(
        inverter_gf24_pipelinedAxDP[5]), .B(inverter_gf24_pipelinedAxDP[4]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_2_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[4]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_5__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[3]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_5__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U3 ( .A(
        inverter_gf24_pipelinedAxDP[3]), .B(inverter_gf24_pipelinedAxDP[2]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_1_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[2]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[9]) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[3]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[8]) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U3 ( .A(
        inverter_gf24_pipelinedAxDP[3]), .B(inverter_gf24_pipelinedAxDP[2]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_1_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[2]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_3__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[3]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_3__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U3 ( .A(
        inverter_gf24_pipelinedAxDP[3]), .B(inverter_gf24_pipelinedAxDP[2]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_1_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[2]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_2__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[1]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_2__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U3 ( .A(
        inverter_gf24_pipelinedAxDP[1]), .B(inverter_gf24_pipelinedAxDP[0]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_0_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[0]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_1__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[1]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_1__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U3 ( .A(
        inverter_gf24_pipelinedAxDP[1]), .B(inverter_gf24_pipelinedAxDP[0]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_0_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[0]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[1]) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[1]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[0]) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U3 ( .A(
        inverter_gf24_pipelinedAxDP[1]), .B(inverter_gf24_pipelinedAxDP[0]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_0_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[0]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n13) );
  XOR2_X1 inverter_gf24_b_mul_e_U32 ( .A(inverter_gf24_b_mul_e_n19), .B(
        inverter_gf24_b_mul_e_n8), .Z(inverter_gf24_b_mul_e_n39) );
  XOR2_X1 inverter_gf24_b_mul_e_U31 ( .A(inverter_gf24_b_mul_e_n22), .B(
        inverter_gf24_b_mul_e_n10), .Z(inverter_gf24_b_mul_e_n38) );
  XOR2_X1 inverter_gf24_b_mul_e_U30 ( .A(inverter_gf24_b_mul_e_n20), .B(
        inverter_gf24_b_mul_e_n12), .Z(inverter_gf24_b_mul_e_n37) );
  XOR2_X1 inverter_gf24_b_mul_e_U29 ( .A(inverter_gf24_b_mul_e_n23), .B(
        inverter_gf24_b_mul_e_n14), .Z(inverter_gf24_b_mul_e_n36) );
  XOR2_X1 inverter_gf24_b_mul_e_U28 ( .A(inverter_gf24_b_mul_e_n21), .B(
        inverter_gf24_b_mul_e_n16), .Z(inverter_gf24_b_mul_e_n35) );
  XOR2_X1 inverter_gf24_b_mul_e_U27 ( .A(inverter_gf24_b_mul_e_n24), .B(
        inverter_gf24_b_mul_e_n18), .Z(inverter_gf24_b_mul_e_n34) );
  XOR2_X1 inverter_gf24_b_mul_e_U26 ( .A(Zinv3xDI[5]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_7__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[15]) );
  XOR2_X1 inverter_gf24_b_mul_e_U25 ( .A(Zinv3xDI[4]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_7__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[14]) );
  XOR2_X1 inverter_gf24_b_mul_e_U24 ( .A(Zinv3xDI[3]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_6__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[13]) );
  XOR2_X1 inverter_gf24_b_mul_e_U23 ( .A(Zinv3xDI[2]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_6__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[12]) );
  XOR2_X1 inverter_gf24_b_mul_e_U22 ( .A(Zinv3xDI[5]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_5__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[11]) );
  XOR2_X1 inverter_gf24_b_mul_e_U21 ( .A(Zinv3xDI[4]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_5__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[10]) );
  XOR2_X1 inverter_gf24_b_mul_e_U20 ( .A(Zinv3xDI[1]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_3__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[7]) );
  XOR2_X1 inverter_gf24_b_mul_e_U19 ( .A(Zinv3xDI[0]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_3__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[6]) );
  XOR2_X1 inverter_gf24_b_mul_e_U18 ( .A(Zinv3xDI[3]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_2__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[5]) );
  XOR2_X1 inverter_gf24_b_mul_e_U17 ( .A(Zinv3xDI[2]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_2__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[4]) );
  XOR2_X1 inverter_gf24_b_mul_e_U16 ( .A(Zinv3xDI[1]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_1__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[3]) );
  XOR2_X1 inverter_gf24_b_mul_e_U15 ( .A(Zinv3xDI[0]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_1__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[2]) );
  INV_X1 inverter_gf24_b_mul_e_U14 ( .A(inverter_gf24_b_mul_e_n42), .ZN(
        InverterOutxD[3]) );
  XOR2_X1 inverter_gf24_b_mul_e_U13 ( .A(inverter_gf24_b_mul_e_n15), .B(
        inverter_gf24_b_mul_e_n35), .Z(inverter_gf24_b_mul_e_n42) );
  INV_X1 inverter_gf24_b_mul_e_U12 ( .A(inverter_gf24_b_mul_e_n41), .ZN(
        InverterOutxD[7]) );
  XOR2_X1 inverter_gf24_b_mul_e_U11 ( .A(inverter_gf24_b_mul_e_n11), .B(
        inverter_gf24_b_mul_e_n37), .Z(inverter_gf24_b_mul_e_n41) );
  INV_X1 inverter_gf24_b_mul_e_U10 ( .A(inverter_gf24_b_mul_e_n40), .ZN(
        InverterOutxD[11]) );
  XOR2_X1 inverter_gf24_b_mul_e_U9 ( .A(inverter_gf24_b_mul_e_n7), .B(
        inverter_gf24_b_mul_e_n39), .Z(inverter_gf24_b_mul_e_n40) );
  INV_X1 inverter_gf24_b_mul_e_U8 ( .A(inverter_gf24_b_mul_e_n27), .ZN(
        InverterOutxD[10]) );
  INV_X1 inverter_gf24_b_mul_e_U7 ( .A(inverter_gf24_b_mul_e_n26), .ZN(
        InverterOutxD[2]) );
  INV_X1 inverter_gf24_b_mul_e_U6 ( .A(inverter_gf24_b_mul_e_n25), .ZN(
        InverterOutxD[6]) );
  XOR2_X1 inverter_gf24_b_mul_e_U5 ( .A(inverter_gf24_b_mul_e_n9), .B(
        inverter_gf24_b_mul_e_n38), .Z(inverter_gf24_b_mul_e_n27) );
  XOR2_X1 inverter_gf24_b_mul_e_U4 ( .A(inverter_gf24_b_mul_e_n17), .B(
        inverter_gf24_b_mul_e_n34), .Z(inverter_gf24_b_mul_e_n26) );
  XOR2_X1 inverter_gf24_b_mul_e_U3 ( .A(inverter_gf24_b_mul_e_n13), .B(
        inverter_gf24_b_mul_e_n36), .Z(inverter_gf24_b_mul_e_n25) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_1__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[2]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n17) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_1__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[3]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n15) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_2__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[4]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n18) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_2__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[5]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n16) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_3__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[6]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n23) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_3__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[7]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n20) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_5__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[10]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n14) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_5__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[11]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n12) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_6__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[12]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n22) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_6__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[13]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n19) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_7__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[14]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n9) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_7__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[15]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n7) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_0__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[0]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n24) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_4__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[8]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n13) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_8__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[16]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n10) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_0__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[1]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n21) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_4__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[9]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n11) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_8__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[17]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n8) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[17]) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[5]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[16]) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U3 ( .A(
        inverter_gf24_pipelinedBxDP[5]), .B(inverter_gf24_pipelinedBxDP[4]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_2_2_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[4]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_7__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[5]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_7__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U3 ( .A(
        inverter_gf24_pipelinedBxDP[5]), .B(inverter_gf24_pipelinedBxDP[4]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_2_1_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[4]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_6__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[5]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_6__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U3 ( .A(
        inverter_gf24_pipelinedBxDP[5]), .B(inverter_gf24_pipelinedBxDP[4]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_2_0_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[4]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_5__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[3]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_5__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U3 ( .A(
        inverter_gf24_pipelinedBxDP[3]), .B(inverter_gf24_pipelinedBxDP[2]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_1_2_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[2]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[9]) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[3]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[8]) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U3 ( .A(
        inverter_gf24_pipelinedBxDP[3]), .B(inverter_gf24_pipelinedBxDP[2]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_1_1_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[2]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_3__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[3]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_3__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U3 ( .A(
        inverter_gf24_pipelinedBxDP[3]), .B(inverter_gf24_pipelinedBxDP[2]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_1_0_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[2]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_2__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[1]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_2__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U3 ( .A(
        inverter_gf24_pipelinedBxDP[1]), .B(inverter_gf24_pipelinedBxDP[0]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_0_2_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[0]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_1__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[1]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_1__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U3 ( .A(
        inverter_gf24_pipelinedBxDP[1]), .B(inverter_gf24_pipelinedBxDP[0]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_0_1_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[0]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[1]) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[1]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[0]) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U3 ( .A(
        inverter_gf24_pipelinedBxDP[1]), .B(inverter_gf24_pipelinedBxDP[0]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_0_0_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[0]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n13) );
  XNOR2_X1 mult_msb_U50 ( .A(mult_msb_n13), .B(mult_msb_n60), .ZN(
        InvUnmappedxD[23]) );
  XOR2_X1 mult_msb_U49 ( .A(mult_msb_n15), .B(mult_msb_n14), .Z(mult_msb_n60)
         );
  XNOR2_X1 mult_msb_U48 ( .A(mult_msb_n16), .B(mult_msb_n59), .ZN(
        InvUnmappedxD[22]) );
  XOR2_X1 mult_msb_U47 ( .A(mult_msb_n18), .B(mult_msb_n17), .Z(mult_msb_n59)
         );
  XNOR2_X1 mult_msb_U46 ( .A(mult_msb_n19), .B(mult_msb_n58), .ZN(
        InvUnmappedxD[21]) );
  XOR2_X1 mult_msb_U45 ( .A(mult_msb_n21), .B(mult_msb_n20), .Z(mult_msb_n58)
         );
  XNOR2_X1 mult_msb_U44 ( .A(mult_msb_n22), .B(mult_msb_n57), .ZN(
        InvUnmappedxD[20]) );
  XOR2_X1 mult_msb_U43 ( .A(mult_msb_n24), .B(mult_msb_n23), .Z(mult_msb_n57)
         );
  XNOR2_X1 mult_msb_U42 ( .A(mult_msb_n25), .B(mult_msb_n56), .ZN(
        InvUnmappedxD[15]) );
  XOR2_X1 mult_msb_U41 ( .A(mult_msb_n27), .B(mult_msb_n26), .Z(mult_msb_n56)
         );
  XNOR2_X1 mult_msb_U40 ( .A(mult_msb_n28), .B(mult_msb_n55), .ZN(
        InvUnmappedxD[14]) );
  XOR2_X1 mult_msb_U39 ( .A(mult_msb_n30), .B(mult_msb_n29), .Z(mult_msb_n55)
         );
  XNOR2_X1 mult_msb_U38 ( .A(mult_msb_n31), .B(mult_msb_n54), .ZN(
        InvUnmappedxD[13]) );
  XOR2_X1 mult_msb_U37 ( .A(mult_msb_n33), .B(mult_msb_n32), .Z(mult_msb_n54)
         );
  XNOR2_X1 mult_msb_U36 ( .A(mult_msb_n34), .B(mult_msb_n53), .ZN(
        InvUnmappedxD[12]) );
  XOR2_X1 mult_msb_U35 ( .A(mult_msb_n36), .B(mult_msb_n35), .Z(mult_msb_n53)
         );
  XNOR2_X1 mult_msb_U34 ( .A(mult_msb_n37), .B(mult_msb_n52), .ZN(
        InvUnmappedxD[7]) );
  XOR2_X1 mult_msb_U33 ( .A(mult_msb_n39), .B(mult_msb_n38), .Z(mult_msb_n52)
         );
  XNOR2_X1 mult_msb_U32 ( .A(mult_msb_n40), .B(mult_msb_n51), .ZN(
        InvUnmappedxD[6]) );
  XOR2_X1 mult_msb_U31 ( .A(mult_msb_n42), .B(mult_msb_n41), .Z(mult_msb_n51)
         );
  XNOR2_X1 mult_msb_U30 ( .A(mult_msb_n43), .B(mult_msb_n50), .ZN(
        InvUnmappedxD[5]) );
  XOR2_X1 mult_msb_U29 ( .A(mult_msb_n45), .B(mult_msb_n44), .Z(mult_msb_n50)
         );
  XNOR2_X1 mult_msb_U28 ( .A(mult_msb_n46), .B(mult_msb_n49), .ZN(
        InvUnmappedxD[4]) );
  XOR2_X1 mult_msb_U27 ( .A(mult_msb_n48), .B(mult_msb_n47), .Z(mult_msb_n49)
         );
  XOR2_X1 mult_msb_U26 ( .A(Zmul2xDI[11]), .B(mult_msb_Xi_mul_Yj_7__3_), .Z(
        mult_msb_FFxDN[31]) );
  XOR2_X1 mult_msb_U25 ( .A(Zmul2xDI[10]), .B(mult_msb_Xi_mul_Yj_7__2_), .Z(
        mult_msb_FFxDN[30]) );
  XOR2_X1 mult_msb_U24 ( .A(Zmul2xDI[9]), .B(mult_msb_Xi_mul_Yj_7__1_), .Z(
        mult_msb_FFxDN[29]) );
  XOR2_X1 mult_msb_U23 ( .A(Zmul2xDI[8]), .B(mult_msb_Xi_mul_Yj_7__0_), .Z(
        mult_msb_FFxDN[28]) );
  XOR2_X1 mult_msb_U22 ( .A(Zmul2xDI[7]), .B(mult_msb_Xi_mul_Yj_6__3_), .Z(
        mult_msb_FFxDN[27]) );
  XOR2_X1 mult_msb_U21 ( .A(Zmul2xDI[6]), .B(mult_msb_Xi_mul_Yj_6__2_), .Z(
        mult_msb_FFxDN[26]) );
  XOR2_X1 mult_msb_U20 ( .A(Zmul2xDI[5]), .B(mult_msb_Xi_mul_Yj_6__1_), .Z(
        mult_msb_FFxDN[25]) );
  XOR2_X1 mult_msb_U19 ( .A(Zmul2xDI[4]), .B(mult_msb_Xi_mul_Yj_6__0_), .Z(
        mult_msb_FFxDN[24]) );
  XOR2_X1 mult_msb_U18 ( .A(Zmul2xDI[11]), .B(mult_msb_Xi_mul_Yj_5__3_), .Z(
        mult_msb_FFxDN[23]) );
  XOR2_X1 mult_msb_U17 ( .A(Zmul2xDI[10]), .B(mult_msb_Xi_mul_Yj_5__2_), .Z(
        mult_msb_FFxDN[22]) );
  XOR2_X1 mult_msb_U16 ( .A(Zmul2xDI[9]), .B(mult_msb_Xi_mul_Yj_5__1_), .Z(
        mult_msb_FFxDN[21]) );
  XOR2_X1 mult_msb_U15 ( .A(Zmul2xDI[8]), .B(mult_msb_Xi_mul_Yj_5__0_), .Z(
        mult_msb_FFxDN[20]) );
  XOR2_X1 mult_msb_U14 ( .A(Zmul2xDI[3]), .B(mult_msb_Xi_mul_Yj_3__3_), .Z(
        mult_msb_FFxDN[15]) );
  XOR2_X1 mult_msb_U13 ( .A(Zmul2xDI[2]), .B(mult_msb_Xi_mul_Yj_3__2_), .Z(
        mult_msb_FFxDN[14]) );
  XOR2_X1 mult_msb_U12 ( .A(Zmul2xDI[1]), .B(mult_msb_Xi_mul_Yj_3__1_), .Z(
        mult_msb_FFxDN[13]) );
  XOR2_X1 mult_msb_U11 ( .A(Zmul2xDI[0]), .B(mult_msb_Xi_mul_Yj_3__0_), .Z(
        mult_msb_FFxDN[12]) );
  XOR2_X1 mult_msb_U10 ( .A(Zmul2xDI[7]), .B(mult_msb_Xi_mul_Yj_2__3_), .Z(
        mult_msb_FFxDN[11]) );
  XOR2_X1 mult_msb_U9 ( .A(Zmul2xDI[6]), .B(mult_msb_Xi_mul_Yj_2__2_), .Z(
        mult_msb_FFxDN[10]) );
  XOR2_X1 mult_msb_U8 ( .A(Zmul2xDI[5]), .B(mult_msb_Xi_mul_Yj_2__1_), .Z(
        mult_msb_FFxDN[9]) );
  XOR2_X1 mult_msb_U7 ( .A(Zmul2xDI[4]), .B(mult_msb_Xi_mul_Yj_2__0_), .Z(
        mult_msb_FFxDN[8]) );
  XOR2_X1 mult_msb_U6 ( .A(Zmul2xDI[3]), .B(mult_msb_Xi_mul_Yj_1__3_), .Z(
        mult_msb_FFxDN[7]) );
  XOR2_X1 mult_msb_U5 ( .A(Zmul2xDI[2]), .B(mult_msb_Xi_mul_Yj_1__2_), .Z(
        mult_msb_FFxDN[6]) );
  XOR2_X1 mult_msb_U4 ( .A(Zmul2xDI[1]), .B(mult_msb_Xi_mul_Yj_1__1_), .Z(
        mult_msb_FFxDN[5]) );
  XOR2_X1 mult_msb_U3 ( .A(Zmul2xDI[0]), .B(mult_msb_Xi_mul_Yj_1__0_), .Z(
        mult_msb_FFxDN[4]) );
  DFF_X1 mult_msb_FFxDP_reg_1__3_ ( .D(mult_msb_FFxDN[7]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n38) );
  DFF_X1 mult_msb_FFxDP_reg_2__3_ ( .D(mult_msb_FFxDN[11]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n39) );
  DFF_X1 mult_msb_FFxDP_reg_3__3_ ( .D(mult_msb_FFxDN[15]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n25) );
  DFF_X1 mult_msb_FFxDP_reg_5__3_ ( .D(mult_msb_FFxDN[23]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n27) );
  DFF_X1 mult_msb_FFxDP_reg_6__3_ ( .D(mult_msb_FFxDN[27]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n13) );
  DFF_X1 mult_msb_FFxDP_reg_7__3_ ( .D(mult_msb_FFxDN[31]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n14) );
  DFF_X1 mult_msb_FFxDP_reg_1__1_ ( .D(mult_msb_FFxDN[5]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n44) );
  DFF_X1 mult_msb_FFxDP_reg_2__1_ ( .D(mult_msb_FFxDN[9]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n45) );
  DFF_X1 mult_msb_FFxDP_reg_3__1_ ( .D(mult_msb_FFxDN[13]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n31) );
  DFF_X1 mult_msb_FFxDP_reg_5__1_ ( .D(mult_msb_FFxDN[21]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n33) );
  DFF_X1 mult_msb_FFxDP_reg_6__1_ ( .D(mult_msb_FFxDN[25]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n19) );
  DFF_X1 mult_msb_FFxDP_reg_7__1_ ( .D(mult_msb_FFxDN[29]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n20) );
  DFF_X1 mult_msb_FFxDP_reg_1__2_ ( .D(mult_msb_FFxDN[6]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n41) );
  DFF_X1 mult_msb_FFxDP_reg_2__2_ ( .D(mult_msb_FFxDN[10]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n42) );
  DFF_X1 mult_msb_FFxDP_reg_3__2_ ( .D(mult_msb_FFxDN[14]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n28) );
  DFF_X1 mult_msb_FFxDP_reg_5__2_ ( .D(mult_msb_FFxDN[22]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n30) );
  DFF_X1 mult_msb_FFxDP_reg_6__2_ ( .D(mult_msb_FFxDN[26]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n16) );
  DFF_X1 mult_msb_FFxDP_reg_7__2_ ( .D(mult_msb_FFxDN[30]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n17) );
  DFF_X1 mult_msb_FFxDP_reg_1__0_ ( .D(mult_msb_FFxDN[4]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n47) );
  DFF_X1 mult_msb_FFxDP_reg_2__0_ ( .D(mult_msb_FFxDN[8]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n48) );
  DFF_X1 mult_msb_FFxDP_reg_3__0_ ( .D(mult_msb_FFxDN[12]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n34) );
  DFF_X1 mult_msb_FFxDP_reg_5__0_ ( .D(mult_msb_FFxDN[20]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n36) );
  DFF_X1 mult_msb_FFxDP_reg_6__0_ ( .D(mult_msb_FFxDN[24]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n22) );
  DFF_X1 mult_msb_FFxDP_reg_7__0_ ( .D(mult_msb_FFxDN[28]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n23) );
  DFF_X1 mult_msb_FFxDP_reg_0__3_ ( .D(mult_msb_FFxDN[3]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n37) );
  DFF_X1 mult_msb_FFxDP_reg_4__3_ ( .D(mult_msb_FFxDN[19]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n26) );
  DFF_X1 mult_msb_FFxDP_reg_8__3_ ( .D(mult_msb_FFxDN[35]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n15) );
  DFF_X1 mult_msb_FFxDP_reg_0__1_ ( .D(mult_msb_FFxDN[1]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n43) );
  DFF_X1 mult_msb_FFxDP_reg_4__1_ ( .D(mult_msb_FFxDN[17]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n32) );
  DFF_X1 mult_msb_FFxDP_reg_8__1_ ( .D(mult_msb_FFxDN[33]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n21) );
  DFF_X1 mult_msb_FFxDP_reg_0__2_ ( .D(mult_msb_FFxDN[2]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n40) );
  DFF_X1 mult_msb_FFxDP_reg_4__2_ ( .D(mult_msb_FFxDN[18]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n29) );
  DFF_X1 mult_msb_FFxDP_reg_8__2_ ( .D(mult_msb_FFxDN[34]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n18) );
  DFF_X1 mult_msb_FFxDP_reg_0__0_ ( .D(mult_msb_FFxDN[0]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n46) );
  DFF_X1 mult_msb_FFxDP_reg_4__0_ ( .D(mult_msb_FFxDN[16]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n35) );
  DFF_X1 mult_msb_FFxDP_reg_8__0_ ( .D(mult_msb_FFxDN[32]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n24) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U29 ( .A(mult_msb_gf4_mul_2_2_n77), .B(
        mult_msb_gf4_mul_2_2_n76), .ZN(mult_msb_FFxDN[35]) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U28 ( .A1(InverterOutxD[11]), .A2(Y0_4xDP[11]), 
        .ZN(mult_msb_gf4_mul_2_2_n76) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U27 ( .A(mult_msb_gf4_mul_2_2_n75), .B(
        mult_msb_gf4_mul_2_2_n74), .Z(mult_msb_gf4_mul_2_2_n77) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U26 ( .A(mult_msb_gf4_mul_2_2_n73), .B(
        mult_msb_gf4_mul_2_2_n72), .ZN(mult_msb_FFxDN[34]) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U25 ( .A1(InverterOutxD[10]), .A2(Y0_4xDP[10]), 
        .ZN(mult_msb_gf4_mul_2_2_n72) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U24 ( .A(mult_msb_gf4_mul_2_2_n74), .B(
        mult_msb_gf4_mul_2_2_n71), .Z(mult_msb_gf4_mul_2_2_n73) );
  NOR2_X1 mult_msb_gf4_mul_2_2_U23 ( .A1(mult_msb_gf4_mul_2_2_n70), .A2(
        mult_msb_gf4_mul_2_2_n69), .ZN(mult_msb_gf4_mul_2_2_n74) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U22 ( .A(InverterOutxD[10]), .B(
        InverterOutxD[11]), .ZN(mult_msb_gf4_mul_2_2_n69) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U21 ( .A(Y0_4xDP[10]), .B(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_2_2_n70) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U20 ( .A(mult_msb_gf4_mul_2_2_n68), .B(
        mult_msb_gf4_mul_2_2_n67), .ZN(mult_msb_FFxDN[33]) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U19 ( .A1(InverterOutxD[9]), .A2(Y0_4xDP[9]), 
        .ZN(mult_msb_gf4_mul_2_2_n67) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U18 ( .A(mult_msb_gf4_mul_2_2_n75), .B(
        mult_msb_gf4_mul_2_2_n66), .Z(mult_msb_gf4_mul_2_2_n68) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U17 ( .A(mult_msb_gf4_mul_2_2_n65), .B(
        mult_msb_gf4_mul_2_2_n64), .ZN(mult_msb_gf4_mul_2_2_n75) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U16 ( .A1(mult_msb_gf4_mul_2_2_n63), .A2(
        mult_msb_gf4_mul_2_2_n62), .ZN(mult_msb_gf4_mul_2_2_n64) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U15 ( .A(mult_msb_gf4_mul_2_2_n61), .B(
        mult_msb_gf4_mul_2_2_n60), .ZN(mult_msb_gf4_mul_2_2_n62) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U14 ( .A(mult_msb_gf4_mul_2_2_n59), .B(
        mult_msb_gf4_mul_2_2_n58), .ZN(mult_msb_gf4_mul_2_2_n63) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U13 ( .A(mult_msb_gf4_mul_2_2_n57), .B(
        mult_msb_gf4_mul_2_2_n56), .ZN(mult_msb_FFxDN[32]) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U12 ( .A1(InverterOutxD[8]), .A2(Y0_4xDP[8]), 
        .ZN(mult_msb_gf4_mul_2_2_n56) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U11 ( .A(mult_msb_gf4_mul_2_2_n66), .B(
        mult_msb_gf4_mul_2_2_n71), .Z(mult_msb_gf4_mul_2_2_n57) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U10 ( .A(mult_msb_gf4_mul_2_2_n55), .B(
        mult_msb_gf4_mul_2_2_n65), .ZN(mult_msb_gf4_mul_2_2_n71) );
  NOR2_X1 mult_msb_gf4_mul_2_2_U9 ( .A1(mult_msb_gf4_mul_2_2_n61), .A2(
        mult_msb_gf4_mul_2_2_n59), .ZN(mult_msb_gf4_mul_2_2_n65) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U8 ( .A(InverterOutxD[8]), .B(
        InverterOutxD[10]), .ZN(mult_msb_gf4_mul_2_2_n59) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U7 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_2_2_n61) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U6 ( .A1(mult_msb_gf4_mul_2_2_n58), .A2(
        mult_msb_gf4_mul_2_2_n60), .ZN(mult_msb_gf4_mul_2_2_n55) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U5 ( .A(Y0_4xDP[9]), .B(Y0_4xDP[11]), .Z(
        mult_msb_gf4_mul_2_2_n60) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U4 ( .A(InverterOutxD[9]), .B(InverterOutxD[11]), .Z(mult_msb_gf4_mul_2_2_n58) );
  NOR2_X1 mult_msb_gf4_mul_2_2_U3 ( .A1(mult_msb_gf4_mul_2_2_n54), .A2(
        mult_msb_gf4_mul_2_2_n53), .ZN(mult_msb_gf4_mul_2_2_n66) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U2 ( .A(InverterOutxD[8]), .B(InverterOutxD[9]), .ZN(mult_msb_gf4_mul_2_2_n53) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U1 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_2_2_n54) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U29 ( .A(mult_msb_gf4_mul_2_1_n77), .B(
        mult_msb_gf4_mul_2_1_n76), .ZN(mult_msb_Xi_mul_Yj_7__3_) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U28 ( .A1(InverterOutxD[11]), .A2(Y0_4xDP[7]), 
        .ZN(mult_msb_gf4_mul_2_1_n76) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U27 ( .A(mult_msb_gf4_mul_2_1_n75), .B(
        mult_msb_gf4_mul_2_1_n74), .Z(mult_msb_gf4_mul_2_1_n77) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U26 ( .A(mult_msb_gf4_mul_2_1_n73), .B(
        mult_msb_gf4_mul_2_1_n72), .ZN(mult_msb_Xi_mul_Yj_7__2_) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U25 ( .A1(InverterOutxD[10]), .A2(Y0_4xDP[6]), 
        .ZN(mult_msb_gf4_mul_2_1_n72) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U24 ( .A(mult_msb_gf4_mul_2_1_n74), .B(
        mult_msb_gf4_mul_2_1_n71), .Z(mult_msb_gf4_mul_2_1_n73) );
  NOR2_X1 mult_msb_gf4_mul_2_1_U23 ( .A1(mult_msb_gf4_mul_2_1_n70), .A2(
        mult_msb_gf4_mul_2_1_n69), .ZN(mult_msb_gf4_mul_2_1_n74) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U22 ( .A(InverterOutxD[10]), .B(
        InverterOutxD[11]), .ZN(mult_msb_gf4_mul_2_1_n69) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U21 ( .A(Y0_4xDP[6]), .B(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_2_1_n70) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U20 ( .A(mult_msb_gf4_mul_2_1_n68), .B(
        mult_msb_gf4_mul_2_1_n67), .ZN(mult_msb_Xi_mul_Yj_7__1_) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U19 ( .A1(InverterOutxD[9]), .A2(Y0_4xDP[5]), 
        .ZN(mult_msb_gf4_mul_2_1_n67) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U18 ( .A(mult_msb_gf4_mul_2_1_n75), .B(
        mult_msb_gf4_mul_2_1_n66), .Z(mult_msb_gf4_mul_2_1_n68) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U17 ( .A(mult_msb_gf4_mul_2_1_n65), .B(
        mult_msb_gf4_mul_2_1_n64), .ZN(mult_msb_gf4_mul_2_1_n75) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U16 ( .A1(mult_msb_gf4_mul_2_1_n63), .A2(
        mult_msb_gf4_mul_2_1_n62), .ZN(mult_msb_gf4_mul_2_1_n64) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U15 ( .A(mult_msb_gf4_mul_2_1_n61), .B(
        mult_msb_gf4_mul_2_1_n60), .ZN(mult_msb_gf4_mul_2_1_n62) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U14 ( .A(mult_msb_gf4_mul_2_1_n59), .B(
        mult_msb_gf4_mul_2_1_n58), .ZN(mult_msb_gf4_mul_2_1_n63) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U13 ( .A(mult_msb_gf4_mul_2_1_n57), .B(
        mult_msb_gf4_mul_2_1_n56), .ZN(mult_msb_Xi_mul_Yj_7__0_) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U12 ( .A1(InverterOutxD[8]), .A2(Y0_4xDP[4]), 
        .ZN(mult_msb_gf4_mul_2_1_n56) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U11 ( .A(mult_msb_gf4_mul_2_1_n66), .B(
        mult_msb_gf4_mul_2_1_n71), .Z(mult_msb_gf4_mul_2_1_n57) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U10 ( .A(mult_msb_gf4_mul_2_1_n55), .B(
        mult_msb_gf4_mul_2_1_n65), .ZN(mult_msb_gf4_mul_2_1_n71) );
  NOR2_X1 mult_msb_gf4_mul_2_1_U9 ( .A1(mult_msb_gf4_mul_2_1_n61), .A2(
        mult_msb_gf4_mul_2_1_n59), .ZN(mult_msb_gf4_mul_2_1_n65) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U8 ( .A(InverterOutxD[8]), .B(
        InverterOutxD[10]), .ZN(mult_msb_gf4_mul_2_1_n59) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U7 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_2_1_n61) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U6 ( .A1(mult_msb_gf4_mul_2_1_n58), .A2(
        mult_msb_gf4_mul_2_1_n60), .ZN(mult_msb_gf4_mul_2_1_n55) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U5 ( .A(Y0_4xDP[5]), .B(Y0_4xDP[7]), .Z(
        mult_msb_gf4_mul_2_1_n60) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U4 ( .A(InverterOutxD[9]), .B(InverterOutxD[11]), .Z(mult_msb_gf4_mul_2_1_n58) );
  NOR2_X1 mult_msb_gf4_mul_2_1_U3 ( .A1(mult_msb_gf4_mul_2_1_n54), .A2(
        mult_msb_gf4_mul_2_1_n53), .ZN(mult_msb_gf4_mul_2_1_n66) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U2 ( .A(InverterOutxD[8]), .B(InverterOutxD[9]), .ZN(mult_msb_gf4_mul_2_1_n53) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U1 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_2_1_n54) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U29 ( .A(mult_msb_gf4_mul_2_0_n77), .B(
        mult_msb_gf4_mul_2_0_n76), .ZN(mult_msb_Xi_mul_Yj_6__3_) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U28 ( .A1(InverterOutxD[11]), .A2(Y0_4xDP[3]), 
        .ZN(mult_msb_gf4_mul_2_0_n76) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U27 ( .A(mult_msb_gf4_mul_2_0_n75), .B(
        mult_msb_gf4_mul_2_0_n74), .Z(mult_msb_gf4_mul_2_0_n77) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U26 ( .A(mult_msb_gf4_mul_2_0_n73), .B(
        mult_msb_gf4_mul_2_0_n72), .ZN(mult_msb_Xi_mul_Yj_6__2_) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U25 ( .A1(InverterOutxD[10]), .A2(Y0_4xDP[2]), 
        .ZN(mult_msb_gf4_mul_2_0_n72) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U24 ( .A(mult_msb_gf4_mul_2_0_n74), .B(
        mult_msb_gf4_mul_2_0_n71), .Z(mult_msb_gf4_mul_2_0_n73) );
  NOR2_X1 mult_msb_gf4_mul_2_0_U23 ( .A1(mult_msb_gf4_mul_2_0_n70), .A2(
        mult_msb_gf4_mul_2_0_n69), .ZN(mult_msb_gf4_mul_2_0_n74) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U22 ( .A(InverterOutxD[10]), .B(
        InverterOutxD[11]), .ZN(mult_msb_gf4_mul_2_0_n69) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U21 ( .A(Y0_4xDP[2]), .B(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_2_0_n70) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U20 ( .A(mult_msb_gf4_mul_2_0_n68), .B(
        mult_msb_gf4_mul_2_0_n67), .ZN(mult_msb_Xi_mul_Yj_6__1_) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U19 ( .A1(InverterOutxD[9]), .A2(Y0_4xDP[1]), 
        .ZN(mult_msb_gf4_mul_2_0_n67) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U18 ( .A(mult_msb_gf4_mul_2_0_n75), .B(
        mult_msb_gf4_mul_2_0_n66), .Z(mult_msb_gf4_mul_2_0_n68) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U17 ( .A(mult_msb_gf4_mul_2_0_n65), .B(
        mult_msb_gf4_mul_2_0_n64), .ZN(mult_msb_gf4_mul_2_0_n75) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U16 ( .A1(mult_msb_gf4_mul_2_0_n63), .A2(
        mult_msb_gf4_mul_2_0_n62), .ZN(mult_msb_gf4_mul_2_0_n64) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U15 ( .A(mult_msb_gf4_mul_2_0_n61), .B(
        mult_msb_gf4_mul_2_0_n60), .ZN(mult_msb_gf4_mul_2_0_n62) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U14 ( .A(mult_msb_gf4_mul_2_0_n59), .B(
        mult_msb_gf4_mul_2_0_n58), .ZN(mult_msb_gf4_mul_2_0_n63) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U13 ( .A(mult_msb_gf4_mul_2_0_n57), .B(
        mult_msb_gf4_mul_2_0_n56), .ZN(mult_msb_Xi_mul_Yj_6__0_) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U12 ( .A1(InverterOutxD[8]), .A2(Y0_4xDP[0]), 
        .ZN(mult_msb_gf4_mul_2_0_n56) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U11 ( .A(mult_msb_gf4_mul_2_0_n66), .B(
        mult_msb_gf4_mul_2_0_n71), .Z(mult_msb_gf4_mul_2_0_n57) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U10 ( .A(mult_msb_gf4_mul_2_0_n55), .B(
        mult_msb_gf4_mul_2_0_n65), .ZN(mult_msb_gf4_mul_2_0_n71) );
  NOR2_X1 mult_msb_gf4_mul_2_0_U9 ( .A1(mult_msb_gf4_mul_2_0_n61), .A2(
        mult_msb_gf4_mul_2_0_n59), .ZN(mult_msb_gf4_mul_2_0_n65) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U8 ( .A(InverterOutxD[8]), .B(
        InverterOutxD[10]), .ZN(mult_msb_gf4_mul_2_0_n59) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U7 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_2_0_n61) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U6 ( .A1(mult_msb_gf4_mul_2_0_n58), .A2(
        mult_msb_gf4_mul_2_0_n60), .ZN(mult_msb_gf4_mul_2_0_n55) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U5 ( .A(Y0_4xDP[1]), .B(Y0_4xDP[3]), .Z(
        mult_msb_gf4_mul_2_0_n60) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U4 ( .A(InverterOutxD[9]), .B(InverterOutxD[11]), .Z(mult_msb_gf4_mul_2_0_n58) );
  NOR2_X1 mult_msb_gf4_mul_2_0_U3 ( .A1(mult_msb_gf4_mul_2_0_n54), .A2(
        mult_msb_gf4_mul_2_0_n53), .ZN(mult_msb_gf4_mul_2_0_n66) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U2 ( .A(InverterOutxD[8]), .B(InverterOutxD[9]), .ZN(mult_msb_gf4_mul_2_0_n53) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U1 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_2_0_n54) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U29 ( .A(mult_msb_gf4_mul_1_2_n77), .B(
        mult_msb_gf4_mul_1_2_n76), .ZN(mult_msb_Xi_mul_Yj_5__3_) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U28 ( .A1(InverterOutxD[7]), .A2(Y0_4xDP[11]), 
        .ZN(mult_msb_gf4_mul_1_2_n76) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U27 ( .A(mult_msb_gf4_mul_1_2_n75), .B(
        mult_msb_gf4_mul_1_2_n74), .Z(mult_msb_gf4_mul_1_2_n77) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U26 ( .A(mult_msb_gf4_mul_1_2_n73), .B(
        mult_msb_gf4_mul_1_2_n72), .ZN(mult_msb_Xi_mul_Yj_5__2_) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U25 ( .A1(InverterOutxD[6]), .A2(Y0_4xDP[10]), 
        .ZN(mult_msb_gf4_mul_1_2_n72) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U24 ( .A(mult_msb_gf4_mul_1_2_n74), .B(
        mult_msb_gf4_mul_1_2_n71), .Z(mult_msb_gf4_mul_1_2_n73) );
  NOR2_X1 mult_msb_gf4_mul_1_2_U23 ( .A1(mult_msb_gf4_mul_1_2_n70), .A2(
        mult_msb_gf4_mul_1_2_n69), .ZN(mult_msb_gf4_mul_1_2_n74) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U22 ( .A(InverterOutxD[6]), .B(
        InverterOutxD[7]), .ZN(mult_msb_gf4_mul_1_2_n69) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U21 ( .A(Y0_4xDP[10]), .B(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_1_2_n70) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U20 ( .A(mult_msb_gf4_mul_1_2_n68), .B(
        mult_msb_gf4_mul_1_2_n67), .ZN(mult_msb_Xi_mul_Yj_5__1_) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U19 ( .A1(InverterOutxD[5]), .A2(Y0_4xDP[9]), 
        .ZN(mult_msb_gf4_mul_1_2_n67) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U18 ( .A(mult_msb_gf4_mul_1_2_n75), .B(
        mult_msb_gf4_mul_1_2_n66), .Z(mult_msb_gf4_mul_1_2_n68) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U17 ( .A(mult_msb_gf4_mul_1_2_n65), .B(
        mult_msb_gf4_mul_1_2_n64), .ZN(mult_msb_gf4_mul_1_2_n75) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U16 ( .A1(mult_msb_gf4_mul_1_2_n63), .A2(
        mult_msb_gf4_mul_1_2_n62), .ZN(mult_msb_gf4_mul_1_2_n64) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U15 ( .A(mult_msb_gf4_mul_1_2_n61), .B(
        mult_msb_gf4_mul_1_2_n60), .ZN(mult_msb_gf4_mul_1_2_n62) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U14 ( .A(mult_msb_gf4_mul_1_2_n59), .B(
        mult_msb_gf4_mul_1_2_n58), .ZN(mult_msb_gf4_mul_1_2_n63) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U13 ( .A(mult_msb_gf4_mul_1_2_n57), .B(
        mult_msb_gf4_mul_1_2_n56), .ZN(mult_msb_Xi_mul_Yj_5__0_) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U12 ( .A1(InverterOutxD[4]), .A2(Y0_4xDP[8]), 
        .ZN(mult_msb_gf4_mul_1_2_n56) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U11 ( .A(mult_msb_gf4_mul_1_2_n66), .B(
        mult_msb_gf4_mul_1_2_n71), .Z(mult_msb_gf4_mul_1_2_n57) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U10 ( .A(mult_msb_gf4_mul_1_2_n55), .B(
        mult_msb_gf4_mul_1_2_n65), .ZN(mult_msb_gf4_mul_1_2_n71) );
  NOR2_X1 mult_msb_gf4_mul_1_2_U9 ( .A1(mult_msb_gf4_mul_1_2_n61), .A2(
        mult_msb_gf4_mul_1_2_n59), .ZN(mult_msb_gf4_mul_1_2_n65) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U8 ( .A(InverterOutxD[4]), .B(InverterOutxD[6]), .ZN(mult_msb_gf4_mul_1_2_n59) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U7 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_1_2_n61) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U6 ( .A1(mult_msb_gf4_mul_1_2_n58), .A2(
        mult_msb_gf4_mul_1_2_n60), .ZN(mult_msb_gf4_mul_1_2_n55) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U5 ( .A(Y0_4xDP[9]), .B(Y0_4xDP[11]), .Z(
        mult_msb_gf4_mul_1_2_n60) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U4 ( .A(InverterOutxD[5]), .B(InverterOutxD[7]), 
        .Z(mult_msb_gf4_mul_1_2_n58) );
  NOR2_X1 mult_msb_gf4_mul_1_2_U3 ( .A1(mult_msb_gf4_mul_1_2_n54), .A2(
        mult_msb_gf4_mul_1_2_n53), .ZN(mult_msb_gf4_mul_1_2_n66) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U2 ( .A(InverterOutxD[4]), .B(InverterOutxD[5]), .ZN(mult_msb_gf4_mul_1_2_n53) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U1 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_1_2_n54) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U29 ( .A(mult_msb_gf4_mul_1_1_n77), .B(
        mult_msb_gf4_mul_1_1_n76), .ZN(mult_msb_FFxDN[19]) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U28 ( .A1(InverterOutxD[7]), .A2(Y0_4xDP[7]), 
        .ZN(mult_msb_gf4_mul_1_1_n76) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U27 ( .A(mult_msb_gf4_mul_1_1_n75), .B(
        mult_msb_gf4_mul_1_1_n74), .Z(mult_msb_gf4_mul_1_1_n77) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U26 ( .A(mult_msb_gf4_mul_1_1_n73), .B(
        mult_msb_gf4_mul_1_1_n72), .ZN(mult_msb_FFxDN[18]) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U25 ( .A1(InverterOutxD[6]), .A2(Y0_4xDP[6]), 
        .ZN(mult_msb_gf4_mul_1_1_n72) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U24 ( .A(mult_msb_gf4_mul_1_1_n74), .B(
        mult_msb_gf4_mul_1_1_n71), .Z(mult_msb_gf4_mul_1_1_n73) );
  NOR2_X1 mult_msb_gf4_mul_1_1_U23 ( .A1(mult_msb_gf4_mul_1_1_n70), .A2(
        mult_msb_gf4_mul_1_1_n69), .ZN(mult_msb_gf4_mul_1_1_n74) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U22 ( .A(InverterOutxD[6]), .B(
        InverterOutxD[7]), .ZN(mult_msb_gf4_mul_1_1_n69) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U21 ( .A(Y0_4xDP[6]), .B(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_1_1_n70) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U20 ( .A(mult_msb_gf4_mul_1_1_n68), .B(
        mult_msb_gf4_mul_1_1_n67), .ZN(mult_msb_FFxDN[17]) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U19 ( .A1(InverterOutxD[5]), .A2(Y0_4xDP[5]), 
        .ZN(mult_msb_gf4_mul_1_1_n67) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U18 ( .A(mult_msb_gf4_mul_1_1_n75), .B(
        mult_msb_gf4_mul_1_1_n66), .Z(mult_msb_gf4_mul_1_1_n68) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U17 ( .A(mult_msb_gf4_mul_1_1_n65), .B(
        mult_msb_gf4_mul_1_1_n64), .ZN(mult_msb_gf4_mul_1_1_n75) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U16 ( .A1(mult_msb_gf4_mul_1_1_n63), .A2(
        mult_msb_gf4_mul_1_1_n62), .ZN(mult_msb_gf4_mul_1_1_n64) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U15 ( .A(mult_msb_gf4_mul_1_1_n61), .B(
        mult_msb_gf4_mul_1_1_n60), .ZN(mult_msb_gf4_mul_1_1_n62) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U14 ( .A(mult_msb_gf4_mul_1_1_n59), .B(
        mult_msb_gf4_mul_1_1_n58), .ZN(mult_msb_gf4_mul_1_1_n63) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U13 ( .A(mult_msb_gf4_mul_1_1_n57), .B(
        mult_msb_gf4_mul_1_1_n56), .ZN(mult_msb_FFxDN[16]) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U12 ( .A1(InverterOutxD[4]), .A2(Y0_4xDP[4]), 
        .ZN(mult_msb_gf4_mul_1_1_n56) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U11 ( .A(mult_msb_gf4_mul_1_1_n66), .B(
        mult_msb_gf4_mul_1_1_n71), .Z(mult_msb_gf4_mul_1_1_n57) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U10 ( .A(mult_msb_gf4_mul_1_1_n55), .B(
        mult_msb_gf4_mul_1_1_n65), .ZN(mult_msb_gf4_mul_1_1_n71) );
  NOR2_X1 mult_msb_gf4_mul_1_1_U9 ( .A1(mult_msb_gf4_mul_1_1_n61), .A2(
        mult_msb_gf4_mul_1_1_n59), .ZN(mult_msb_gf4_mul_1_1_n65) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U8 ( .A(InverterOutxD[4]), .B(InverterOutxD[6]), .ZN(mult_msb_gf4_mul_1_1_n59) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U7 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_1_1_n61) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U6 ( .A1(mult_msb_gf4_mul_1_1_n58), .A2(
        mult_msb_gf4_mul_1_1_n60), .ZN(mult_msb_gf4_mul_1_1_n55) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U5 ( .A(Y0_4xDP[5]), .B(Y0_4xDP[7]), .Z(
        mult_msb_gf4_mul_1_1_n60) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U4 ( .A(InverterOutxD[5]), .B(InverterOutxD[7]), 
        .Z(mult_msb_gf4_mul_1_1_n58) );
  NOR2_X1 mult_msb_gf4_mul_1_1_U3 ( .A1(mult_msb_gf4_mul_1_1_n54), .A2(
        mult_msb_gf4_mul_1_1_n53), .ZN(mult_msb_gf4_mul_1_1_n66) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U2 ( .A(InverterOutxD[4]), .B(InverterOutxD[5]), .ZN(mult_msb_gf4_mul_1_1_n53) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U1 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_1_1_n54) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U29 ( .A(mult_msb_gf4_mul_1_0_n77), .B(
        mult_msb_gf4_mul_1_0_n76), .ZN(mult_msb_Xi_mul_Yj_3__3_) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U28 ( .A1(InverterOutxD[7]), .A2(Y0_4xDP[3]), 
        .ZN(mult_msb_gf4_mul_1_0_n76) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U27 ( .A(mult_msb_gf4_mul_1_0_n75), .B(
        mult_msb_gf4_mul_1_0_n74), .Z(mult_msb_gf4_mul_1_0_n77) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U26 ( .A(mult_msb_gf4_mul_1_0_n73), .B(
        mult_msb_gf4_mul_1_0_n72), .ZN(mult_msb_Xi_mul_Yj_3__2_) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U25 ( .A1(InverterOutxD[6]), .A2(Y0_4xDP[2]), 
        .ZN(mult_msb_gf4_mul_1_0_n72) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U24 ( .A(mult_msb_gf4_mul_1_0_n74), .B(
        mult_msb_gf4_mul_1_0_n71), .Z(mult_msb_gf4_mul_1_0_n73) );
  NOR2_X1 mult_msb_gf4_mul_1_0_U23 ( .A1(mult_msb_gf4_mul_1_0_n70), .A2(
        mult_msb_gf4_mul_1_0_n69), .ZN(mult_msb_gf4_mul_1_0_n74) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U22 ( .A(InverterOutxD[6]), .B(
        InverterOutxD[7]), .ZN(mult_msb_gf4_mul_1_0_n69) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U21 ( .A(Y0_4xDP[2]), .B(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_1_0_n70) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U20 ( .A(mult_msb_gf4_mul_1_0_n68), .B(
        mult_msb_gf4_mul_1_0_n67), .ZN(mult_msb_Xi_mul_Yj_3__1_) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U19 ( .A1(InverterOutxD[5]), .A2(Y0_4xDP[1]), 
        .ZN(mult_msb_gf4_mul_1_0_n67) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U18 ( .A(mult_msb_gf4_mul_1_0_n75), .B(
        mult_msb_gf4_mul_1_0_n66), .Z(mult_msb_gf4_mul_1_0_n68) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U17 ( .A(mult_msb_gf4_mul_1_0_n65), .B(
        mult_msb_gf4_mul_1_0_n64), .ZN(mult_msb_gf4_mul_1_0_n75) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U16 ( .A1(mult_msb_gf4_mul_1_0_n63), .A2(
        mult_msb_gf4_mul_1_0_n62), .ZN(mult_msb_gf4_mul_1_0_n64) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U15 ( .A(mult_msb_gf4_mul_1_0_n61), .B(
        mult_msb_gf4_mul_1_0_n60), .ZN(mult_msb_gf4_mul_1_0_n62) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U14 ( .A(mult_msb_gf4_mul_1_0_n59), .B(
        mult_msb_gf4_mul_1_0_n58), .ZN(mult_msb_gf4_mul_1_0_n63) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U13 ( .A(mult_msb_gf4_mul_1_0_n57), .B(
        mult_msb_gf4_mul_1_0_n56), .ZN(mult_msb_Xi_mul_Yj_3__0_) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U12 ( .A1(InverterOutxD[4]), .A2(Y0_4xDP[0]), 
        .ZN(mult_msb_gf4_mul_1_0_n56) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U11 ( .A(mult_msb_gf4_mul_1_0_n66), .B(
        mult_msb_gf4_mul_1_0_n71), .Z(mult_msb_gf4_mul_1_0_n57) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U10 ( .A(mult_msb_gf4_mul_1_0_n55), .B(
        mult_msb_gf4_mul_1_0_n65), .ZN(mult_msb_gf4_mul_1_0_n71) );
  NOR2_X1 mult_msb_gf4_mul_1_0_U9 ( .A1(mult_msb_gf4_mul_1_0_n61), .A2(
        mult_msb_gf4_mul_1_0_n59), .ZN(mult_msb_gf4_mul_1_0_n65) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U8 ( .A(InverterOutxD[4]), .B(InverterOutxD[6]), .ZN(mult_msb_gf4_mul_1_0_n59) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U7 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_1_0_n61) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U6 ( .A1(mult_msb_gf4_mul_1_0_n58), .A2(
        mult_msb_gf4_mul_1_0_n60), .ZN(mult_msb_gf4_mul_1_0_n55) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U5 ( .A(Y0_4xDP[1]), .B(Y0_4xDP[3]), .Z(
        mult_msb_gf4_mul_1_0_n60) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U4 ( .A(InverterOutxD[5]), .B(InverterOutxD[7]), 
        .Z(mult_msb_gf4_mul_1_0_n58) );
  NOR2_X1 mult_msb_gf4_mul_1_0_U3 ( .A1(mult_msb_gf4_mul_1_0_n54), .A2(
        mult_msb_gf4_mul_1_0_n53), .ZN(mult_msb_gf4_mul_1_0_n66) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U2 ( .A(InverterOutxD[4]), .B(InverterOutxD[5]), .ZN(mult_msb_gf4_mul_1_0_n53) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U1 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_1_0_n54) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U29 ( .A(mult_msb_gf4_mul_0_2_n77), .B(
        mult_msb_gf4_mul_0_2_n76), .ZN(mult_msb_Xi_mul_Yj_2__3_) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U28 ( .A1(InverterOutxD[3]), .A2(Y0_4xDP[11]), 
        .ZN(mult_msb_gf4_mul_0_2_n76) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U27 ( .A(mult_msb_gf4_mul_0_2_n75), .B(
        mult_msb_gf4_mul_0_2_n74), .Z(mult_msb_gf4_mul_0_2_n77) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U26 ( .A(mult_msb_gf4_mul_0_2_n73), .B(
        mult_msb_gf4_mul_0_2_n72), .ZN(mult_msb_Xi_mul_Yj_2__2_) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U25 ( .A1(InverterOutxD[2]), .A2(Y0_4xDP[10]), 
        .ZN(mult_msb_gf4_mul_0_2_n72) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U24 ( .A(mult_msb_gf4_mul_0_2_n74), .B(
        mult_msb_gf4_mul_0_2_n71), .Z(mult_msb_gf4_mul_0_2_n73) );
  NOR2_X1 mult_msb_gf4_mul_0_2_U23 ( .A1(mult_msb_gf4_mul_0_2_n70), .A2(
        mult_msb_gf4_mul_0_2_n69), .ZN(mult_msb_gf4_mul_0_2_n74) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U22 ( .A(InverterOutxD[2]), .B(
        InverterOutxD[3]), .ZN(mult_msb_gf4_mul_0_2_n69) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U21 ( .A(Y0_4xDP[10]), .B(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_0_2_n70) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U20 ( .A(mult_msb_gf4_mul_0_2_n68), .B(
        mult_msb_gf4_mul_0_2_n67), .ZN(mult_msb_Xi_mul_Yj_2__1_) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U19 ( .A1(InverterOutxD[1]), .A2(Y0_4xDP[9]), 
        .ZN(mult_msb_gf4_mul_0_2_n67) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U18 ( .A(mult_msb_gf4_mul_0_2_n75), .B(
        mult_msb_gf4_mul_0_2_n66), .Z(mult_msb_gf4_mul_0_2_n68) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U17 ( .A(mult_msb_gf4_mul_0_2_n65), .B(
        mult_msb_gf4_mul_0_2_n64), .ZN(mult_msb_gf4_mul_0_2_n75) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U16 ( .A1(mult_msb_gf4_mul_0_2_n63), .A2(
        mult_msb_gf4_mul_0_2_n62), .ZN(mult_msb_gf4_mul_0_2_n64) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U15 ( .A(mult_msb_gf4_mul_0_2_n61), .B(
        mult_msb_gf4_mul_0_2_n60), .ZN(mult_msb_gf4_mul_0_2_n62) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U14 ( .A(mult_msb_gf4_mul_0_2_n59), .B(
        mult_msb_gf4_mul_0_2_n58), .ZN(mult_msb_gf4_mul_0_2_n63) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U13 ( .A(mult_msb_gf4_mul_0_2_n57), .B(
        mult_msb_gf4_mul_0_2_n56), .ZN(mult_msb_Xi_mul_Yj_2__0_) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U12 ( .A1(InverterOutxD[0]), .A2(Y0_4xDP[8]), 
        .ZN(mult_msb_gf4_mul_0_2_n56) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U11 ( .A(mult_msb_gf4_mul_0_2_n66), .B(
        mult_msb_gf4_mul_0_2_n71), .Z(mult_msb_gf4_mul_0_2_n57) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U10 ( .A(mult_msb_gf4_mul_0_2_n55), .B(
        mult_msb_gf4_mul_0_2_n65), .ZN(mult_msb_gf4_mul_0_2_n71) );
  NOR2_X1 mult_msb_gf4_mul_0_2_U9 ( .A1(mult_msb_gf4_mul_0_2_n61), .A2(
        mult_msb_gf4_mul_0_2_n59), .ZN(mult_msb_gf4_mul_0_2_n65) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U8 ( .A(InverterOutxD[0]), .B(InverterOutxD[2]), .ZN(mult_msb_gf4_mul_0_2_n59) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U7 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_0_2_n61) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U6 ( .A1(mult_msb_gf4_mul_0_2_n58), .A2(
        mult_msb_gf4_mul_0_2_n60), .ZN(mult_msb_gf4_mul_0_2_n55) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U5 ( .A(Y0_4xDP[9]), .B(Y0_4xDP[11]), .Z(
        mult_msb_gf4_mul_0_2_n60) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U4 ( .A(InverterOutxD[1]), .B(InverterOutxD[3]), 
        .Z(mult_msb_gf4_mul_0_2_n58) );
  NOR2_X1 mult_msb_gf4_mul_0_2_U3 ( .A1(mult_msb_gf4_mul_0_2_n54), .A2(
        mult_msb_gf4_mul_0_2_n53), .ZN(mult_msb_gf4_mul_0_2_n66) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U2 ( .A(InverterOutxD[0]), .B(InverterOutxD[1]), .ZN(mult_msb_gf4_mul_0_2_n53) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U1 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_0_2_n54) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U29 ( .A(mult_msb_gf4_mul_0_1_n77), .B(
        mult_msb_gf4_mul_0_1_n76), .ZN(mult_msb_Xi_mul_Yj_1__3_) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U28 ( .A1(InverterOutxD[3]), .A2(Y0_4xDP[7]), 
        .ZN(mult_msb_gf4_mul_0_1_n76) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U27 ( .A(mult_msb_gf4_mul_0_1_n75), .B(
        mult_msb_gf4_mul_0_1_n74), .Z(mult_msb_gf4_mul_0_1_n77) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U26 ( .A(mult_msb_gf4_mul_0_1_n73), .B(
        mult_msb_gf4_mul_0_1_n72), .ZN(mult_msb_Xi_mul_Yj_1__2_) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U25 ( .A1(InverterOutxD[2]), .A2(Y0_4xDP[6]), 
        .ZN(mult_msb_gf4_mul_0_1_n72) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U24 ( .A(mult_msb_gf4_mul_0_1_n74), .B(
        mult_msb_gf4_mul_0_1_n71), .Z(mult_msb_gf4_mul_0_1_n73) );
  NOR2_X1 mult_msb_gf4_mul_0_1_U23 ( .A1(mult_msb_gf4_mul_0_1_n70), .A2(
        mult_msb_gf4_mul_0_1_n69), .ZN(mult_msb_gf4_mul_0_1_n74) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U22 ( .A(InverterOutxD[2]), .B(
        InverterOutxD[3]), .ZN(mult_msb_gf4_mul_0_1_n69) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U21 ( .A(Y0_4xDP[6]), .B(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_0_1_n70) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U20 ( .A(mult_msb_gf4_mul_0_1_n68), .B(
        mult_msb_gf4_mul_0_1_n67), .ZN(mult_msb_Xi_mul_Yj_1__1_) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U19 ( .A1(InverterOutxD[1]), .A2(Y0_4xDP[5]), 
        .ZN(mult_msb_gf4_mul_0_1_n67) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U18 ( .A(mult_msb_gf4_mul_0_1_n75), .B(
        mult_msb_gf4_mul_0_1_n66), .Z(mult_msb_gf4_mul_0_1_n68) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U17 ( .A(mult_msb_gf4_mul_0_1_n65), .B(
        mult_msb_gf4_mul_0_1_n64), .ZN(mult_msb_gf4_mul_0_1_n75) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U16 ( .A1(mult_msb_gf4_mul_0_1_n63), .A2(
        mult_msb_gf4_mul_0_1_n62), .ZN(mult_msb_gf4_mul_0_1_n64) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U15 ( .A(mult_msb_gf4_mul_0_1_n61), .B(
        mult_msb_gf4_mul_0_1_n60), .ZN(mult_msb_gf4_mul_0_1_n62) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U14 ( .A(mult_msb_gf4_mul_0_1_n59), .B(
        mult_msb_gf4_mul_0_1_n58), .ZN(mult_msb_gf4_mul_0_1_n63) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U13 ( .A(mult_msb_gf4_mul_0_1_n57), .B(
        mult_msb_gf4_mul_0_1_n56), .ZN(mult_msb_Xi_mul_Yj_1__0_) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U12 ( .A1(InverterOutxD[0]), .A2(Y0_4xDP[4]), 
        .ZN(mult_msb_gf4_mul_0_1_n56) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U11 ( .A(mult_msb_gf4_mul_0_1_n66), .B(
        mult_msb_gf4_mul_0_1_n71), .Z(mult_msb_gf4_mul_0_1_n57) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U10 ( .A(mult_msb_gf4_mul_0_1_n55), .B(
        mult_msb_gf4_mul_0_1_n65), .ZN(mult_msb_gf4_mul_0_1_n71) );
  NOR2_X1 mult_msb_gf4_mul_0_1_U9 ( .A1(mult_msb_gf4_mul_0_1_n61), .A2(
        mult_msb_gf4_mul_0_1_n59), .ZN(mult_msb_gf4_mul_0_1_n65) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U8 ( .A(InverterOutxD[0]), .B(InverterOutxD[2]), .ZN(mult_msb_gf4_mul_0_1_n59) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U7 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_0_1_n61) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U6 ( .A1(mult_msb_gf4_mul_0_1_n58), .A2(
        mult_msb_gf4_mul_0_1_n60), .ZN(mult_msb_gf4_mul_0_1_n55) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U5 ( .A(Y0_4xDP[5]), .B(Y0_4xDP[7]), .Z(
        mult_msb_gf4_mul_0_1_n60) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U4 ( .A(InverterOutxD[1]), .B(InverterOutxD[3]), 
        .Z(mult_msb_gf4_mul_0_1_n58) );
  NOR2_X1 mult_msb_gf4_mul_0_1_U3 ( .A1(mult_msb_gf4_mul_0_1_n54), .A2(
        mult_msb_gf4_mul_0_1_n53), .ZN(mult_msb_gf4_mul_0_1_n66) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U2 ( .A(InverterOutxD[0]), .B(InverterOutxD[1]), .ZN(mult_msb_gf4_mul_0_1_n53) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U1 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_0_1_n54) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U29 ( .A(mult_msb_gf4_mul_0_0_n77), .B(
        mult_msb_gf4_mul_0_0_n76), .ZN(mult_msb_FFxDN[3]) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U28 ( .A1(InverterOutxD[3]), .A2(Y0_4xDP[3]), 
        .ZN(mult_msb_gf4_mul_0_0_n76) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U27 ( .A(mult_msb_gf4_mul_0_0_n75), .B(
        mult_msb_gf4_mul_0_0_n74), .Z(mult_msb_gf4_mul_0_0_n77) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U26 ( .A(mult_msb_gf4_mul_0_0_n73), .B(
        mult_msb_gf4_mul_0_0_n72), .ZN(mult_msb_FFxDN[2]) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U25 ( .A1(InverterOutxD[2]), .A2(Y0_4xDP[2]), 
        .ZN(mult_msb_gf4_mul_0_0_n72) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U24 ( .A(mult_msb_gf4_mul_0_0_n74), .B(
        mult_msb_gf4_mul_0_0_n71), .Z(mult_msb_gf4_mul_0_0_n73) );
  NOR2_X1 mult_msb_gf4_mul_0_0_U23 ( .A1(mult_msb_gf4_mul_0_0_n70), .A2(
        mult_msb_gf4_mul_0_0_n69), .ZN(mult_msb_gf4_mul_0_0_n74) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U22 ( .A(InverterOutxD[2]), .B(
        InverterOutxD[3]), .ZN(mult_msb_gf4_mul_0_0_n69) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U21 ( .A(Y0_4xDP[2]), .B(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_0_0_n70) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U20 ( .A(mult_msb_gf4_mul_0_0_n68), .B(
        mult_msb_gf4_mul_0_0_n67), .ZN(mult_msb_FFxDN[1]) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U19 ( .A1(InverterOutxD[1]), .A2(Y0_4xDP[1]), 
        .ZN(mult_msb_gf4_mul_0_0_n67) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U18 ( .A(mult_msb_gf4_mul_0_0_n75), .B(
        mult_msb_gf4_mul_0_0_n66), .Z(mult_msb_gf4_mul_0_0_n68) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U17 ( .A(mult_msb_gf4_mul_0_0_n65), .B(
        mult_msb_gf4_mul_0_0_n64), .ZN(mult_msb_gf4_mul_0_0_n75) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U16 ( .A1(mult_msb_gf4_mul_0_0_n63), .A2(
        mult_msb_gf4_mul_0_0_n62), .ZN(mult_msb_gf4_mul_0_0_n64) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U15 ( .A(mult_msb_gf4_mul_0_0_n61), .B(
        mult_msb_gf4_mul_0_0_n60), .ZN(mult_msb_gf4_mul_0_0_n62) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U14 ( .A(mult_msb_gf4_mul_0_0_n59), .B(
        mult_msb_gf4_mul_0_0_n58), .ZN(mult_msb_gf4_mul_0_0_n63) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U13 ( .A(mult_msb_gf4_mul_0_0_n57), .B(
        mult_msb_gf4_mul_0_0_n56), .ZN(mult_msb_FFxDN[0]) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U12 ( .A1(InverterOutxD[0]), .A2(Y0_4xDP[0]), 
        .ZN(mult_msb_gf4_mul_0_0_n56) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U11 ( .A(mult_msb_gf4_mul_0_0_n66), .B(
        mult_msb_gf4_mul_0_0_n71), .Z(mult_msb_gf4_mul_0_0_n57) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U10 ( .A(mult_msb_gf4_mul_0_0_n55), .B(
        mult_msb_gf4_mul_0_0_n65), .ZN(mult_msb_gf4_mul_0_0_n71) );
  NOR2_X1 mult_msb_gf4_mul_0_0_U9 ( .A1(mult_msb_gf4_mul_0_0_n61), .A2(
        mult_msb_gf4_mul_0_0_n59), .ZN(mult_msb_gf4_mul_0_0_n65) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U8 ( .A(InverterOutxD[0]), .B(InverterOutxD[2]), .ZN(mult_msb_gf4_mul_0_0_n59) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U7 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_0_0_n61) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U6 ( .A1(mult_msb_gf4_mul_0_0_n58), .A2(
        mult_msb_gf4_mul_0_0_n60), .ZN(mult_msb_gf4_mul_0_0_n55) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U5 ( .A(Y0_4xDP[1]), .B(Y0_4xDP[3]), .Z(
        mult_msb_gf4_mul_0_0_n60) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U4 ( .A(InverterOutxD[1]), .B(InverterOutxD[3]), 
        .Z(mult_msb_gf4_mul_0_0_n58) );
  NOR2_X1 mult_msb_gf4_mul_0_0_U3 ( .A1(mult_msb_gf4_mul_0_0_n54), .A2(
        mult_msb_gf4_mul_0_0_n53), .ZN(mult_msb_gf4_mul_0_0_n66) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U2 ( .A(InverterOutxD[0]), .B(InverterOutxD[1]), .ZN(mult_msb_gf4_mul_0_0_n53) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U1 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_0_0_n54) );
  XNOR2_X1 mult_lsb_U50 ( .A(mult_lsb_n96), .B(mult_lsb_n60), .ZN(
        InvUnmappedxD[19]) );
  XOR2_X1 mult_lsb_U49 ( .A(mult_lsb_n94), .B(mult_lsb_n95), .Z(mult_lsb_n60)
         );
  XNOR2_X1 mult_lsb_U48 ( .A(mult_lsb_n93), .B(mult_lsb_n59), .ZN(
        InvUnmappedxD[18]) );
  XOR2_X1 mult_lsb_U47 ( .A(mult_lsb_n91), .B(mult_lsb_n92), .Z(mult_lsb_n59)
         );
  XNOR2_X1 mult_lsb_U46 ( .A(mult_lsb_n90), .B(mult_lsb_n58), .ZN(
        InvUnmappedxD[17]) );
  XOR2_X1 mult_lsb_U45 ( .A(mult_lsb_n88), .B(mult_lsb_n89), .Z(mult_lsb_n58)
         );
  XNOR2_X1 mult_lsb_U44 ( .A(mult_lsb_n87), .B(mult_lsb_n57), .ZN(
        InvUnmappedxD[16]) );
  XOR2_X1 mult_lsb_U43 ( .A(mult_lsb_n85), .B(mult_lsb_n86), .Z(mult_lsb_n57)
         );
  XNOR2_X1 mult_lsb_U42 ( .A(mult_lsb_n84), .B(mult_lsb_n56), .ZN(
        InvUnmappedxD[11]) );
  XOR2_X1 mult_lsb_U41 ( .A(mult_lsb_n82), .B(mult_lsb_n83), .Z(mult_lsb_n56)
         );
  XNOR2_X1 mult_lsb_U40 ( .A(mult_lsb_n81), .B(mult_lsb_n55), .ZN(
        InvUnmappedxD[10]) );
  XOR2_X1 mult_lsb_U39 ( .A(mult_lsb_n79), .B(mult_lsb_n80), .Z(mult_lsb_n55)
         );
  XNOR2_X1 mult_lsb_U38 ( .A(mult_lsb_n78), .B(mult_lsb_n54), .ZN(
        InvUnmappedxD[9]) );
  XOR2_X1 mult_lsb_U37 ( .A(mult_lsb_n76), .B(mult_lsb_n77), .Z(mult_lsb_n54)
         );
  XNOR2_X1 mult_lsb_U36 ( .A(mult_lsb_n75), .B(mult_lsb_n53), .ZN(
        InvUnmappedxD[8]) );
  XOR2_X1 mult_lsb_U35 ( .A(mult_lsb_n73), .B(mult_lsb_n74), .Z(mult_lsb_n53)
         );
  XNOR2_X1 mult_lsb_U34 ( .A(mult_lsb_n72), .B(mult_lsb_n52), .ZN(
        InvUnmappedxD[3]) );
  XOR2_X1 mult_lsb_U33 ( .A(mult_lsb_n70), .B(mult_lsb_n71), .Z(mult_lsb_n52)
         );
  XNOR2_X1 mult_lsb_U32 ( .A(mult_lsb_n69), .B(mult_lsb_n51), .ZN(
        InvUnmappedxD[2]) );
  XOR2_X1 mult_lsb_U31 ( .A(mult_lsb_n67), .B(mult_lsb_n68), .Z(mult_lsb_n51)
         );
  XNOR2_X1 mult_lsb_U30 ( .A(mult_lsb_n66), .B(mult_lsb_n50), .ZN(
        InvUnmappedxD[1]) );
  XOR2_X1 mult_lsb_U29 ( .A(mult_lsb_n64), .B(mult_lsb_n65), .Z(mult_lsb_n50)
         );
  XNOR2_X1 mult_lsb_U28 ( .A(mult_lsb_n63), .B(mult_lsb_n49), .ZN(
        InvUnmappedxD[0]) );
  XOR2_X1 mult_lsb_U27 ( .A(mult_lsb_n61), .B(mult_lsb_n62), .Z(mult_lsb_n49)
         );
  XOR2_X1 mult_lsb_U26 ( .A(Zmul3xDI[11]), .B(mult_lsb_Xi_mul_Yj_7__3_), .Z(
        mult_lsb_FFxDN[31]) );
  XOR2_X1 mult_lsb_U25 ( .A(Zmul3xDI[10]), .B(mult_lsb_Xi_mul_Yj_7__2_), .Z(
        mult_lsb_FFxDN[30]) );
  XOR2_X1 mult_lsb_U24 ( .A(Zmul3xDI[9]), .B(mult_lsb_Xi_mul_Yj_7__1_), .Z(
        mult_lsb_FFxDN[29]) );
  XOR2_X1 mult_lsb_U23 ( .A(Zmul3xDI[8]), .B(mult_lsb_Xi_mul_Yj_7__0_), .Z(
        mult_lsb_FFxDN[28]) );
  XOR2_X1 mult_lsb_U22 ( .A(Zmul3xDI[7]), .B(mult_lsb_Xi_mul_Yj_6__3_), .Z(
        mult_lsb_FFxDN[27]) );
  XOR2_X1 mult_lsb_U21 ( .A(Zmul3xDI[6]), .B(mult_lsb_Xi_mul_Yj_6__2_), .Z(
        mult_lsb_FFxDN[26]) );
  XOR2_X1 mult_lsb_U20 ( .A(Zmul3xDI[5]), .B(mult_lsb_Xi_mul_Yj_6__1_), .Z(
        mult_lsb_FFxDN[25]) );
  XOR2_X1 mult_lsb_U19 ( .A(Zmul3xDI[4]), .B(mult_lsb_Xi_mul_Yj_6__0_), .Z(
        mult_lsb_FFxDN[24]) );
  XOR2_X1 mult_lsb_U18 ( .A(Zmul3xDI[11]), .B(mult_lsb_Xi_mul_Yj_5__3_), .Z(
        mult_lsb_FFxDN[23]) );
  XOR2_X1 mult_lsb_U17 ( .A(Zmul3xDI[10]), .B(mult_lsb_Xi_mul_Yj_5__2_), .Z(
        mult_lsb_FFxDN[22]) );
  XOR2_X1 mult_lsb_U16 ( .A(Zmul3xDI[9]), .B(mult_lsb_Xi_mul_Yj_5__1_), .Z(
        mult_lsb_FFxDN[21]) );
  XOR2_X1 mult_lsb_U15 ( .A(Zmul3xDI[8]), .B(mult_lsb_Xi_mul_Yj_5__0_), .Z(
        mult_lsb_FFxDN[20]) );
  XOR2_X1 mult_lsb_U14 ( .A(Zmul3xDI[3]), .B(mult_lsb_Xi_mul_Yj_3__3_), .Z(
        mult_lsb_FFxDN[15]) );
  XOR2_X1 mult_lsb_U13 ( .A(Zmul3xDI[2]), .B(mult_lsb_Xi_mul_Yj_3__2_), .Z(
        mult_lsb_FFxDN[14]) );
  XOR2_X1 mult_lsb_U12 ( .A(Zmul3xDI[1]), .B(mult_lsb_Xi_mul_Yj_3__1_), .Z(
        mult_lsb_FFxDN[13]) );
  XOR2_X1 mult_lsb_U11 ( .A(Zmul3xDI[0]), .B(mult_lsb_Xi_mul_Yj_3__0_), .Z(
        mult_lsb_FFxDN[12]) );
  XOR2_X1 mult_lsb_U10 ( .A(Zmul3xDI[7]), .B(mult_lsb_Xi_mul_Yj_2__3_), .Z(
        mult_lsb_FFxDN[11]) );
  XOR2_X1 mult_lsb_U9 ( .A(Zmul3xDI[6]), .B(mult_lsb_Xi_mul_Yj_2__2_), .Z(
        mult_lsb_FFxDN[10]) );
  XOR2_X1 mult_lsb_U8 ( .A(Zmul3xDI[5]), .B(mult_lsb_Xi_mul_Yj_2__1_), .Z(
        mult_lsb_FFxDN[9]) );
  XOR2_X1 mult_lsb_U7 ( .A(Zmul3xDI[4]), .B(mult_lsb_Xi_mul_Yj_2__0_), .Z(
        mult_lsb_FFxDN[8]) );
  XOR2_X1 mult_lsb_U6 ( .A(Zmul3xDI[3]), .B(mult_lsb_Xi_mul_Yj_1__3_), .Z(
        mult_lsb_FFxDN[7]) );
  XOR2_X1 mult_lsb_U5 ( .A(Zmul3xDI[2]), .B(mult_lsb_Xi_mul_Yj_1__2_), .Z(
        mult_lsb_FFxDN[6]) );
  XOR2_X1 mult_lsb_U4 ( .A(Zmul3xDI[1]), .B(mult_lsb_Xi_mul_Yj_1__1_), .Z(
        mult_lsb_FFxDN[5]) );
  XOR2_X1 mult_lsb_U3 ( .A(Zmul3xDI[0]), .B(mult_lsb_Xi_mul_Yj_1__0_), .Z(
        mult_lsb_FFxDN[4]) );
  DFF_X1 mult_lsb_FFxDP_reg_1__3_ ( .D(mult_lsb_FFxDN[7]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n71) );
  DFF_X1 mult_lsb_FFxDP_reg_2__3_ ( .D(mult_lsb_FFxDN[11]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n70) );
  DFF_X1 mult_lsb_FFxDP_reg_3__3_ ( .D(mult_lsb_FFxDN[15]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n84) );
  DFF_X1 mult_lsb_FFxDP_reg_5__3_ ( .D(mult_lsb_FFxDN[23]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n82) );
  DFF_X1 mult_lsb_FFxDP_reg_6__3_ ( .D(mult_lsb_FFxDN[27]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n96) );
  DFF_X1 mult_lsb_FFxDP_reg_7__3_ ( .D(mult_lsb_FFxDN[31]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n95) );
  DFF_X1 mult_lsb_FFxDP_reg_1__1_ ( .D(mult_lsb_FFxDN[5]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n65) );
  DFF_X1 mult_lsb_FFxDP_reg_2__1_ ( .D(mult_lsb_FFxDN[9]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n64) );
  DFF_X1 mult_lsb_FFxDP_reg_3__1_ ( .D(mult_lsb_FFxDN[13]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n78) );
  DFF_X1 mult_lsb_FFxDP_reg_5__1_ ( .D(mult_lsb_FFxDN[21]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n76) );
  DFF_X1 mult_lsb_FFxDP_reg_6__1_ ( .D(mult_lsb_FFxDN[25]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n90) );
  DFF_X1 mult_lsb_FFxDP_reg_7__1_ ( .D(mult_lsb_FFxDN[29]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n89) );
  DFF_X1 mult_lsb_FFxDP_reg_1__2_ ( .D(mult_lsb_FFxDN[6]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n68) );
  DFF_X1 mult_lsb_FFxDP_reg_2__2_ ( .D(mult_lsb_FFxDN[10]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n67) );
  DFF_X1 mult_lsb_FFxDP_reg_3__2_ ( .D(mult_lsb_FFxDN[14]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n81) );
  DFF_X1 mult_lsb_FFxDP_reg_5__2_ ( .D(mult_lsb_FFxDN[22]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n79) );
  DFF_X1 mult_lsb_FFxDP_reg_6__2_ ( .D(mult_lsb_FFxDN[26]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n93) );
  DFF_X1 mult_lsb_FFxDP_reg_7__2_ ( .D(mult_lsb_FFxDN[30]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n92) );
  DFF_X1 mult_lsb_FFxDP_reg_1__0_ ( .D(mult_lsb_FFxDN[4]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n62) );
  DFF_X1 mult_lsb_FFxDP_reg_2__0_ ( .D(mult_lsb_FFxDN[8]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n61) );
  DFF_X1 mult_lsb_FFxDP_reg_3__0_ ( .D(mult_lsb_FFxDN[12]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n75) );
  DFF_X1 mult_lsb_FFxDP_reg_5__0_ ( .D(mult_lsb_FFxDN[20]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n73) );
  DFF_X1 mult_lsb_FFxDP_reg_6__0_ ( .D(mult_lsb_FFxDN[24]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n87) );
  DFF_X1 mult_lsb_FFxDP_reg_7__0_ ( .D(mult_lsb_FFxDN[28]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n86) );
  DFF_X1 mult_lsb_FFxDP_reg_0__3_ ( .D(mult_lsb_FFxDN[3]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n72) );
  DFF_X1 mult_lsb_FFxDP_reg_4__3_ ( .D(mult_lsb_FFxDN[19]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n83) );
  DFF_X1 mult_lsb_FFxDP_reg_8__3_ ( .D(mult_lsb_FFxDN[35]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n94) );
  DFF_X1 mult_lsb_FFxDP_reg_0__1_ ( .D(mult_lsb_FFxDN[1]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n66) );
  DFF_X1 mult_lsb_FFxDP_reg_4__1_ ( .D(mult_lsb_FFxDN[17]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n77) );
  DFF_X1 mult_lsb_FFxDP_reg_8__1_ ( .D(mult_lsb_FFxDN[33]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n88) );
  DFF_X1 mult_lsb_FFxDP_reg_0__2_ ( .D(mult_lsb_FFxDN[2]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n69) );
  DFF_X1 mult_lsb_FFxDP_reg_4__2_ ( .D(mult_lsb_FFxDN[18]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n80) );
  DFF_X1 mult_lsb_FFxDP_reg_8__2_ ( .D(mult_lsb_FFxDN[34]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n91) );
  DFF_X1 mult_lsb_FFxDP_reg_0__0_ ( .D(mult_lsb_FFxDN[0]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n63) );
  DFF_X1 mult_lsb_FFxDP_reg_4__0_ ( .D(mult_lsb_FFxDN[16]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n74) );
  DFF_X1 mult_lsb_FFxDP_reg_8__0_ ( .D(mult_lsb_FFxDN[32]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n85) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U29 ( .A(mult_lsb_gf4_mul_2_2_n77), .B(
        mult_lsb_gf4_mul_2_2_n76), .ZN(mult_lsb_FFxDN[35]) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U28 ( .A1(InverterOutxD[11]), .A2(Y1_4xDP[11]), 
        .ZN(mult_lsb_gf4_mul_2_2_n76) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U27 ( .A(mult_lsb_gf4_mul_2_2_n75), .B(
        mult_lsb_gf4_mul_2_2_n74), .Z(mult_lsb_gf4_mul_2_2_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U26 ( .A(mult_lsb_gf4_mul_2_2_n73), .B(
        mult_lsb_gf4_mul_2_2_n72), .ZN(mult_lsb_FFxDN[34]) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U25 ( .A1(InverterOutxD[10]), .A2(Y1_4xDP[10]), 
        .ZN(mult_lsb_gf4_mul_2_2_n72) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U24 ( .A(mult_lsb_gf4_mul_2_2_n74), .B(
        mult_lsb_gf4_mul_2_2_n71), .Z(mult_lsb_gf4_mul_2_2_n73) );
  NOR2_X1 mult_lsb_gf4_mul_2_2_U23 ( .A1(mult_lsb_gf4_mul_2_2_n70), .A2(
        mult_lsb_gf4_mul_2_2_n69), .ZN(mult_lsb_gf4_mul_2_2_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U22 ( .A(InverterOutxD[10]), .B(
        InverterOutxD[11]), .ZN(mult_lsb_gf4_mul_2_2_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U21 ( .A(Y1_4xDP[10]), .B(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_2_2_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U20 ( .A(mult_lsb_gf4_mul_2_2_n68), .B(
        mult_lsb_gf4_mul_2_2_n67), .ZN(mult_lsb_FFxDN[33]) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U19 ( .A1(InverterOutxD[9]), .A2(Y1_4xDP[9]), 
        .ZN(mult_lsb_gf4_mul_2_2_n67) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U18 ( .A(mult_lsb_gf4_mul_2_2_n75), .B(
        mult_lsb_gf4_mul_2_2_n66), .Z(mult_lsb_gf4_mul_2_2_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U17 ( .A(mult_lsb_gf4_mul_2_2_n65), .B(
        mult_lsb_gf4_mul_2_2_n64), .ZN(mult_lsb_gf4_mul_2_2_n75) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U16 ( .A1(mult_lsb_gf4_mul_2_2_n63), .A2(
        mult_lsb_gf4_mul_2_2_n62), .ZN(mult_lsb_gf4_mul_2_2_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U15 ( .A(mult_lsb_gf4_mul_2_2_n61), .B(
        mult_lsb_gf4_mul_2_2_n60), .ZN(mult_lsb_gf4_mul_2_2_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U14 ( .A(mult_lsb_gf4_mul_2_2_n59), .B(
        mult_lsb_gf4_mul_2_2_n58), .ZN(mult_lsb_gf4_mul_2_2_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U13 ( .A(mult_lsb_gf4_mul_2_2_n57), .B(
        mult_lsb_gf4_mul_2_2_n56), .ZN(mult_lsb_FFxDN[32]) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U12 ( .A1(InverterOutxD[8]), .A2(Y1_4xDP[8]), 
        .ZN(mult_lsb_gf4_mul_2_2_n56) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U11 ( .A(mult_lsb_gf4_mul_2_2_n66), .B(
        mult_lsb_gf4_mul_2_2_n71), .Z(mult_lsb_gf4_mul_2_2_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U10 ( .A(mult_lsb_gf4_mul_2_2_n55), .B(
        mult_lsb_gf4_mul_2_2_n65), .ZN(mult_lsb_gf4_mul_2_2_n71) );
  NOR2_X1 mult_lsb_gf4_mul_2_2_U9 ( .A1(mult_lsb_gf4_mul_2_2_n61), .A2(
        mult_lsb_gf4_mul_2_2_n59), .ZN(mult_lsb_gf4_mul_2_2_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U8 ( .A(InverterOutxD[8]), .B(
        InverterOutxD[10]), .ZN(mult_lsb_gf4_mul_2_2_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U7 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_2_2_n61) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U6 ( .A1(mult_lsb_gf4_mul_2_2_n58), .A2(
        mult_lsb_gf4_mul_2_2_n60), .ZN(mult_lsb_gf4_mul_2_2_n55) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U5 ( .A(Y1_4xDP[9]), .B(Y1_4xDP[11]), .Z(
        mult_lsb_gf4_mul_2_2_n60) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U4 ( .A(InverterOutxD[9]), .B(InverterOutxD[11]), .Z(mult_lsb_gf4_mul_2_2_n58) );
  NOR2_X1 mult_lsb_gf4_mul_2_2_U3 ( .A1(mult_lsb_gf4_mul_2_2_n54), .A2(
        mult_lsb_gf4_mul_2_2_n53), .ZN(mult_lsb_gf4_mul_2_2_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U2 ( .A(InverterOutxD[8]), .B(InverterOutxD[9]), .ZN(mult_lsb_gf4_mul_2_2_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U1 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_2_2_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U29 ( .A(mult_lsb_gf4_mul_2_1_n77), .B(
        mult_lsb_gf4_mul_2_1_n76), .ZN(mult_lsb_Xi_mul_Yj_7__3_) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U28 ( .A1(InverterOutxD[11]), .A2(Y1_4xDP[7]), 
        .ZN(mult_lsb_gf4_mul_2_1_n76) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U27 ( .A(mult_lsb_gf4_mul_2_1_n75), .B(
        mult_lsb_gf4_mul_2_1_n74), .Z(mult_lsb_gf4_mul_2_1_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U26 ( .A(mult_lsb_gf4_mul_2_1_n73), .B(
        mult_lsb_gf4_mul_2_1_n72), .ZN(mult_lsb_Xi_mul_Yj_7__2_) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U25 ( .A1(InverterOutxD[10]), .A2(Y1_4xDP[6]), 
        .ZN(mult_lsb_gf4_mul_2_1_n72) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U24 ( .A(mult_lsb_gf4_mul_2_1_n74), .B(
        mult_lsb_gf4_mul_2_1_n71), .Z(mult_lsb_gf4_mul_2_1_n73) );
  NOR2_X1 mult_lsb_gf4_mul_2_1_U23 ( .A1(mult_lsb_gf4_mul_2_1_n70), .A2(
        mult_lsb_gf4_mul_2_1_n69), .ZN(mult_lsb_gf4_mul_2_1_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U22 ( .A(InverterOutxD[10]), .B(
        InverterOutxD[11]), .ZN(mult_lsb_gf4_mul_2_1_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U21 ( .A(Y1_4xDP[6]), .B(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_2_1_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U20 ( .A(mult_lsb_gf4_mul_2_1_n68), .B(
        mult_lsb_gf4_mul_2_1_n67), .ZN(mult_lsb_Xi_mul_Yj_7__1_) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U19 ( .A1(InverterOutxD[9]), .A2(Y1_4xDP[5]), 
        .ZN(mult_lsb_gf4_mul_2_1_n67) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U18 ( .A(mult_lsb_gf4_mul_2_1_n75), .B(
        mult_lsb_gf4_mul_2_1_n66), .Z(mult_lsb_gf4_mul_2_1_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U17 ( .A(mult_lsb_gf4_mul_2_1_n65), .B(
        mult_lsb_gf4_mul_2_1_n64), .ZN(mult_lsb_gf4_mul_2_1_n75) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U16 ( .A1(mult_lsb_gf4_mul_2_1_n63), .A2(
        mult_lsb_gf4_mul_2_1_n62), .ZN(mult_lsb_gf4_mul_2_1_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U15 ( .A(mult_lsb_gf4_mul_2_1_n61), .B(
        mult_lsb_gf4_mul_2_1_n60), .ZN(mult_lsb_gf4_mul_2_1_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U14 ( .A(mult_lsb_gf4_mul_2_1_n59), .B(
        mult_lsb_gf4_mul_2_1_n58), .ZN(mult_lsb_gf4_mul_2_1_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U13 ( .A(mult_lsb_gf4_mul_2_1_n57), .B(
        mult_lsb_gf4_mul_2_1_n56), .ZN(mult_lsb_Xi_mul_Yj_7__0_) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U12 ( .A1(InverterOutxD[8]), .A2(Y1_4xDP[4]), 
        .ZN(mult_lsb_gf4_mul_2_1_n56) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U11 ( .A(mult_lsb_gf4_mul_2_1_n66), .B(
        mult_lsb_gf4_mul_2_1_n71), .Z(mult_lsb_gf4_mul_2_1_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U10 ( .A(mult_lsb_gf4_mul_2_1_n55), .B(
        mult_lsb_gf4_mul_2_1_n65), .ZN(mult_lsb_gf4_mul_2_1_n71) );
  NOR2_X1 mult_lsb_gf4_mul_2_1_U9 ( .A1(mult_lsb_gf4_mul_2_1_n61), .A2(
        mult_lsb_gf4_mul_2_1_n59), .ZN(mult_lsb_gf4_mul_2_1_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U8 ( .A(InverterOutxD[8]), .B(
        InverterOutxD[10]), .ZN(mult_lsb_gf4_mul_2_1_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U7 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_2_1_n61) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U6 ( .A1(mult_lsb_gf4_mul_2_1_n58), .A2(
        mult_lsb_gf4_mul_2_1_n60), .ZN(mult_lsb_gf4_mul_2_1_n55) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U5 ( .A(Y1_4xDP[5]), .B(Y1_4xDP[7]), .Z(
        mult_lsb_gf4_mul_2_1_n60) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U4 ( .A(InverterOutxD[9]), .B(InverterOutxD[11]), .Z(mult_lsb_gf4_mul_2_1_n58) );
  NOR2_X1 mult_lsb_gf4_mul_2_1_U3 ( .A1(mult_lsb_gf4_mul_2_1_n54), .A2(
        mult_lsb_gf4_mul_2_1_n53), .ZN(mult_lsb_gf4_mul_2_1_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U2 ( .A(InverterOutxD[8]), .B(InverterOutxD[9]), .ZN(mult_lsb_gf4_mul_2_1_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U1 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_2_1_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U29 ( .A(mult_lsb_gf4_mul_2_0_n77), .B(
        mult_lsb_gf4_mul_2_0_n76), .ZN(mult_lsb_Xi_mul_Yj_6__3_) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U28 ( .A1(InverterOutxD[11]), .A2(Y1_4xDP[3]), 
        .ZN(mult_lsb_gf4_mul_2_0_n76) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U27 ( .A(mult_lsb_gf4_mul_2_0_n75), .B(
        mult_lsb_gf4_mul_2_0_n74), .Z(mult_lsb_gf4_mul_2_0_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U26 ( .A(mult_lsb_gf4_mul_2_0_n73), .B(
        mult_lsb_gf4_mul_2_0_n72), .ZN(mult_lsb_Xi_mul_Yj_6__2_) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U25 ( .A1(InverterOutxD[10]), .A2(Y1_4xDP[2]), 
        .ZN(mult_lsb_gf4_mul_2_0_n72) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U24 ( .A(mult_lsb_gf4_mul_2_0_n74), .B(
        mult_lsb_gf4_mul_2_0_n71), .Z(mult_lsb_gf4_mul_2_0_n73) );
  NOR2_X1 mult_lsb_gf4_mul_2_0_U23 ( .A1(mult_lsb_gf4_mul_2_0_n70), .A2(
        mult_lsb_gf4_mul_2_0_n69), .ZN(mult_lsb_gf4_mul_2_0_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U22 ( .A(InverterOutxD[10]), .B(
        InverterOutxD[11]), .ZN(mult_lsb_gf4_mul_2_0_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U21 ( .A(Y1_4xDP[2]), .B(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_2_0_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U20 ( .A(mult_lsb_gf4_mul_2_0_n68), .B(
        mult_lsb_gf4_mul_2_0_n67), .ZN(mult_lsb_Xi_mul_Yj_6__1_) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U19 ( .A1(InverterOutxD[9]), .A2(Y1_4xDP[1]), 
        .ZN(mult_lsb_gf4_mul_2_0_n67) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U18 ( .A(mult_lsb_gf4_mul_2_0_n75), .B(
        mult_lsb_gf4_mul_2_0_n66), .Z(mult_lsb_gf4_mul_2_0_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U17 ( .A(mult_lsb_gf4_mul_2_0_n65), .B(
        mult_lsb_gf4_mul_2_0_n64), .ZN(mult_lsb_gf4_mul_2_0_n75) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U16 ( .A1(mult_lsb_gf4_mul_2_0_n63), .A2(
        mult_lsb_gf4_mul_2_0_n62), .ZN(mult_lsb_gf4_mul_2_0_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U15 ( .A(mult_lsb_gf4_mul_2_0_n61), .B(
        mult_lsb_gf4_mul_2_0_n60), .ZN(mult_lsb_gf4_mul_2_0_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U14 ( .A(mult_lsb_gf4_mul_2_0_n59), .B(
        mult_lsb_gf4_mul_2_0_n58), .ZN(mult_lsb_gf4_mul_2_0_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U13 ( .A(mult_lsb_gf4_mul_2_0_n57), .B(
        mult_lsb_gf4_mul_2_0_n56), .ZN(mult_lsb_Xi_mul_Yj_6__0_) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U12 ( .A1(InverterOutxD[8]), .A2(Y1_4xDP[0]), 
        .ZN(mult_lsb_gf4_mul_2_0_n56) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U11 ( .A(mult_lsb_gf4_mul_2_0_n66), .B(
        mult_lsb_gf4_mul_2_0_n71), .Z(mult_lsb_gf4_mul_2_0_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U10 ( .A(mult_lsb_gf4_mul_2_0_n55), .B(
        mult_lsb_gf4_mul_2_0_n65), .ZN(mult_lsb_gf4_mul_2_0_n71) );
  NOR2_X1 mult_lsb_gf4_mul_2_0_U9 ( .A1(mult_lsb_gf4_mul_2_0_n61), .A2(
        mult_lsb_gf4_mul_2_0_n59), .ZN(mult_lsb_gf4_mul_2_0_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U8 ( .A(InverterOutxD[8]), .B(
        InverterOutxD[10]), .ZN(mult_lsb_gf4_mul_2_0_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U7 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_2_0_n61) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U6 ( .A1(mult_lsb_gf4_mul_2_0_n58), .A2(
        mult_lsb_gf4_mul_2_0_n60), .ZN(mult_lsb_gf4_mul_2_0_n55) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U5 ( .A(Y1_4xDP[1]), .B(Y1_4xDP[3]), .Z(
        mult_lsb_gf4_mul_2_0_n60) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U4 ( .A(InverterOutxD[9]), .B(InverterOutxD[11]), .Z(mult_lsb_gf4_mul_2_0_n58) );
  NOR2_X1 mult_lsb_gf4_mul_2_0_U3 ( .A1(mult_lsb_gf4_mul_2_0_n54), .A2(
        mult_lsb_gf4_mul_2_0_n53), .ZN(mult_lsb_gf4_mul_2_0_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U2 ( .A(InverterOutxD[8]), .B(InverterOutxD[9]), .ZN(mult_lsb_gf4_mul_2_0_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U1 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_2_0_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U29 ( .A(mult_lsb_gf4_mul_1_2_n77), .B(
        mult_lsb_gf4_mul_1_2_n76), .ZN(mult_lsb_Xi_mul_Yj_5__3_) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U28 ( .A1(InverterOutxD[7]), .A2(Y1_4xDP[11]), 
        .ZN(mult_lsb_gf4_mul_1_2_n76) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U27 ( .A(mult_lsb_gf4_mul_1_2_n75), .B(
        mult_lsb_gf4_mul_1_2_n74), .Z(mult_lsb_gf4_mul_1_2_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U26 ( .A(mult_lsb_gf4_mul_1_2_n73), .B(
        mult_lsb_gf4_mul_1_2_n72), .ZN(mult_lsb_Xi_mul_Yj_5__2_) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U25 ( .A1(InverterOutxD[6]), .A2(Y1_4xDP[10]), 
        .ZN(mult_lsb_gf4_mul_1_2_n72) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U24 ( .A(mult_lsb_gf4_mul_1_2_n74), .B(
        mult_lsb_gf4_mul_1_2_n71), .Z(mult_lsb_gf4_mul_1_2_n73) );
  NOR2_X1 mult_lsb_gf4_mul_1_2_U23 ( .A1(mult_lsb_gf4_mul_1_2_n70), .A2(
        mult_lsb_gf4_mul_1_2_n69), .ZN(mult_lsb_gf4_mul_1_2_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U22 ( .A(InverterOutxD[6]), .B(
        InverterOutxD[7]), .ZN(mult_lsb_gf4_mul_1_2_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U21 ( .A(Y1_4xDP[10]), .B(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_1_2_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U20 ( .A(mult_lsb_gf4_mul_1_2_n68), .B(
        mult_lsb_gf4_mul_1_2_n67), .ZN(mult_lsb_Xi_mul_Yj_5__1_) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U19 ( .A1(InverterOutxD[5]), .A2(Y1_4xDP[9]), 
        .ZN(mult_lsb_gf4_mul_1_2_n67) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U18 ( .A(mult_lsb_gf4_mul_1_2_n75), .B(
        mult_lsb_gf4_mul_1_2_n66), .Z(mult_lsb_gf4_mul_1_2_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U17 ( .A(mult_lsb_gf4_mul_1_2_n65), .B(
        mult_lsb_gf4_mul_1_2_n64), .ZN(mult_lsb_gf4_mul_1_2_n75) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U16 ( .A1(mult_lsb_gf4_mul_1_2_n63), .A2(
        mult_lsb_gf4_mul_1_2_n62), .ZN(mult_lsb_gf4_mul_1_2_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U15 ( .A(mult_lsb_gf4_mul_1_2_n61), .B(
        mult_lsb_gf4_mul_1_2_n60), .ZN(mult_lsb_gf4_mul_1_2_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U14 ( .A(mult_lsb_gf4_mul_1_2_n59), .B(
        mult_lsb_gf4_mul_1_2_n58), .ZN(mult_lsb_gf4_mul_1_2_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U13 ( .A(mult_lsb_gf4_mul_1_2_n57), .B(
        mult_lsb_gf4_mul_1_2_n56), .ZN(mult_lsb_Xi_mul_Yj_5__0_) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U12 ( .A1(InverterOutxD[4]), .A2(Y1_4xDP[8]), 
        .ZN(mult_lsb_gf4_mul_1_2_n56) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U11 ( .A(mult_lsb_gf4_mul_1_2_n66), .B(
        mult_lsb_gf4_mul_1_2_n71), .Z(mult_lsb_gf4_mul_1_2_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U10 ( .A(mult_lsb_gf4_mul_1_2_n55), .B(
        mult_lsb_gf4_mul_1_2_n65), .ZN(mult_lsb_gf4_mul_1_2_n71) );
  NOR2_X1 mult_lsb_gf4_mul_1_2_U9 ( .A1(mult_lsb_gf4_mul_1_2_n61), .A2(
        mult_lsb_gf4_mul_1_2_n59), .ZN(mult_lsb_gf4_mul_1_2_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U8 ( .A(InverterOutxD[4]), .B(InverterOutxD[6]), .ZN(mult_lsb_gf4_mul_1_2_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U7 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_1_2_n61) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U6 ( .A1(mult_lsb_gf4_mul_1_2_n58), .A2(
        mult_lsb_gf4_mul_1_2_n60), .ZN(mult_lsb_gf4_mul_1_2_n55) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U5 ( .A(Y1_4xDP[9]), .B(Y1_4xDP[11]), .Z(
        mult_lsb_gf4_mul_1_2_n60) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U4 ( .A(InverterOutxD[5]), .B(InverterOutxD[7]), 
        .Z(mult_lsb_gf4_mul_1_2_n58) );
  NOR2_X1 mult_lsb_gf4_mul_1_2_U3 ( .A1(mult_lsb_gf4_mul_1_2_n54), .A2(
        mult_lsb_gf4_mul_1_2_n53), .ZN(mult_lsb_gf4_mul_1_2_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U2 ( .A(InverterOutxD[4]), .B(InverterOutxD[5]), .ZN(mult_lsb_gf4_mul_1_2_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U1 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_1_2_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U29 ( .A(mult_lsb_gf4_mul_1_1_n77), .B(
        mult_lsb_gf4_mul_1_1_n76), .ZN(mult_lsb_FFxDN[19]) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U28 ( .A1(InverterOutxD[7]), .A2(Y1_4xDP[7]), 
        .ZN(mult_lsb_gf4_mul_1_1_n76) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U27 ( .A(mult_lsb_gf4_mul_1_1_n75), .B(
        mult_lsb_gf4_mul_1_1_n74), .Z(mult_lsb_gf4_mul_1_1_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U26 ( .A(mult_lsb_gf4_mul_1_1_n73), .B(
        mult_lsb_gf4_mul_1_1_n72), .ZN(mult_lsb_FFxDN[18]) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U25 ( .A1(InverterOutxD[6]), .A2(Y1_4xDP[6]), 
        .ZN(mult_lsb_gf4_mul_1_1_n72) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U24 ( .A(mult_lsb_gf4_mul_1_1_n74), .B(
        mult_lsb_gf4_mul_1_1_n71), .Z(mult_lsb_gf4_mul_1_1_n73) );
  NOR2_X1 mult_lsb_gf4_mul_1_1_U23 ( .A1(mult_lsb_gf4_mul_1_1_n70), .A2(
        mult_lsb_gf4_mul_1_1_n69), .ZN(mult_lsb_gf4_mul_1_1_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U22 ( .A(InverterOutxD[6]), .B(
        InverterOutxD[7]), .ZN(mult_lsb_gf4_mul_1_1_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U21 ( .A(Y1_4xDP[6]), .B(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_1_1_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U20 ( .A(mult_lsb_gf4_mul_1_1_n68), .B(
        mult_lsb_gf4_mul_1_1_n67), .ZN(mult_lsb_FFxDN[17]) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U19 ( .A1(InverterOutxD[5]), .A2(Y1_4xDP[5]), 
        .ZN(mult_lsb_gf4_mul_1_1_n67) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U18 ( .A(mult_lsb_gf4_mul_1_1_n75), .B(
        mult_lsb_gf4_mul_1_1_n66), .Z(mult_lsb_gf4_mul_1_1_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U17 ( .A(mult_lsb_gf4_mul_1_1_n65), .B(
        mult_lsb_gf4_mul_1_1_n64), .ZN(mult_lsb_gf4_mul_1_1_n75) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U16 ( .A1(mult_lsb_gf4_mul_1_1_n63), .A2(
        mult_lsb_gf4_mul_1_1_n62), .ZN(mult_lsb_gf4_mul_1_1_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U15 ( .A(mult_lsb_gf4_mul_1_1_n61), .B(
        mult_lsb_gf4_mul_1_1_n60), .ZN(mult_lsb_gf4_mul_1_1_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U14 ( .A(mult_lsb_gf4_mul_1_1_n59), .B(
        mult_lsb_gf4_mul_1_1_n58), .ZN(mult_lsb_gf4_mul_1_1_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U13 ( .A(mult_lsb_gf4_mul_1_1_n57), .B(
        mult_lsb_gf4_mul_1_1_n56), .ZN(mult_lsb_FFxDN[16]) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U12 ( .A1(InverterOutxD[4]), .A2(Y1_4xDP[4]), 
        .ZN(mult_lsb_gf4_mul_1_1_n56) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U11 ( .A(mult_lsb_gf4_mul_1_1_n66), .B(
        mult_lsb_gf4_mul_1_1_n71), .Z(mult_lsb_gf4_mul_1_1_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U10 ( .A(mult_lsb_gf4_mul_1_1_n55), .B(
        mult_lsb_gf4_mul_1_1_n65), .ZN(mult_lsb_gf4_mul_1_1_n71) );
  NOR2_X1 mult_lsb_gf4_mul_1_1_U9 ( .A1(mult_lsb_gf4_mul_1_1_n61), .A2(
        mult_lsb_gf4_mul_1_1_n59), .ZN(mult_lsb_gf4_mul_1_1_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U8 ( .A(InverterOutxD[4]), .B(InverterOutxD[6]), .ZN(mult_lsb_gf4_mul_1_1_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U7 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_1_1_n61) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U6 ( .A1(mult_lsb_gf4_mul_1_1_n58), .A2(
        mult_lsb_gf4_mul_1_1_n60), .ZN(mult_lsb_gf4_mul_1_1_n55) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U5 ( .A(Y1_4xDP[5]), .B(Y1_4xDP[7]), .Z(
        mult_lsb_gf4_mul_1_1_n60) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U4 ( .A(InverterOutxD[5]), .B(InverterOutxD[7]), 
        .Z(mult_lsb_gf4_mul_1_1_n58) );
  NOR2_X1 mult_lsb_gf4_mul_1_1_U3 ( .A1(mult_lsb_gf4_mul_1_1_n54), .A2(
        mult_lsb_gf4_mul_1_1_n53), .ZN(mult_lsb_gf4_mul_1_1_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U2 ( .A(InverterOutxD[4]), .B(InverterOutxD[5]), .ZN(mult_lsb_gf4_mul_1_1_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U1 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_1_1_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U29 ( .A(mult_lsb_gf4_mul_1_0_n77), .B(
        mult_lsb_gf4_mul_1_0_n76), .ZN(mult_lsb_Xi_mul_Yj_3__3_) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U28 ( .A1(InverterOutxD[7]), .A2(Y1_4xDP[3]), 
        .ZN(mult_lsb_gf4_mul_1_0_n76) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U27 ( .A(mult_lsb_gf4_mul_1_0_n75), .B(
        mult_lsb_gf4_mul_1_0_n74), .Z(mult_lsb_gf4_mul_1_0_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U26 ( .A(mult_lsb_gf4_mul_1_0_n73), .B(
        mult_lsb_gf4_mul_1_0_n72), .ZN(mult_lsb_Xi_mul_Yj_3__2_) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U25 ( .A1(InverterOutxD[6]), .A2(Y1_4xDP[2]), 
        .ZN(mult_lsb_gf4_mul_1_0_n72) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U24 ( .A(mult_lsb_gf4_mul_1_0_n74), .B(
        mult_lsb_gf4_mul_1_0_n71), .Z(mult_lsb_gf4_mul_1_0_n73) );
  NOR2_X1 mult_lsb_gf4_mul_1_0_U23 ( .A1(mult_lsb_gf4_mul_1_0_n70), .A2(
        mult_lsb_gf4_mul_1_0_n69), .ZN(mult_lsb_gf4_mul_1_0_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U22 ( .A(InverterOutxD[6]), .B(
        InverterOutxD[7]), .ZN(mult_lsb_gf4_mul_1_0_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U21 ( .A(Y1_4xDP[2]), .B(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_1_0_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U20 ( .A(mult_lsb_gf4_mul_1_0_n68), .B(
        mult_lsb_gf4_mul_1_0_n67), .ZN(mult_lsb_Xi_mul_Yj_3__1_) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U19 ( .A1(InverterOutxD[5]), .A2(Y1_4xDP[1]), 
        .ZN(mult_lsb_gf4_mul_1_0_n67) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U18 ( .A(mult_lsb_gf4_mul_1_0_n75), .B(
        mult_lsb_gf4_mul_1_0_n66), .Z(mult_lsb_gf4_mul_1_0_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U17 ( .A(mult_lsb_gf4_mul_1_0_n65), .B(
        mult_lsb_gf4_mul_1_0_n64), .ZN(mult_lsb_gf4_mul_1_0_n75) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U16 ( .A1(mult_lsb_gf4_mul_1_0_n63), .A2(
        mult_lsb_gf4_mul_1_0_n62), .ZN(mult_lsb_gf4_mul_1_0_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U15 ( .A(mult_lsb_gf4_mul_1_0_n61), .B(
        mult_lsb_gf4_mul_1_0_n60), .ZN(mult_lsb_gf4_mul_1_0_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U14 ( .A(mult_lsb_gf4_mul_1_0_n59), .B(
        mult_lsb_gf4_mul_1_0_n58), .ZN(mult_lsb_gf4_mul_1_0_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U13 ( .A(mult_lsb_gf4_mul_1_0_n57), .B(
        mult_lsb_gf4_mul_1_0_n56), .ZN(mult_lsb_Xi_mul_Yj_3__0_) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U12 ( .A1(InverterOutxD[4]), .A2(Y1_4xDP[0]), 
        .ZN(mult_lsb_gf4_mul_1_0_n56) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U11 ( .A(mult_lsb_gf4_mul_1_0_n66), .B(
        mult_lsb_gf4_mul_1_0_n71), .Z(mult_lsb_gf4_mul_1_0_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U10 ( .A(mult_lsb_gf4_mul_1_0_n55), .B(
        mult_lsb_gf4_mul_1_0_n65), .ZN(mult_lsb_gf4_mul_1_0_n71) );
  NOR2_X1 mult_lsb_gf4_mul_1_0_U9 ( .A1(mult_lsb_gf4_mul_1_0_n61), .A2(
        mult_lsb_gf4_mul_1_0_n59), .ZN(mult_lsb_gf4_mul_1_0_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U8 ( .A(InverterOutxD[4]), .B(InverterOutxD[6]), .ZN(mult_lsb_gf4_mul_1_0_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U7 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_1_0_n61) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U6 ( .A1(mult_lsb_gf4_mul_1_0_n58), .A2(
        mult_lsb_gf4_mul_1_0_n60), .ZN(mult_lsb_gf4_mul_1_0_n55) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U5 ( .A(Y1_4xDP[1]), .B(Y1_4xDP[3]), .Z(
        mult_lsb_gf4_mul_1_0_n60) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U4 ( .A(InverterOutxD[5]), .B(InverterOutxD[7]), 
        .Z(mult_lsb_gf4_mul_1_0_n58) );
  NOR2_X1 mult_lsb_gf4_mul_1_0_U3 ( .A1(mult_lsb_gf4_mul_1_0_n54), .A2(
        mult_lsb_gf4_mul_1_0_n53), .ZN(mult_lsb_gf4_mul_1_0_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U2 ( .A(InverterOutxD[4]), .B(InverterOutxD[5]), .ZN(mult_lsb_gf4_mul_1_0_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U1 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_1_0_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U29 ( .A(mult_lsb_gf4_mul_0_2_n77), .B(
        mult_lsb_gf4_mul_0_2_n76), .ZN(mult_lsb_Xi_mul_Yj_2__3_) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U28 ( .A1(InverterOutxD[3]), .A2(Y1_4xDP[11]), 
        .ZN(mult_lsb_gf4_mul_0_2_n76) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U27 ( .A(mult_lsb_gf4_mul_0_2_n75), .B(
        mult_lsb_gf4_mul_0_2_n74), .Z(mult_lsb_gf4_mul_0_2_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U26 ( .A(mult_lsb_gf4_mul_0_2_n73), .B(
        mult_lsb_gf4_mul_0_2_n72), .ZN(mult_lsb_Xi_mul_Yj_2__2_) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U25 ( .A1(InverterOutxD[2]), .A2(Y1_4xDP[10]), 
        .ZN(mult_lsb_gf4_mul_0_2_n72) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U24 ( .A(mult_lsb_gf4_mul_0_2_n74), .B(
        mult_lsb_gf4_mul_0_2_n71), .Z(mult_lsb_gf4_mul_0_2_n73) );
  NOR2_X1 mult_lsb_gf4_mul_0_2_U23 ( .A1(mult_lsb_gf4_mul_0_2_n70), .A2(
        mult_lsb_gf4_mul_0_2_n69), .ZN(mult_lsb_gf4_mul_0_2_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U22 ( .A(InverterOutxD[2]), .B(
        InverterOutxD[3]), .ZN(mult_lsb_gf4_mul_0_2_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U21 ( .A(Y1_4xDP[10]), .B(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_0_2_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U20 ( .A(mult_lsb_gf4_mul_0_2_n68), .B(
        mult_lsb_gf4_mul_0_2_n67), .ZN(mult_lsb_Xi_mul_Yj_2__1_) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U19 ( .A1(InverterOutxD[1]), .A2(Y1_4xDP[9]), 
        .ZN(mult_lsb_gf4_mul_0_2_n67) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U18 ( .A(mult_lsb_gf4_mul_0_2_n75), .B(
        mult_lsb_gf4_mul_0_2_n66), .Z(mult_lsb_gf4_mul_0_2_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U17 ( .A(mult_lsb_gf4_mul_0_2_n65), .B(
        mult_lsb_gf4_mul_0_2_n64), .ZN(mult_lsb_gf4_mul_0_2_n75) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U16 ( .A1(mult_lsb_gf4_mul_0_2_n63), .A2(
        mult_lsb_gf4_mul_0_2_n62), .ZN(mult_lsb_gf4_mul_0_2_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U15 ( .A(mult_lsb_gf4_mul_0_2_n61), .B(
        mult_lsb_gf4_mul_0_2_n60), .ZN(mult_lsb_gf4_mul_0_2_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U14 ( .A(mult_lsb_gf4_mul_0_2_n59), .B(
        mult_lsb_gf4_mul_0_2_n58), .ZN(mult_lsb_gf4_mul_0_2_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U13 ( .A(mult_lsb_gf4_mul_0_2_n57), .B(
        mult_lsb_gf4_mul_0_2_n56), .ZN(mult_lsb_Xi_mul_Yj_2__0_) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U12 ( .A1(InverterOutxD[0]), .A2(Y1_4xDP[8]), 
        .ZN(mult_lsb_gf4_mul_0_2_n56) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U11 ( .A(mult_lsb_gf4_mul_0_2_n66), .B(
        mult_lsb_gf4_mul_0_2_n71), .Z(mult_lsb_gf4_mul_0_2_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U10 ( .A(mult_lsb_gf4_mul_0_2_n55), .B(
        mult_lsb_gf4_mul_0_2_n65), .ZN(mult_lsb_gf4_mul_0_2_n71) );
  NOR2_X1 mult_lsb_gf4_mul_0_2_U9 ( .A1(mult_lsb_gf4_mul_0_2_n61), .A2(
        mult_lsb_gf4_mul_0_2_n59), .ZN(mult_lsb_gf4_mul_0_2_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U8 ( .A(InverterOutxD[0]), .B(InverterOutxD[2]), .ZN(mult_lsb_gf4_mul_0_2_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U7 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_0_2_n61) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U6 ( .A1(mult_lsb_gf4_mul_0_2_n58), .A2(
        mult_lsb_gf4_mul_0_2_n60), .ZN(mult_lsb_gf4_mul_0_2_n55) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U5 ( .A(Y1_4xDP[9]), .B(Y1_4xDP[11]), .Z(
        mult_lsb_gf4_mul_0_2_n60) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U4 ( .A(InverterOutxD[1]), .B(InverterOutxD[3]), 
        .Z(mult_lsb_gf4_mul_0_2_n58) );
  NOR2_X1 mult_lsb_gf4_mul_0_2_U3 ( .A1(mult_lsb_gf4_mul_0_2_n54), .A2(
        mult_lsb_gf4_mul_0_2_n53), .ZN(mult_lsb_gf4_mul_0_2_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U2 ( .A(InverterOutxD[0]), .B(InverterOutxD[1]), .ZN(mult_lsb_gf4_mul_0_2_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U1 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_0_2_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U29 ( .A(mult_lsb_gf4_mul_0_1_n77), .B(
        mult_lsb_gf4_mul_0_1_n76), .ZN(mult_lsb_Xi_mul_Yj_1__3_) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U28 ( .A1(InverterOutxD[3]), .A2(Y1_4xDP[7]), 
        .ZN(mult_lsb_gf4_mul_0_1_n76) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U27 ( .A(mult_lsb_gf4_mul_0_1_n75), .B(
        mult_lsb_gf4_mul_0_1_n74), .Z(mult_lsb_gf4_mul_0_1_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U26 ( .A(mult_lsb_gf4_mul_0_1_n73), .B(
        mult_lsb_gf4_mul_0_1_n72), .ZN(mult_lsb_Xi_mul_Yj_1__2_) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U25 ( .A1(InverterOutxD[2]), .A2(Y1_4xDP[6]), 
        .ZN(mult_lsb_gf4_mul_0_1_n72) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U24 ( .A(mult_lsb_gf4_mul_0_1_n74), .B(
        mult_lsb_gf4_mul_0_1_n71), .Z(mult_lsb_gf4_mul_0_1_n73) );
  NOR2_X1 mult_lsb_gf4_mul_0_1_U23 ( .A1(mult_lsb_gf4_mul_0_1_n70), .A2(
        mult_lsb_gf4_mul_0_1_n69), .ZN(mult_lsb_gf4_mul_0_1_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U22 ( .A(InverterOutxD[2]), .B(
        InverterOutxD[3]), .ZN(mult_lsb_gf4_mul_0_1_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U21 ( .A(Y1_4xDP[6]), .B(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_0_1_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U20 ( .A(mult_lsb_gf4_mul_0_1_n68), .B(
        mult_lsb_gf4_mul_0_1_n67), .ZN(mult_lsb_Xi_mul_Yj_1__1_) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U19 ( .A1(InverterOutxD[1]), .A2(Y1_4xDP[5]), 
        .ZN(mult_lsb_gf4_mul_0_1_n67) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U18 ( .A(mult_lsb_gf4_mul_0_1_n75), .B(
        mult_lsb_gf4_mul_0_1_n66), .Z(mult_lsb_gf4_mul_0_1_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U17 ( .A(mult_lsb_gf4_mul_0_1_n65), .B(
        mult_lsb_gf4_mul_0_1_n64), .ZN(mult_lsb_gf4_mul_0_1_n75) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U16 ( .A1(mult_lsb_gf4_mul_0_1_n63), .A2(
        mult_lsb_gf4_mul_0_1_n62), .ZN(mult_lsb_gf4_mul_0_1_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U15 ( .A(mult_lsb_gf4_mul_0_1_n61), .B(
        mult_lsb_gf4_mul_0_1_n60), .ZN(mult_lsb_gf4_mul_0_1_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U14 ( .A(mult_lsb_gf4_mul_0_1_n59), .B(
        mult_lsb_gf4_mul_0_1_n58), .ZN(mult_lsb_gf4_mul_0_1_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U13 ( .A(mult_lsb_gf4_mul_0_1_n57), .B(
        mult_lsb_gf4_mul_0_1_n56), .ZN(mult_lsb_Xi_mul_Yj_1__0_) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U12 ( .A1(InverterOutxD[0]), .A2(Y1_4xDP[4]), 
        .ZN(mult_lsb_gf4_mul_0_1_n56) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U11 ( .A(mult_lsb_gf4_mul_0_1_n66), .B(
        mult_lsb_gf4_mul_0_1_n71), .Z(mult_lsb_gf4_mul_0_1_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U10 ( .A(mult_lsb_gf4_mul_0_1_n55), .B(
        mult_lsb_gf4_mul_0_1_n65), .ZN(mult_lsb_gf4_mul_0_1_n71) );
  NOR2_X1 mult_lsb_gf4_mul_0_1_U9 ( .A1(mult_lsb_gf4_mul_0_1_n61), .A2(
        mult_lsb_gf4_mul_0_1_n59), .ZN(mult_lsb_gf4_mul_0_1_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U8 ( .A(InverterOutxD[0]), .B(InverterOutxD[2]), .ZN(mult_lsb_gf4_mul_0_1_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U7 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_0_1_n61) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U6 ( .A1(mult_lsb_gf4_mul_0_1_n58), .A2(
        mult_lsb_gf4_mul_0_1_n60), .ZN(mult_lsb_gf4_mul_0_1_n55) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U5 ( .A(Y1_4xDP[5]), .B(Y1_4xDP[7]), .Z(
        mult_lsb_gf4_mul_0_1_n60) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U4 ( .A(InverterOutxD[1]), .B(InverterOutxD[3]), 
        .Z(mult_lsb_gf4_mul_0_1_n58) );
  NOR2_X1 mult_lsb_gf4_mul_0_1_U3 ( .A1(mult_lsb_gf4_mul_0_1_n54), .A2(
        mult_lsb_gf4_mul_0_1_n53), .ZN(mult_lsb_gf4_mul_0_1_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U2 ( .A(InverterOutxD[0]), .B(InverterOutxD[1]), .ZN(mult_lsb_gf4_mul_0_1_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U1 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_0_1_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U29 ( .A(mult_lsb_gf4_mul_0_0_n77), .B(
        mult_lsb_gf4_mul_0_0_n76), .ZN(mult_lsb_FFxDN[3]) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U28 ( .A1(InverterOutxD[3]), .A2(Y1_4xDP[3]), 
        .ZN(mult_lsb_gf4_mul_0_0_n76) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U27 ( .A(mult_lsb_gf4_mul_0_0_n75), .B(
        mult_lsb_gf4_mul_0_0_n74), .Z(mult_lsb_gf4_mul_0_0_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U26 ( .A(mult_lsb_gf4_mul_0_0_n73), .B(
        mult_lsb_gf4_mul_0_0_n72), .ZN(mult_lsb_FFxDN[2]) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U25 ( .A1(InverterOutxD[2]), .A2(Y1_4xDP[2]), 
        .ZN(mult_lsb_gf4_mul_0_0_n72) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U24 ( .A(mult_lsb_gf4_mul_0_0_n74), .B(
        mult_lsb_gf4_mul_0_0_n71), .Z(mult_lsb_gf4_mul_0_0_n73) );
  NOR2_X1 mult_lsb_gf4_mul_0_0_U23 ( .A1(mult_lsb_gf4_mul_0_0_n70), .A2(
        mult_lsb_gf4_mul_0_0_n69), .ZN(mult_lsb_gf4_mul_0_0_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U22 ( .A(InverterOutxD[2]), .B(
        InverterOutxD[3]), .ZN(mult_lsb_gf4_mul_0_0_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U21 ( .A(Y1_4xDP[2]), .B(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_0_0_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U20 ( .A(mult_lsb_gf4_mul_0_0_n68), .B(
        mult_lsb_gf4_mul_0_0_n67), .ZN(mult_lsb_FFxDN[1]) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U19 ( .A1(InverterOutxD[1]), .A2(Y1_4xDP[1]), 
        .ZN(mult_lsb_gf4_mul_0_0_n67) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U18 ( .A(mult_lsb_gf4_mul_0_0_n75), .B(
        mult_lsb_gf4_mul_0_0_n66), .Z(mult_lsb_gf4_mul_0_0_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U17 ( .A(mult_lsb_gf4_mul_0_0_n65), .B(
        mult_lsb_gf4_mul_0_0_n64), .ZN(mult_lsb_gf4_mul_0_0_n75) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U16 ( .A1(mult_lsb_gf4_mul_0_0_n63), .A2(
        mult_lsb_gf4_mul_0_0_n62), .ZN(mult_lsb_gf4_mul_0_0_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U15 ( .A(mult_lsb_gf4_mul_0_0_n61), .B(
        mult_lsb_gf4_mul_0_0_n60), .ZN(mult_lsb_gf4_mul_0_0_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U14 ( .A(mult_lsb_gf4_mul_0_0_n59), .B(
        mult_lsb_gf4_mul_0_0_n58), .ZN(mult_lsb_gf4_mul_0_0_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U13 ( .A(mult_lsb_gf4_mul_0_0_n57), .B(
        mult_lsb_gf4_mul_0_0_n56), .ZN(mult_lsb_FFxDN[0]) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U12 ( .A1(InverterOutxD[0]), .A2(Y1_4xDP[0]), 
        .ZN(mult_lsb_gf4_mul_0_0_n56) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U11 ( .A(mult_lsb_gf4_mul_0_0_n66), .B(
        mult_lsb_gf4_mul_0_0_n71), .Z(mult_lsb_gf4_mul_0_0_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U10 ( .A(mult_lsb_gf4_mul_0_0_n55), .B(
        mult_lsb_gf4_mul_0_0_n65), .ZN(mult_lsb_gf4_mul_0_0_n71) );
  NOR2_X1 mult_lsb_gf4_mul_0_0_U9 ( .A1(mult_lsb_gf4_mul_0_0_n61), .A2(
        mult_lsb_gf4_mul_0_0_n59), .ZN(mult_lsb_gf4_mul_0_0_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U8 ( .A(InverterOutxD[0]), .B(InverterOutxD[2]), .ZN(mult_lsb_gf4_mul_0_0_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U7 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_0_0_n61) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U6 ( .A1(mult_lsb_gf4_mul_0_0_n58), .A2(
        mult_lsb_gf4_mul_0_0_n60), .ZN(mult_lsb_gf4_mul_0_0_n55) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U5 ( .A(Y1_4xDP[1]), .B(Y1_4xDP[3]), .Z(
        mult_lsb_gf4_mul_0_0_n60) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U4 ( .A(InverterOutxD[1]), .B(InverterOutxD[3]), 
        .Z(mult_lsb_gf4_mul_0_0_n58) );
  NOR2_X1 mult_lsb_gf4_mul_0_0_U3 ( .A1(mult_lsb_gf4_mul_0_0_n54), .A2(
        mult_lsb_gf4_mul_0_0_n53), .ZN(mult_lsb_gf4_mul_0_0_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U2 ( .A(InverterOutxD[0]), .B(InverterOutxD[1]), .ZN(mult_lsb_gf4_mul_0_0_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U1 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_0_0_n54) );
endmodule

